PK   j
mWݵ�2>  ��    cirkitFile.json�}[�%�q�_1J�[e!yK2����~�%X��A3(�USpO�lu�d���f��S]y��/O0O�f��tU�� F����������s������ӧ�w�)w�c����z�����秏�/���\����w�?g/��s�5�~������ˣs6X[�Yߴ:�u�g��yV�NV����c~���:[S�]_Zj]��U����Y��Uk|�u���j�JYI k�,�nċ��9�9��s٪��Yg��U�ɕ+h�M�6mWd�(lf{�gU����:�M�h����� kn������}V�9�kCt�f��k�}|���ه�����\N��+��we�m��L]Z��$�9�h�ۦwY_Z/��lT��]��rZׅ�f ��nU�7��LI�,���yf�ЗM����,�@�9�V��}^�����lW��.��ja����%@�쑄�;	��fuV{�ɌW.��'Ȯt�6y�V�)[Ӳ*Z22G�d-�Q(Zq$
��(�ӽ��U�!�2Mf���`�:k��zG�k�B�Ӻ���m�h֢���|�N��]�t��U��{�y�+yc�/�מ�iۛ���/rOWeUgU��iڶ�$����,�hќE��K	h�F� �	Eh/���^Ⱥ{Y� �^ʺ�\�_	��
�����֟���l=I�:��@��R�E�JgN�A� ��uFH4��2�MC�N��YYu&���f�qN7un�U����-��s<��	�YW�}f-�P��ȼ�JZ��胒-O+Тq{��܊C�E
'c���$Qd�LL���h�U5�I$'�t�N�Z������V6g!���X*C�A��� �γ�;��V�2�91WD��Y�uF���i]��ߠ����UN�y� :��۲���m�ʘ�2�:�F2c�D�q��y��Z�j;[f%��B�*�Ӳ��?��@)�U�,S
X�4]y�Q��t�Ug��\Q��VG-7��� ˖��xJb��FV�=�,Ӛ�lL�u�������k^���C��,[n���ou�mFf�PvY�$�j��w�8��� dn�}����rbMN,�:W1o�ʔ�q�2&�dwv��ܜ��fO4vE,I�m�@��p��͂hL �۬�SUӄ����SY["����!�N�|Xh�F��'�1oi�,��E�T��]Y�s�Ȅ�,27�^�
UI��`�H&Q��K�,IYu�J�3C��ː���m8�N��q^䇺����{|�u��uΝ�Y���#�D�Y���1mո��}q.��'�J��:��Ŵ�;�D|�0��>I���%	u0}A�T�`.Q�$\�[���D��/�Ht��!�C]G���]��y�ڈ ���Z���[�=��`ޜp A.��n�V\qr	� -�"W����Kr�q���ɰ��Ӣ<Gu��m�ی��K�So��L���i����m�h�A��$����SQC�p��%�y'P�^&ͺ�!w�4g��VМ��I@��;�BZ�S4��@�	h^r��r$�9��E��B���?��%r�^��N([`��Dd�����y�3h��5ǎ@=�WLLK~/�Ǽ�bR�䅉c�m��&�<316Ɩ$��]��/zmM����l��$q�]V��f�z��&�(�x����,+i�Z�d��Y��5UF�m�4�d�����1����m� 2Gbm�IH7}fl�g6DVR�&���Z�����l���@l��E(I(l�W}ը��s�{C�[����� d^����5��[��ܲA�±2�t@&���`����F.C�2�9fFe
 �,�'�M���	�Y�}��� �h�9��7W<+�`lH��ܜ��]��A�g��@�m�����P�#VW>b�1?f��[m0�@��έ6��3d5�;g9 =��Q��b�1'dN�=��9�g.��̙��@'n���,I�5�>dI@s�10lGp�pD��	X ��d^�c"V� ��0��)#��_D�����	 �~$�m)@������ �~$ ���/�i����ӳ0��ݯ���q�B�&��*υ��$��$�حuA%E]F�:�(:	.&�(vk���:룠�r�g�潡Q�P�F����<0;�f�Y_4�L\��匓2�$�p�lS1�Hh���=Bs�����e4�J\�u!��=BS����F9�iכR0��F�$�'%$�L2�����z��'.I1���1Y�f��e��$	p��&4�H�Q�#es���!뫋�I0���9:��fu7O �}c}u�L	p��#4�F�Q654�Ć��H0��9B�BD\H�c��{fk��#0��ݯ<	�����$
�3B"��Mnp����WW�����(o�(js0��slPן`�M\�P���E��Q7
B���>
ھ>
���Gh���ꢑ�	pټ�8��l� 4*=�(i�eSf@�಩���	Ftsl�X�ЈԈKE<KBu����MqҐ�n���&�4$��а
[�p�f
��o��p���S�0޶�I�-�s\$�C�m�p�ẁ%\���a��Fh8�o�"�른�7y1��~{��t	p�[w�~�k[/1X�ن$K0ʶ%�Zgzh��:.h�Ն%��J0ʶU�m��S�������l
Wh�ƫ3M�`��p0@(�(n���$e���l�:08f�ׁ�.	pٜ��qO��$�00$�(����ؘH� ����/�h�B\�.w�n���%�@��l�]�A?�m����|�Q6� Qo��uA=����wQg��lR�?�`��$3ڴ/������N0�����꥓zA쾼<W�������$��$�حQ`/h�(��{A�G�\]�Z>��������G��|��=����l��-es]`/h�(��{A�GI�.�g����R$�'%$�LCu��7��4��ЯJC�j��a/h�(��{A�G��%�zu�Z>����^��Q6W�����y`/h�(�{{A�G��#�Z>���^��Q���z}]P/h�(�T�zA��{A�Gٜ���_@/h�(�������M/��|�M\`/h�(��zA�G��dQ/��Q`/h�(�3����lލ��|��u���壤Y�M���������^��Q6us�:�%"�4Ի���^�	�IC�ۺ9��`�44���JC�:�D<8�4T��P�NC�:�4T��P�NC�&�M*���壤�0ق^��Q +4��n}@���l[BP/���F��WG����u/�Z>ʶ6�zA���zA�Gٶ(�^��Q6o%�Z>��8�-e��zA�G쒠�:�B���lsL�z�c�^��Q��2��|�4�l[�P/h�(�3B����F�Z>J\�o{�Z>�&߅���l*I��|�Mz���壤�e�va/h�(�T{A�G٤:�Z>ʦb{A'������{����2A?>��y�������s������ǧ���������/��!���.dm-�:�
c详m���U�W\!���]S�"�A�}�@Y�ʔ��O�u���v!��2�v��â�ˬ�H�����r��ޙ�oM�U#�l�e���A�]^wM�&/��`�,x�L�Vhr[��酐�}� ��\�ʛ�X����$��YmB�馭��p��mr�An��ކL[C�htT"٭�T][�J�4w�!Ȗ��If�����!����i���"�θ�u1.��3�����}�EUt��hF�TE�Ua]����Ga�z��̬v[{뛐g͗��UV�C�s��P[ݭ�Y ��}_�d��!�u_�rݓ�mC�[��h�9C���mٜ���rބ�_vY�4����o�����]��9�P�B@a�ծuߨ�������'�8��=1(S��>f�{M�EoK*IV5.'�۪�MY5YFےSa�B~�9����3��eh��]��t#F��fu�w���hZ�֡��6t"5+�|령�RhV6� sٖ�,��!�6�?���v�`��5I�}Q���]���'\XR�w��@��Y�-�ꪐU$�Ғ�ti���!�*�ՠ~c�/�5Q���4��+�1yo3SF�����g�����h_����ɪ"� �A����PIsrG;���zr�m|?�+�ӶE�UQ$���1���c�ٜz�6�t`ڮӶoY�����9E����N� 3�/4g�<K Cs�'B%m�V�w�7��]C'۵*+�V�D�}U��@n����s�	��E�vWhJ_�<�M%�N"�3÷�9����� �V["�"u�Sd=5�j\�tzi��͊�T�Fm�fE��@��*l|Yet�+:�m��H�^U6�Mk���`�,��@���CF�>Fˀ�f���04f>` ��矬�!��2�	�u�V�6���d>:4ZKZU�z������H�}��%�9��]}UsY)ɜ�S�b�2gjF��3OGP$���esf��e �s˲>���6�z=dv�`���ϳ�������pK�q��C�e@0t�z�앁\���`d���(����X6�e!�Ĕ@�N��U��	�5�%HF�h�N�� �|r��f�L�' �Z��� ��#�ޒ�,7�@#�$���h,�M�ϲ�W��\�`����r d0�� ��� ̻s d0����=���&�ZH�{���-9��ey\��,,���K�>�Ci��}̤���Gl4�eYY1W%��Z"�p�1,�gdǒT^Oc��L�����UF��ݦ7Y(�&�iLgr�x�*X`d3��X�6�ŚK �Vv(>���7��t���1n�v-�n�Ό��BU�g�+h�X�
�MS#�j⊕u�:Z_K�CP�����5��Eh0g0f��L��e���⦯����}��X��a������a����x
���pd,n�Ű��(\���,��8;�_����~���@�<D�>^����h���LU\M��&�x/Ȓ9��S�l��8��L�!Ym�q��8�X���3dLL��G���AuY�(��*J��|�\��1Y	٧�sCh���%�)�����Ȳw+ٜ%ou`�F�6�.�:ˍ3$ř&��>k�is_�z�\Ho�R�a-�3�ڲ9�|��̞*0��y������CƼ���
%`��N%��y '�y�Bxs�0ǯ�d�2�)��C|0��:�3�JW�pY[�(�(I��*��im��sOɜ!�2
㬀�C�RY�V[�� �29L�C^��6����@K�����E/���9�(Ƶ�gM�D�ҐAfvZ��>��$���t�\ZhB�n-0��{Af��̫ߘ
f�=���)Y`�`b��r�����"��Q���dw��W�� K��8 �,p@�'��~��֌���y�r�,�KR���O����c������#5��	o>>�a�g9��r�	���#,+�?$!��]�c#���En����c���^E���W�E�n�%��A�7����W�E��un�F\��l�B"�B� �[d5�3"a�k�1�8_E���y"���o�-R��#p����H��w�2�A6�����-@S�3[�ͮ�MpXC�&I��=@�XV1�77�vk �@��_��0y��
���i��}W���+�Ѝ���SXE�e�-����f*������MT1����m�e7��q��-���nPoc�[��X�NnP}C�	�E8C ��!G@X��0�����:C �|��	oP�C�ª��&7(�!�a��TX��0Њr��=C �ﱎ�-�|�bp�jrV$Lg���-j�8�����&��F�S(F@��p�E����Nev21R[�1+^��&�骙�����*vG(�d��K�?t-L����WB~ϸ��qm�Cu;�^�\�_Lu<N� ���>�	�������1R���(F��q�W�H_��oSG���~�I�ȯG����:R����'�W������6,(�z�V�&��k��o���YIH� =P��I.#���Q�1�2&>���o˛n�(�+G@�+m�[�ꕯ��b�ar�UnQ�W��2��ܢ���)�AQ����+G@X�w�[T��# L���@z���	0���c ��ΌoPX���&�ii`9+F�h��-�����1����U8�z��F>4'�aIa9+�9����a��3|h���n���a�ŇC ��t���H��	0&^gƷ�O|�I�ǋ�j��Է(Z|�����#���i%c�X$,h��G|����&��7^߃T9�# ,v���-j���ߠ�1�~���G�a���u���J�w������7���+B�82������ՠI!_�[��9�~�[��&럂	vF�h��c� ���4 $]�E�u��u���A9s�P*�j���-����Y��P���}C��1��0֥0W
��#6�Xo��M��e"�r�z�B9޺���DA�,B���W���8=��&@�H��-k��[�%��v)xd ����F&���6�!2�F������%��!����9w��ˊF�F�� ������kS�r��� �>�����J��C��)$��.��b1�w[a?7p':pv�4]�N$��@̉�wx�%��y�g��XY������F�1�Iԑi��`��r����
�����\,t�z �*���@������r�LF��x���zgZ�G���Cp�e��|[=Dp��(�-`��-!�d�����82�N �7��-����� ��;��	6�� �B��������f!�W���qDx��(ȷ�&!�)�	'<2$�� �t�
����2�aek�^��Λ��M���d #B��ft��O�8_�=[p�P��%�1�@�'t�Q������S��~��ڶ��n3�ʊ�i�ִ1%��u=Q���b���@���|�p�R�B W�ot��D�s�Cs�0@�!�$4�[�zW�U�"p���j�0��S9;KA��~'ӭ�Ƒ�{��!\��	yIlF���+ ��mUQ ��(R�jR]]l3:�ob.#p$�O I��u�rζMﲾ0:����Fe}ݕ�(G��ǭ�QuB`ӷJ��ClIƇ#�Ua[�o�r	!�$1'@$IL��VB�ǾhI�4���e�qh�e�˼���g��j�V��K����\A��Ib�䴔=yJ����|��%�I���z�7Hax`8 ��q��$���(M^��P8Ar�$y�Aޙ�[��_�p��@"����������O��_����ן?��i�ǗO�_�ڻ���L���]>�c��L�2��h8M�=��
��XƊF�͆�d�[X{�{�|�-����x6��=�
%�W,O`r�:|�$5:;0�t8-�n����f�F�T_f�1,�g�I����cvLy��X�a6#�qwI�[X;���Ef�I
Y̹9W8��	�_�{a� �_
��\:���"n`� +�6�
����ș��b�Y�;����ӳ#/Age���3��[�W��<�04�;�;��ٌ�$�I�~堀�"f{���A����fY���uSQ��I�K�X>tT���ú��|ƕ��N�R�NL�?�,#��%�ɂE<�ɂ�f�e<=9c���͆c��n	3x,Rs���R��n�_��ѵ3ΆcN�;�Kt�Μ���XOt8� ���D�n�&���� ��|e9��Pa���C���_]�s��4܊� �b% �|�n4I�r>�0�'j��Ɠ�I@J�k&l��@J���u-�D�5З�F���d�i h*T�F�q��cd1��*�%0���1}C@���'�}5]���Q�:Z\5�cW�T&1+|t�@�`r=T( k_��(X��A���
J��r���I��a�j��Lt=S�Bwφ�2La9ē�`�X���Lh�L�X-�v�y+2���!í�P��,�#���#�e���Q+��T��,���p�E�P.��J�`0,얄U�Aw���C�J�s�z1� ����u`�~Ի�D�>������b����bY���H09�N��,��`R�L����,��p:�N�Ds���G�����0�
j�CQ�0�����[�q@7qT���[��裤{�@��Cíؽ��e���a�I�[�{ӱ�����q��-@ >�p�������%�D�D���p�8X/w��sq ��x> uD\l;"�s<��w��Gj��-���F0��'j�n&35L�c�q_Z]^ĥfu �ke<@�
x�:!^�N�s��N��o0ꀸ �: ��c�����2~�@�����s�XSS��+6,�9|x���5{9��`�^���1<���c��0�"!��9!V�Y'�z7���^����6F,X�Xrb�@����|��{�Ԁ><:_�N9���f�N��;]�W>;cq~�8=�"G�<�?����$W|�^�X�H#��$2���^e��92�A�<�8A͑�2�ߑ�_l�L�	�%���͐Q9��J�I<o%.��}�`F�����V���@\��cx���9�*�P%)+�п���e)
$&���I׌O�ccE�0�/0�q�wYݠ4�����E�K�ޯ�dn$�}^ A�]}`�ȍj�w<AO�����dX�a3GFt89�0�d�M!�;���̱�[0DH��8ǆ�l��,�c�Ýo0No��c!0sd8�}X$nsdx������̑�tɸ��m�x�$qh�#Sr�	s����̐����tI|3��p��;C��4�&��}�$n�sd���䓸<η�[0���cF�2���`6+�����e>����>כ�V��AO����%Ck<8C��L��ݢ��n�nQ�v�M,27(J;�w9��Ea��i℺[��x"]o�Xbp�4y�RP�ۘ#�[�-�ݢ6Ό�p�ܢ8�N��I��6���OI�G%�V�p��-j?̎"�Ƿ�1�Ÿ��I9�6��q�� 3l8~���+�#���g����������m>����9���ҽ����0��Ο���?��O��)�>����p4��.�����|3�o���ο]&��3�\�}���������xz^q�V̿]VSϗS_�S���\�`�s0xf�\��9<s�g�]�g����ӷr��^�����^���	�\�����\�����^��y?{�g�]�g������T�9��C�
o��2��Oj�Z^O���쬝﬽�]��˘fa���9��o�^�����?]�hNE�2�Y��nj�O]�D��D]�D��D_���I����~�T=��O�O��>�D�֝m�VgeUE��m��w]�+j�P��0���ߞ�t�?����_'��!x����W/�k��ï~������婋.��ϟ>?�<}�H�����*��d�!�te^҈�"���fU)e	S[
]e�/l�5��tC^ݻ��kZ����_��ͩ�O~����P�N�}��~�<=7��$I��}P�{�!�q��}Y����A�����{a���cǇܕ��C���04{i�8�Q���@�؇�n����K�(�B��I�����^��O���{�|��zP��csk��	mk�8z��D�����v�Z�_�8Y8�#I�Y�E���Ժr����R��jޓ�H+s���7?o�xw���������8ej���������O������Շ/��ͯ3��"����':!w���?~��o>�7��𹣏�����T�^����/O�-��>ڗ���_��y���=����W\~�s��������i$��Aِ�Ņ���;���)���x~-i���"Su]Fd���W��Ս�16 PI1�7����b�q��?�~�7RJBJ%1��TIb��G�+|����m"C�J���G��({b1��N�����IC���3��8x�>py�4E
Mi�����s�(�dpO�1���'���?�<�՜\�
}�(�n.
\���bG�SM�x�{ҽK��7:#�Bg���n�붝.�4]�AF�.Lf����V�E��s��C�ő�HbRg�Q�//�%T�K��s!����x!誉ds�����n
[<(S��N�h����y��kB��:#Q����mV�]��m�٢�]�g�E��YӤMHrT�(�ȍ;��w�`�E<,���R8�v&d�.�[�-�P�*�*W�nC�f,��C&��&�):���?�r�`�>�`z~	��p��o�
��S!��7�mZ�7k��9Б|C8ڴ���ɢ�����\�YԦ�����\4"(*R�p�I�Q������K�����|���o�����Y��Kx��|��Fu�|���t�S+�4���Sa�O��U��t��Қ�e�^��U����˟�f?���{|���*�^�=�7�3v�ܕ�^��I��tq�:g�N�d�	1$�g�����]�;�9L?��G�
�ΧT�B�s/�2S>~�}Ћ�w�����'X�2P$*��ʮ�=��,�ܟ�K3ZJe��+���"���$2{�(+���F�N�j&M"����Ǣ�!\'"���ZhV�忥fJM��������gvl�f�YX@n����i�Bp>�������u!�Y(+���p�ef�*"K9�,[n�~�2��R���d}����>�y�6��3�L�Q�?hbD�G�����BI��bX	}�TՓ n�6�cG�X�If0&:i�������,���ycI��[3�MRu"��P�.*��/�I������럈,+�(uw=�v��1�������$u(���Q��/� y�~~L0�����*�=�gR�]<ϧ�?jg��v:S����)���Ѥ�h���~�B�����pdζ�2DS�$d�By�J���Al� v�,�y,������Fw$�.���o�bƽ���b��Sp�����F2�Μ��g�`��uZ��	*�"�/3�5t��e �G>Q}���d��2A�T ���9�]
�N��.x{�u���P�2:�_1s�93��2�/�2�VgZuV��Y�ٝ���A�u�;��e������5����}p�����H��ɷ���\$��yA+�I�7�˴7U޵�m������ � �����S9��:?�U��^Jp��.�
�@�[���tq��>��#�R�L��D^?}rD0v,�Ç��!U��H�.��q�%�@Ȼ��m|m+b
�TL��jb�!F}�Z�<Ӝ�L����F��{~�Ïs&���$�Nu��v'1��襑�ʉh%��D�2���]�/|:�uy�9K�#�t�bҪ�th��c:�<�Fm��x5M�J��fZv�����R	�)�w��C�_�਒��$hjuVcF7�n�<��Q�%ᯨ��W��U��'jq3��r5��):�����b@�>�'��F�2�%��k3���h�]��4%��J<���=�Jt�C��R-����$}����2�(�#�҅�����HװfF�PFI�ii�!�<��֓|>���Oީ/ߊ7+\P;�/��cXf���X��W�ם6v*\f���<��/K�\j�4˥vK3��7�׏Ks^��Į�������[��K%_(� (��WR=\C��?�K��+�_�����F���I�D���$��H�W$��UYW:����?T���+_��t]7�y(�.����y�>�G��	k���9sxu�f◇��|��W��vֽ��S�BǛ)�%&\d<�R���P����p�O��_����M��xe��7�R��3ᡠ-	gَ��5����j�)T�3�-]�U^O��}cl��f��P�M�ʴ��Yf� bϏ5��&B^�$�D�Ic�/�t5M�ƫY��I>���'�3�F�a���TW=��h)SxF�"��hu&du_�м��g��>M�����*����iVY�g�ϕ�j��vn�A�"�.�S��0��۔���s������'C�ҷ�d�vS���i=cBo�mu�y�	��|���DS�����{�`��-i9ט����{ͬ>�f���%n�U�˿v��N(��!�O_�}�*C�i�*AD��Et���g"<D�`*'=���>�!&����PxR��Z�6�O\�A���C�<ņ>_�g|���*и��K�s\��C��=�*P��?���ӏ��ǰ��g&n�˗�����~��ݯ����U��m�`9B�޻��?��{�GҔ׍'	���_&�mGw��\�)�siB�f�1(�2bSnp��'qh����Y��,H����ȳuԖ�c�/rS���\ty�i�e��*'���$R��X[�4��C�E)O���u�VЕ\ÉɄӗ��	������c�ι��$�旇r�2d�)��
�S�����IYu��+��.����A��J�cd������$C^�_�(�v���҂�;�6g Q�-
e�r������Q�ʸchF������>�.�3d�:���F?��Q	M��`^%x��I��J_�x䯣چ�RGZ"%ۛ.��wYa�N��$ ??JH�~H%=��]��Oq��L|�VSc(}A��1x�ӗ��D��$1������'\�/�rlnC$�?=�/?ʅ�ͧ��~�+�~K�<�7v�-�����5�A�B"Ϗ]���(��>w//���Oݟ�'1��o��{����������_�v�����I���_~��������ׇ�����PP.�a���O�K���������Ǘ�V/?c���￿�A���?�n0|��������Uo����~��y��k��~o+�y����Q���j�����/D�cRT6'1$E,}>D�X�w�������mf0˔8i52s~mU�mfL
&�DX]�4v������Ƙ�_��I��/7+��m6��|+L��8v����"�����?�х�KG�#��Z�3~�H�f˔q��R��,W�ʀQ(cv;)c�r�8��*��/�Y�/����`�P@@X�L$�����5D$����Z�Xt�aq7���2)g���L/�.�,�ٷECXU������5���}���)��k����6�n�{Q��ޗ�
�j�4S9CE���G�c���v�Ub�ދ*w`�7��vj&�-S�ݷE�Xm�w�8v�J�!\�ʸe��^o��T��������������kz�oS�Ê�������F�ئ���loڍmz�-����U���e����ݷEEX�������u���C���7.�a�ߏg�����-ϯk�g����;�+��mPMo��v���m8v;�mv	���xC�v��S��z���ǎUKr��qz�EnI��$b=��f��5s�r�q��,z("/Q��"�B�<%R��ޕ��0��ǎx��9k��۞��@%�v�@��1;���x�r��1��C[���O`�u�_j�Lh��E�SJֺLgH-Z�qKe�N�6�����b��6S�g�Tџ��8�m�>)��t���[*��)`�w~ڌ��>�f��c:���.���v�A�O��|���n��6~!cU�q)WN�+�iFj��e͚}[4y>�~P�ihv�44$	���f�����1Im↩mv�Km#�L��W��4é�!�aB����ލ*w`�7��<pYל{��}cT�x>�U�ؽ+UE+cA��1�A<�R+�8������ڤ+���z/b�<�ލY����F�ӫlg�3�,�@҅2-U��mj��i�����䘡m��2��oB`�utd#�~N�MG�Y[��t��k���F��Z��Td _�I��-��(�>0X+.̢��?eQ��Q{��uS�j�'���&!]��fq�R$ M�)������u�fp��-���Jz�t���O������b�ï[�]|�f�\&K?��5+�f��!
lK9cv�Y;���M,�a�( SVr��SQ�@o�� �7�'$:��8��L�3i9�nh;ø��,m�����i60�0H?LN��K��vӥø��&N���6c-��4lg?���
���%�#)]b^Ӑ�59]�n�;��M���fv�@�q" ��Y�t��F	�<�,�<V�.]'ڨ�uF���i]����Q��󈣖���J?��:���>�5K��@�-0�Rn�؁��8v;�<����i������3�̥�������cRRek��sj����n�a�'�x�V���>��4���q���Ԃv
�1�m��������3u�c��Ie�7B䤝_N%9�M6s����;H���JH	�]��"���퍝�]L��Oo����J��Њ����Ҫ{B8w��x��	�x�{c�c�q�{jg�2�0QI�f�v�H9���#n5��3(#EYw�j8j������ceƻΥ�/�i6Ϝ��cA���c��~w���c]��N�%�~0e�f\����0�V,t�ƶֵtߨ��k]���
�ˮ(�U�I�`Awv�Y�$��6m�l�ד� `���(�v�!x��Tƒ�i�SK�c�?�E�	�f˦W=~WE�qI2NU~W�%�� ]Ӫ���{�hj ��n'���?ח��i�e������1)v��p3o���PK�i��8֌�-'�޼Y�k
��:�;L�;PK�`�2��n��������K �}�ā���#��rr�K ����u����@�n�%wj�X�U��iU FԜ��V�,|'�0�OYhv�LI i Gn��G-CHb�_>�XA�����F9җ��ݪ:%h5*��r(�QC�&8v�ꔌ��9Ĵ2iU0U��hv���	)#u����q�%d�I�&�q�e�W6.����"W��μY�
�H�c̊�Ύ���������ݏ�����f��H��q`3�1��? q@U1���;ԓ��"��ԓ��b�H��B�rY�\�h6�?�ծIrBVX`fk�����h*���Z�f����S��M��^Gf�@o�SB�9H��q��z�!��b�.�eKM]s����hߗ���8lk��S�T>/�0�C�rUzǴJ@CP�L�HMB;P{W
��tc�2���Yf���f�-+�S� ����3��|ȧ�R'8�����]V�P����`3�Rc�y�5�{L"�S�!��,V�w`��Ō���i3&5��PE��r�Mݔ�f��8�	��wI�:�8m�5w[ہZ*/�+�Z��+�q��J��,�_�G��݌%�q=3��aRU�I*;��0~��K@���S����;PKe-����ǔ��CY�X݃ء+�U��ܤ~؎��������y���<TB3u��>TZ;uq%�؇ܔ>?'�R�T�,���$Jl7w?5�l����.wh�h�0�O;�Hw�����z"،'R0�LE��B9�����Z
X;��~߱4^��p�컿�'��t���W�k��Ҝ�ހ�z4�!�@��������C���lc&�O�f��[yH%��zцQKe!�jϧR���Sl�r&���h�Le��!��&EB�[S'�����	8��'1cL��"���xL_�����n��-N�V���6U���+��RJ���ּ����!�fiZ�i֌��:��ML�Y3��M���as�􄙇�}7�L����Z��M�t߱w%����=��*x]��i�.n�'͸�㌕`3���Ǽ�$�?~����>|�M���K��T}�|�]$���O��k��������O?��K���8��r���PK   �cW�����8 �I /   images/13784fae-2b69-4ff3-9746-a43cbc14e23a.png���7����D�D��D��	�k�{�u�!D�-z�h���3��� �`�2�6��w���'\�~�΃s�s�{���k�=U�GL����(�Ք������H����/���!qQR�SWR����rtqw��*������#|MDN���N�X�M���#*�(j���d��z-r�
�Տ#�,��!@P)�zO���\N������-rI���"����{�ȥw���
���j�St����?����-��KV�� �O�w?�Prd��:��z;y?�f/}�!�4&"�%%i,�%'_5cdx��9`H'(x�&(�.�J���h���c�����Y9>'�d{kꮞ���d$,�x H!';	�ї�}Գ"�`�Q��l�h�h�hF��yyU�=<|<<ueE� �#�S��I�z���uut����C��<����ԋ'�{�@#b��Z�p��Qq����B�s���\�UhW����+1���s�����G\�DE`/k''sB'�Bέp-F;���������?������?�?�DW�{�H����?q�Q���E�������@z�"��iuu~�Ԕqf��!�G�C�f�¨��"G�*ٍ�@  d&
��� ��:V^^���5�c���$d)��4���Ǯ���(�Kuh�ּ��s�1�l����}���l�^GM��X�媄v��� w�u����A��c�W6IB�`l�
����됭����@��!D���C��_�� ʹ w����heeX�16.Kd�`���ް���p�����Y����/\�l���D���oR-�v�����n�UO���*��X�#vܭ�(� \ɥ�b��X_�/�ǃ��ސ����wm�'��
%�� Pc�kD��K�Z8�L�{�xK���TA�Yhy8Eq}qSr�vX�Ⱥ&}y���M<���o�����=����$�V����@08���Jw�a�-g)D�Ep� �J$e{|������к�yբ� /;�M'�@�ATx�$��J�Ww�(���:X��T����+ޑr��xa-R��4t^#s������F�ӆ���>%}�mMkP�p�|w}�ݟ�ӯ�|H���U"�
��iQPa(����sQlvaW�u�� #���U��11�iDêۊy����L�]����ς�w�j���U;���:{�U�nA. ED�@7�쓌���?�NR#]�=�_����-bKB��WD�2���2�-�Sx��ۻ�*Ȯ {�1�k�nHׇ��W�v9
o�f61�聙K��e �bn�nvxX=�æ|Uy\���_�MҭH@ DD�3byx�O�hBT���C#{U�S|����̋����f��ZL������{ҋ�s�DE���������:U�"X����04��M`.i�Z��|�_Sb{A/��i\{8s��QM��:åCJ��T��I���x~�2(��l�E��'E��������ದ:�4U�y���ޱ#����BK���1��1�,{%�?H�k�#;�b���p�	g��x~A�T񢡓Z����ݹȻI� m^�lsa\[�-ιN@ԩx�{Qƀ.>X5��_2sⓟ���MU�6޼���c ���e?�	��z��O�g$����f^�s�C��R~��28E����B�����=��;Lt�G�>��M�l��;�uI`0B�����/�W�~S���$�)���5X>�����!J�%d��]��K��!��ՈV82=`�ז� �\�^UѪl���ۻfw��wtd'�2&�R㐽�1Z��3v��U���
@�n���]p���>�������j�&���F����Ǧ���O�>�������TJD˯�[�6*)�O���'QV֍�27�д�)QR(������݀-��8�s�1s؉Xq�9	�j9 ���#�ww�b�8�	�_l"؞�4.�~��d���Zt�X�����:�&�����Q?�>b�u�bV#`8kl��KR�q���Z|�֒~���f��=������!�3�'-�ӡC)��D<jo�����ǵ�0�������[Ug��7�;|��w��L����c�a�dd�܏E܇{9�9�Y��}B��7fF�z�YY�O�y��Ԟл���U)d`��O=L�:��Y��b���G�L��xN�K�������)������ӹ5�n��V����30�i�����2����J�%�J�Y$�rjq����z����ɳm����9ttt�}��x�i/x��KE֣{aR����3���r���h�*Xު�M��&uE@�V�iD\�HѾ.�܁Qfc}��.��O`)k����n�I-t��p@�pE�xW��)�Y|[X����ѭ,�ꔨk0߷�>$$t8���	�����m:����Ί��IA��?�"��3��h��ٶ�&�^-��k�����AS^�s{�������]�9H{����s��gӅ~�����W��[
�[Z��[I��;�h����#�]�m�Ϗ�Ԙ$v���Cs�T�^��gh��-��͟�R%�$��&	���i3�9�d��_l�:GH��6���Ȁw7���ݯ3���˷ĝ�����+p³�⫿&���S@Ѝ�H����M��$yЏ���v�1�����wM 0X��j��ʁk2�y�t�����D���	����h[�b?W�n�QNPZ�2�c���L�L]�R[8ͦW��Fd�4���6��^t"�xt��[ݘ���~��1�*���7C4�N�e����Vx�n��4{�ܩ���*�Q�(#�Θ� �t�߯k�z7��c:p�v|���u�e�ӛ3����˲^���
Q��AW�e�@~
"��	��Q�Y^����m�ER�Q�S�(������.������[�ыO=���7]H��吊�I�n��y��a6+��J�lٺ;�eZpCfS���X\NR2dg������P�B�Lh��㪫֚���R>}68�����#��~�t�U飘���.��0,VV�%�o��5�X��6ʂ�t���yd:w��s`����v�^r\�`��VQ�ƴJP��;�_`s�X���fyF����ׂ��6���C�Km��:�����۷���}�#����ǒ��G�YM����r^�<�I<&�oþn���4Y▏��r�|�����l~�\��"[Ĥ���.>0F��I�έ��p[�j=|Jl�l���g^��j�"�-+�Tm�Ŷ
�� ������TQr�e�����kH�+�-�[�����=A������H���g%s\q����8���[����\�v����Wx_��C0F���(���_U~QKQz�|S$&f���N����ܥY�5�ǻ����Ԍm���f#7���t�����K�����~�&�
^�]���ZY� /ɀ����
V�h��B:bguj��L�A�>���Ƀ&���_�ߍ�)U=�11���Z��%���)K`����I'g۹�w�]/���V2� ��
,�v3L|�d�G{U�S�p��8�����U9ܹ�9�Q)㌪��D�R�L��@b90�"ڹ�(�GV�y�_x�l�۹k�#(���8�㵃3��W�l�P���MS�^��7�<D����ijsz^o�L,��!����>�L�kh��S�x�0�2ROE���V��l���@�%�%��G~s%q�D����p���1�قD�t�V��(3�ɛ��_�<e����!7e�I�Sq�=�c��K����`)����d�g����҉��g8f+��Y�LqLK��%�))���U��� �"���[=?m���q������e��a씏ceמ��8V���T7�Y����#��?�3>NX�>��l���D�$qg�S���Ͱ�R`xܣ	�Ds����A���-�E�7j=�h,�����U׉*ї�C�]k�	���U88�gtz%ojZ��GY�U>\:2H,2�0�y:�+���H�`�������)Y����Ta��3af��	��%��������kau�<u7��K��R�`�,��94�8��xD�p�\6�-�۠��2�l����f��p���n�B��šE����e��Ĳ���&D�p��w�Ȫ&#A���t�p���p( :t�x�M���������¨�t�g1!H��f ��v4&�0��:pE����:Gi��[i��2��Kխ+T%o�6��ʒwm��t�~m~;*�ټy3�QY;���O��Ή%ڤDl-S�|BT#��c�SV=�&Ͻ��H D��������Q	�B{�+k�Kă����M�G��SP4�Y��+�U���Y�dj���hRR��� ����՝0}�����P�
m�����eP���DC~k�WPv�|��Hϓ��]G�/�@�%�ȯj��q��?�EO�,nv�j��K���㮈��#w-r�o����q=,�P����������Tf��eI�-
����;R��6�F�ƙ�޶�,�����\`�����	�s#��%F>��j���
�ඞdٻ�e�w�m������5q�{T!�" �X�����s�v�*tc��6b�m<{0���/����1X�y�_f|�7�Z���:�&S���*g$���_<rCe���n]PQV���VfT����'7ݫO�{mݭ^�g˪�y� CEіӣ�-�J�WU�)��� �ŎQ�Vw���c�q��c��F���#,̝Gs���F��#���tQ�P��GW1��"�`��9(�3Yq���2n���u	���]�� .zto8JΝ������O������=J������^ƒ�ÏW�7l�F�٫jT�H1U�[������Zu建��~T���V �݋H	�WbX�B�شa=^R�˙{βj�y�KE�]�pi�����{XC�S�V_T1n.���#~o�$հ؅D"��q��u�$)I�).NVM��fV�Ds���r%6��q�✧i|��Dkgn�Ov�%�r����zx������$�O�<<2��q7��`1������:剹C��J�LC�b�b2��]���:�1	��"���7���u����ɐ��Z�9���
=W➖dvK����0��x�Xrr�p�c����Sǲ�qYYH�7��p�
����5�n��3:m�Uh"�S�T��h��C�M3I7�9r��,�`�Z�UNEҹH�1�]��������K�_UPB5՚w��n||�Vڷ���e�?u�hXᆮE������P:�Ϗ�%���d۾%��
��,u4��$_W)0�O`�u}�G��p}��$��s��Q��T���x�X8�/Ç囖&��?�����׭�N�4Yb4�K�q	�N�"M(=&�����E���ݶ������WT�����E���؊��A�I����L	nB-�)�~����Fx���Z)0m���R�؊i��K�zc-�6�>�~f@�5zHՅ���Te��0�ٸr<���^��^Qq>
�N=��h�զ�ǉ�p)!��z�(@NI~��Q���Ru��t�Z۬l��}&:�P�a�7<d+�t� �Q�E��Z�A��SX�un[j��6B?�"�'"��s��:sw�������0�w��I)����������,�	�wD7U�||!\��I�'}%���g{0���}-(��MDH������������t��I�$�e�á A `_׭�,��=������UT䠑��͙m��+6r� #��*�0�t(�=|�.`���$�:< �>n�3*r]�.�?
˓���u=�@<�1�bd�ʿ���D�L:��6�́�*��d;�<h{�=��]~w?���]��l�w��34���X2���(���f��W{�@&CY-p���b�`A���*��_񚬟�_�>��g�VG�	ӓk-�i��c���eG�ꠙ�9�!��2���N�
yR�z����?'��>�̹_��po���נ��]]�㼭Ǎ��8�
�H�9��� �8 ?�uL��`�>�,��,VQyMt�a�����kx�i��ql������*����@��̄���a�x����݈����C �M����.$4��K#[,���|������U�(���2�}��r`�F��(Μ�n�3��y�\7Wo��5��mv-w�)!�Qk�R�5�G�ݚ�����@59�+�r�������=��C�LN߇C%xjʅ�8�)�?�M�Gǲ�G$���Q���:��,�*+�q�I��iC��[;?�z.�K�?\"������d��n{�o���m��q��8ŠW�0$��P�����Z�*|M-SW�����9�?D�/$��V>g�G��9���J��0/}���,�9��ϠS����b��Z�mH��}2��Cz�Y��?�G��U^p���e��3�[���=36<7��?���K���c0/�F�5-�V�$��ԙ�r�(7��;"��;�G��N�s�`�2<v�A�o�޶fWm����Ѿ>�#��qsj]�������ě��׏��[SL͹2)~�nEGg�7��s��
\��0)z�S�R;j!��A<Y��!��4�X���B";�n���](x�m<9�/<J�>J]�����.,"���&�Zm��/�%2���EG�K�W�$���9!�"4ز��
vѷ�Ȥ��|%$�����n��)藧�vM��<�#t�Q[.��V�]M��˳J��>5��O[0�~_�*��o���M�=�m���/��n���h���\�J:��~P��PԟtS��B=](�$.��+<~.�>>0��Ì���r
ڃg[�L��34�:��У��e����4|�]�!���~��Nxd�%���L�G-O�O
x�=Wgɥ�M��s���a?+ʈ���ĺv�&�!{A�=�,-�+煮B���	���Ŷݯ�_wc'+�o��R�~�fݒA�$���� �����/z���d�[ЃXh��0BL	m��H�hk��|��w�];23Cn�@�P��o"�:)�:!��,��`���V8<��P�'?;�y��<88�d_
�%��W�o��[M!.�qS�Ǣ0J�����to��4�	�2I8��<)kY���+B
�%6�3fk�w�WO.�_��p��߯�;c�_Xל�r����ʪ3������Z�çw�`超>";��6j�ʵ34�F�si"0��nAA�+���v���ʜh���\��>����Ϥ4����^�\�~K��y��``��p�������PƋ���btt����l�E��r�,嗝 ��i{/���R�ԃ��O
Mp�I��5�y޳'�#T)�"g�n�uv�5�)��a��C�?7�Ƌm�y̄�'�T`E ��H���w GlX��슩f[}�桦�4�dڷ"����&ߙ�E�C���DB�ښ�+A�_��V��AD�VR�� x���Q�Fs?����$��*:�
��z��s�Z{�E��Xu4���� <u�&W5�!�g�GӴdd~�nۇTlK����}ź�,�.gҙloyV�lr:��Y�Q�h�ά�ö�x�G7x{ ^V���9�����#'(�ތ����J*a��\��C�>)"����X}��h�b~:��������*�Ֆ�	pfh}�`��Ώ�ˠ�1X��v�A�n��*���N�a����>����[%睽��4�*Q�;��y����=�1��yDس
�$0񩛠��VEIzI$,���$���C�MIVv���G��Sw����&/���Fܕ��/��'��3�͗$k�Qȱ7���aO����s´��P��t_��K��fu���E5k��-�sKu��dX��t���)���f|_��V��$��ۣ˱�og�uՊÌ��V�{�k7G�va��E�w����篘!ѐo%�)��0�8������x���m\�%�)�b2]�{�%t���������{�������l��ߍ��6N������Ko���������\����v0���K�;��2�<���ߜf@-�2����u)�XT��{�*�}��k1���b���#��73<l��i�t�{B�Ɗ��B_�HJɀ����NE:vs�Cr>S��bYS�_1��2����Rƛ$w�2VL�2��G����>�к��.:�s1�����x9k���%�#�S�Y�� ���GG�s�dQ��ȣPT�:%�LYL{oɎI��U��1�yTZ�@�Atc3�G�-��9E�Zw����Kd�wkJ���UY��4F�O]sK�ר�ef���ο�-���-�%p�RY�얮��Mu��\�\lJ��p����P�bhFh����cK-d׌�6������+=�e*ߑ꿣��֚_�����v 4&�����|�5�{��'P�7���E�@@k��d����߳F�	/aӋ�Z�%�a�,�<��_rF���;��������
v:��.��f<l!#T�N�(�M�T�Z��f�q 
���e쳠�c��h8q��p;����"�����s��`�*R�'_�s���?JP�x���d������[\
@�$�����4E=�M- ��9������kU�]�M�V��
��v�@��Gu#^�b����]���|
��>}��af?���
��g��"^=֨:|4�kY[@]@ǭ����<ld��HPz�ό��zh�b����+�[;�?� M��gm�`񇸸)�S���DL]z��f�����x��x��U#��R����R�j?�2�3�8����h��4��Hn���<����^��Ͳ�P�p3�.�޴�X���3kA&��FdD����2�P3_T���R�E�<����/q��<��O�n|�%cwc�DQ)4�`�O��i'Q�ҦTX6���^\�3�;
&�B��47Gy�n��^3A�	��*��)��ݦ�o�x���&g���.��3���y��}^��R�33�0���aŔ��7�ݶ������r8�R5�jױD�6��X���je�W�y+�2��b(+l,��~/�!��!�&�)����oB`��[�g��Ȁv�M"U |�%����șX�$���~�}������6��lB�b{��Ŗ��Z~�0���}��ު��U��	Ct�w�z$ c��e'���*��B�n{R�z�R�]���I]-�"�j�7�S�#�BNt��H_`>�A6�8yR���8���t��;9X9h��+�|�q�/�4u�M��~��mf�ȣtF���k>�>�,�LeM���_���灶%/�� �����(O�
�tqS��5�R��$�>��n�c4<��N�����O���G�Ց��e�-�Ԣ7���E��������F��7hvu�o*L���(9ϖ�\F����{�e[Ϝ
�N�C�{{j�T���-)1_)�ٲ�j���n�߽[��G�@h���(���,�t�Z��������������ce��q��8�	�S�z�**k� @��Eg�"��-��/澝nRw:�-$zr$s3��ӓ���ύ�.Pz��Z��爫�R��o��l;�R@ݿ��:[
�d=�z *��`Rm02m��	Z%w�����T�paw��m�h}Gر>7����ۋ8�h�/N���J��"�g?ُW�x�_oQ�ݨ���@�o=����~V��l���6��QB�nZZ�ku���ab Z�^{�t_@�*��Cy�>ޏ�k��Y:�+g����M��f��,ox�h��c�?��	�O�����|B����II��q������OH�ꑲ�_����ǹY)�F��CD����aGt闅� ��*3c�������o�-�DA�>���.c-�$VD��Ry���
��[ټY.��Z�^�Ye������{�b��B*V6�*K-?:���C�먟sq�>���̺v�l�ev5��M��g��裃wT;�GH�(�5/���TV߀2~�A��J%/��Um�(!h����XY^
�n'ܦ8V�D�t�N��4V���e����O���_RF���G�_aj%g�	#�fs�V�pψ���_MV}�F�3��?Z.��g�4�?|5j�,Ș�Q���'�;*Ry�[1v������v;�}L�f�[3�B�K%�GSt�~X�K+1��6N��:#J�KT�������(sUF�3���F��� ��y�qO<}D#-bF�Υg$/�³K��9�v�#;Y�����?èF3�u�~'�r;ו;}N9��� P ����T9��{�*�yF�[�2�9��+Hw��k�V8�p��QXd�m�^sIv
�4�����_�|f橅!W�-�;1�@�X4����Ʒ�"���"��<�]"T��/�ßM�T�}�"*���:Tώ���.S#m� �zt��e,S���*��vX>wL��{�iכ�f"Gh��V�PCEGl����3#�Q��[��^��~T��c�6�x��i�֩z����PYy��D��3���A%�(J���?�V�˖% �a�}S롁;jX�M��;e0N#�L��`gKQ�@�����!#�W�:�і�Nl�[~�8�M��x���ϝ4	8�{�:]��rsڿW�v�R�.�,s- ��5�%�&
�ssZW�u�
w�_-f�� _J����'-̠��T���A�o@��'O���kS6E�%�ȗ�2�=6Ui�kW$:��% ����L�o
,A|^]��,������C2-�<�T�k��dV{Yd��Ɣ��u�go�&Ӓׇ�_���4��`��.�LJ���i~�*n�[�����t� @�Re���?��wݸ*��i�T-��ws"9�9]h?Y�L��-��C7�	/:��[�����sw:WO��u�vt����p��T�ѻ`��g0y�����b�Ƚ���ȩ�dU(�{vX��h�#���(z$��0ןe�9�Ӵ^�t�D�����}}�<�֚=(��/���I�����Ȇ*��	�&ٻ�F�:O�o��\��Yq��Mܨ��>0-��:�N�a�9t���%{9�U�0�W��O�bsV?YU��Y�j��HA�"��}檂�^��4�
q��QBF�m��&	�͕,�Q�.�#`�����J���2�O�̧~�-��ȁ��T=��5���W$�D�ب��A�`~7�8���5�\gd�X��%�����<(��=*a��y�P�
+�)c19�c��J�WN'	1	A�fj��[E���u�Qn�>w�;fS��n�$��Q�坧�'=��z��ք/`������%[~��}�:q)�r�D��Z��6�N�XR��tPw�G���3:�m��d.h.��g��
���2��!OR(cf�uw�*��\���c��1��d:)�Z�a� ���W<1_��9f�*(��q�J�<���/�/�W��$�$��yZ���ο1e'���Z��6;%�2#q:���:�n�ɂ\�`p	Cn7������,����ãl�JO�2��=���łF�m�{D�T?^Q=�*�Z���!Y����rD�w;0J�<��<G��pYaR#�{qq7�G�7��~�o�w6p��5mËb�q�1�0��a+�zI�Yv������LGE���P�{ySԳ~����j��Y���j�K�f���-��=��U�(Dt(�^ߞb������i0���uk���ڴƩC�v���H�Mᅗ'4}?�x�u9V�;W.ʟ���`��Ӈ����"�a���K���8��X��v!���Z�eۿ]b��^?�"�	 ��B�^�̅�Ҧ�ž뚈3uq�}Yj ��J �!�Ȏ�Eg f�.�w���<H߰2��	���P�h����YJ=qx]ӂ��m�ڂv�4��+ڪTIU	6`����&[�T���u�ؕt1n�ě{f����5�No����Fc������A�i�ݧ �'��j��^�9���9I�+ƝR}v�4Bb/%@�^�!���f�KK� ����Ft�c��"y������D�>}���Z"�����Fv�V���JO��F��������44����W�F=���	��-�X g�e�<�$E�o�7��y�m�<Ga5��!�vz���wL C1XM����n�Fc�o�KZxѣ[�y6k�-P31g��r�}d�ek��r�#�5X�i$)���EuTW��nMZ���$�}�L�{��W��DD~�PP���r�!7���/*����L���0�!���M7�%ѥ���O�.콢��a,��ѬǛ���b��%����N�kx�5y����1n2��Z�w�>��İ?�b�C�8���i��,Xٖ�=������O	�H�*q5U�z�萌�-!��\��or2d���t+5��s��\H�.&R���ӆ����,&���M����l���NK������t;G�w���V�C������Wv�"#{_C��ֆ�f�G��n��X�陔�l8�����]��8�0�axE�,/ǁ�V��X��n�6�Zʨ��8F��\ �nW��������Wę�Bn�2$�r^$�e����j,ؒP\q%u[�#�q���*<&-������W��VVf�Ul�#.�m���"k���yR�Ѓ�݁@P��Z����#�}J7%�a"'�O-���[�X�a"5����}�F֑��c����1g�o� Β���N�Kըl�]]%�'�"���A�H��sr\!�f4Q�u �	���;�K�18�ݖs�����V7qΧ>�K#�r� � ���0���ag��y�cʖ��[��Ul��\Q�iP{��L�#x�xMv�= �e�F̘�R���O������ve#��mJ�.p3GMR�q�<4d�(��C�͂�<�Z������ t��<z�����������~��O�r����?����i�C�m'���j0}��A0��d�Ǚ8>��A$�Zͱ�@屰��4��n-F>�ޖ��%�(��2K �O����8�w\�MZ{��T�8��D�(�1�������6}$ ���=S�������Ji�+���8Լ)"LWv��U��l�"%��Sf,e�{me>�3�h�����M9Q�X�ȭ4�G�?�5l{���������S��_c��ԇ��H��|
zBl�Rc�x�q�Y���P��mE���1՜��*�4>;���4���iM|�MCIlz��D!Rz4��Fh/�/�����f�mʭ�/x�!�ȏ�w��zCt������E��]�̫��˞7��n?�A������V`Q����9Y���0�T���6H�}��K�=��8�6�����J��L�m��|z9�9Cj���{V�͓W��������\�z�X�tt�.�z_����
�R���k^̰�X��3$K^6�X�C���*ο�t��ʿ�*�:3��35_=p�Q�L H�ŗ�X�ҷE�ח����7&g�A"��A�-IΪ3�eB(��'�-����+�\0����� s��"���Z�ͣ�N7���s�Ǌ5]��(<�{��_���{欁��P0�O������J��^G6Ǚ?�ƥ��T���K����o�������I���W.�"!��P	b�2��zr�-I�f���8_�s�d��K���a�"�`�G�vM��͔�J� ��r:6M��*����̪�S9zuf�7;0�W�B�񹏭�žvD�ؒԄ�%ߛh��A(�R��=�-t�3[¥[1ڸ�����vb;ʌ|]:9-��K�n���"�1��[��� ?ѺDQ��h���\7%�����DČ*{��>�x6�3;��*�!6Bu�[ufZ�d�w��߮��7�m5��T��m����T������pܨ�5O��?K!�B�y�b 葽����x���4��@�V(����.LoK8Yl�p�Ö>	ƿ^/d�n�e�z�lD��b��=9��"���u ��74�Oa(F~}�66����nL��9D�� Y�4��g�}h$�����@��-+�e�x�P.���!��^��^�x��������=�A�U��{yX��ja5Y�w"�f+[�E�bu�}:�b��V��/%VY��\����^΂�;giq���ҕ\hΑͦPv����g������GG��?3čH��r�*��MS�٫����@�5��_n)RF?5H�t���t@$��5l��v���o�`'���]�yJ�C�19[�/-�;^�M�x`�C�l2Lwf�R+��eA$�͛�`Z�g��/|@}�����C���a���f�"�y3
�Tna�g�y�����؊���'��:6vվth�y����wH��ۗp�����dj^�m�XJ��BB�rF�:m�S���#�F{0}���q���<�a �/Gϐ�&��dA<�xA�����&�8�D�t�+���5�����ՙ�B�ON��'@s���v�O~��g�xEx�����]��w_�P{Gϑ9#W�i��w��؏�I}ø�I�%q&9��FL��𰝲��E�n�/�g�аPU\>n���6����[���W9��&��#6�����7����r�;�����e۬�}�@���\H��+�k�puW��4�!����i��ߗ���R+)Qf\<����,��Pa|�����@{՟c��k�t�oۈ��v���4b���G�ɣ�:S�L����V�����
���+���r^m*��&7r�zCc�	s?C[[0�a9��$��P��vE�l�6��]���k܄M�j7Ý���e��iKͺ�?R�B��̒�����j^�`�a�Q!���t`�����e��[����l�9�|�����KO����D|�r�><Oe*�j�4ry��B�h���������wm������m�Gͼ1a-���E-ñ0�������]ˎȴ�(�>Z��Z�5��]m�u���}��]��qh��|�k�?&]��g����(��孓��p�C�Mn�.�?���TYWq��&�r��g�
I[�r]~�G���ɽǷ��=u
�!F�0k5äL��#��<��*.Gq�"�2�1l��V�O �<sZs�*a��0����'�(+��Z��/�#6����7~Te��Y�#�N��S%�^ra���Q�N�i�nBL; �j��U~�)��ث�n2Ҵ�e�]����I�=��$2�|M�W�90n��xD�p�C�J4�L����"%h/���"�?p�u1�{����J�;��(���<e��ϒ�b�m(���S�7�XЪm�^��ur`<(���(T~T�֘vDp�I7��.A�hx�˖�p��X��ۢ�,�T3�Կ�������3����v�9��8��^�y��t��%r��/!���t�{]<;h�]j�Q�jo ��t�R�z�4��xlh�1_��36����ԗ�>���8��ATv=c�
呿P?ۊ�&���Z|M�S�9:KcY�o��|�!�ĿRņz��+s���d����Z���g�?M��7�@���b9���]��$�䑌�)���x�{��%>�$j[�f�Ϝt�7���X+W�O�m3�x"Q���9u�p�|�$<�������-a�'���D��~r��on�4.tʫi���JOBZ����-]�N�� �&D��^�9`)[�� HB�~����%7��n��V!*U@�������l�"yz�~?��*���}mE�
�̺a��8��f[ha�q�6�$Oi�d��A&��`�w,�v����.^�d���w�Л�o��"�n�dҼ�nf6�K�#R�pS�����r����S*�"�@�Հ�4�3���� `�7��$$���)@�|hl��J�:��uGa;����-���z6�n���{���;��	�g�*�'�c�b���	T��Z�S&�:�?d%Tlj�'�'�?�	���.n?��e7��H��HWLĳ%��6#��#�-i��#dʆ��|����Ky3���q�(!�,wb���["ۋn��ٗN=f8A�G��Ǉ����<��յ��?��;mf/�,ī��f�yD;J.NV�3P�Up���)�Z+	h��kE�x�K%-DЗ��.��ڥ|b�����Bc�4�Ҏ��:uiY=����n�\��tZ$�ʽ�4s<��k"8;r�&ة�k1��gX�KD�{�d�#�@b�hG싴�GiE3�C��b<�e��{��vbŃ3 ����6v�eU!�w��T��,�Q�J��_Dɋg�QJ�A�i%��n��Y����C�G�Ԏ 'Zb�7��_���Zl׍
�Gɦ`��oa("������v9�6?˔!���é�$#w�39!�#kǾݪ:a�)�B���{����(,�u�L�[aQ2�����+�҉=��|,�K�-r��@�򡼢�T�J��Ik��z�����խ�O�K���L���	��#F[J�yP!_u)�s���t��d북X����B�n_��%�����QG_㾺s�d�����x��^46�k�+o=��N������>^�,�5��.�s�wk�>��;Ъm����ܮo�w����a�m���܆���t��S�Կ�l4j��D�� �3��Z\Bw�q/� �q�j|
�J"KV��_�$��H)ND�sXkrc�r},��e$#�I���d�|����t��_�H���6F�~�ʆG���:��Ag̯J4��w{�갂R@X;��x�3k��Do�0�a�$rrwf���TG�$���pU�F:H�#.9�P�!c�o��C55�ź�A�=
yj�2R���	�á�lȒ�,
	��
���.�=N��&�a<r8�ƾ�-�D.E{�S��#���"gL����3{%���7���sYY~���U�ׁ�1q�!����־�H� �*�8��׼�3�@��f������1��N�Ző��a�J�s&����Aj?��nr��v;���dpV�������������?�2�i=d�/W�M��H����04ѓu�B։#_��9m��;Hl�6��=��;WΥ�6����CQ��Ork��ŵ�8>hk]\��t�� �"|�3������k��HL=��`,߫����@�=�&�!�*�������ԤA:s��@?<p�ZZ��b���V�Ps���8��k0�WY4���DqXca�Z)#�8e/}��~X�P,.�%ޤ5�:�Zdy?���iY Q<�#i��� �Hb��5_(�F.��Y��pJL�Q蕴�F%׋��۝��r){�NK[Y]B�g>���n[�:#���#���i��U�bOP?����6�0�ylQ:'��_���u��<�پ�IP������D� j��y#����A2#�!/+k+���v�}�^������F�H�ݥ���Y�Y����`q� ��h�a�R�G��ym��m�F;����ae����׬5Z��4֘Av=�i��j`p�ϰ�v�������>����r�¿�h��b���'e0�F��Ӟ�	�F{����![KD^���&��"T�)FD#8{�� ��]�Z΅���A1RU(�l+*�"O��/��C�p�-���I;���y�bwm��<!!���P�qX3�;�Z�+rOP�Fk�M��R$51�4��KSB;(k!���u���jzȲ#�hS�'�/�Lr�m����o��D���m:�PT�~� �{��d���'�*��b,�-��X׀d7������FMׁ�5��Q��:��IY��ނ�5	���} �LK�{���;�%�U3��RWd�}׿���{spO�K�����;�	�o�]��q�7{1���1��w�fSvI�^Ľw��Sn�_���i��3d��5e���âs�i��Ak�|�{H��'�p]3>�����B�6��p�zz��L��+d�S��V���`@�[�v�8��0��3�5�h�t#ǏN���0�c#=��#�*>׈�C`}�ѓ�2a��A��j���2{me1�ߺ��o�F�!�i�=<���D�:�q�bh�t|,���2-u�Ř�1����DH�k��"���<�G���*�H	�T.� �9�ٍC��A��{������Y���=(�Z�d:���>^gz�s��[i�܎����i(PD}l�:}�wX�d��DcoXsچ٤=��`�L���JD�A+��w"�gA��wR��l���V*�X�y�h�D;�L�*�0��)L�P�� ����������j��7��/��/�g�y&F;6�ܮt���P&�]~���|��X𖦙7�m�����|x�: ~��>�����U
����a��=�U�e��@2�|�
{������������޷�n�{a�Clo����l؇�ch�u�d�4�F�UcP1�\|� o������eh�!&���q�����B��en�`XC�m�uy�{�+�n��FT�Β�����q�S���8!@�v�2*�;�*X�$6F�zlL��(�u����*��樓#�b*�1JoB���V��1���3�Y�o#'1���Z,l���y��-r�U���:YÙsj�0U"�0k��;�ZD�*p�F��	�>J�UƯ��.eX�#�7��� 4�?�4O:rd:�H�7/P�9�F�)9���L�z���p�HW:}����E�Xt��N�9��kF�B��`�?V9��Q�,��&N�'��4����^�LC�v�*Ñ��_��/�O�3�O���q�Ȳ"@U	�tr�`�^�C����V��_1�U5GԩۗF�k��KvԽ��+U��s
-��v'@ bv�zM�GK@#�g�ڿ}�n��m]����7�Ҿ��,��}��5����6���Y22�
�[x�.�rU��L��}�H���?��_x?����dz���r�Y�=88N����u�������8�<m-i�jGP��G��4��D
�z��:R�(�.��zwѭ�歬X]^ A���K�S~���l���Ɏq D2#��Rr��6����u�{��a��68�6-�lo�]zPy�<Z����_���[�PP��.�~U����5���8[�f�H����oP/����T��1���H�`���Ƣ�L�	��$�\A}�Z�u�ǏF �C]x�L�yl�A>1bc��,:濓�����s��#�/R�.n{I!+#�@�^�M��6\K6�d��	/~e��*#q	=K���<y.M;K�Y��M�BpS3���p�BW����u�k�jinɮF1�e!�4��0[���bZv��Ĉ`�����hL5|*������ג���5��æIr�ݝ0�YI�gC]e6��ǉVZ}a=В.��BC��ȝ�l'�sP�K?hI������㭿Śb|rݭ�(r�O�v���|����a���}�V9��&���R�����"B���.?��]#5��ܽ�h�2��m#�p��W�飇L��Ž��_�������H@>Rm5��p�T���g+Zm�0����g=�=>��O���F�W�S���>F�F��
�����)֎e��z�)�xT��xy����Y�����Bʦ�����{���j)e�G��0�D��8{C��uf�����	�:k=q��*�D) �V"B�}�W�e����Eh\u:�:�|��(�H�.ryj���<�%\L�M���ӆ����Wn��M^���60r��M�Q:��Rѵ@�f$Ԓ
Y\�F�O}Li���2Dc������Bx~�SO<���s�k<�H������`44iGZհV9G�+y�4ٗ���5�^ƿ�s��X��$��'[9�k_}�=⇰<z����Ƒ#��̊J8a��P8f���Վ��my��|��S���,ci�4� �5�0�$�4����һL*m������A�ך{6��%�{�^�:�"�e������1�O��'�`%��0��;Ic���({k8ݴ���2K�g]�{M�,�M�6��*��s��w�kw+��R����mZ�A'��vr�1x@8-����Fv!:?|�h(T_�(&H#n'�1_]�w��Y��~P������&^�<GŰ����L_�����ݜ~=���k��Ȼ٫^��>��_#�����k�p�&�u�� ��� D*d�,��6�P�E�� �t�p��=�	�D�}1�ƙ�*I/�#��J(S�q��[�S2����IjQ1��9=���mfjU����ZH�G������%��V^ј�Ly�>�ܝ>	ѫO~��6NQ�c..�&j�9�����h��S32~�c���H�Qˆ��_T8�R����t�D��Q`l�\%��Ijɀ�6z�'?���ٓȏ�
�s�F�a��1�D+��`��.����$�iIl";B
=�cjl"�2=��G�$.�1"�'��={�p&�p�&���SO�5���B����5\���9��0�>d�Au�x.:\�U׏<�i����~�\?��zm5��]2.�f�'�]f?l2P��^�9�T����%���&7us^OQ�מ��%�{�n�жc�s�9�l�}��O�"�U-����p=��W�\50~[聳���7߾@�E	��ވS������aM�]3�
B[c�n�\��,����u��F�t��9:;6\�x�������BT���u�|�,)	ۦx�\����+d�4Kj9W�|�5t�9s�ph�%&z�no�� ��hF4B��W��j��(�ZON�3�7?:F�w��&cYޕ��]-�?�;�!Z��c֝�|�m�S�����-&I��g�A2�s}h��z����c���_�+�kv3���4�b�<(˄��r@�I9��#�W��-7���n��(,<s��6�x�v8rκ�#��Ní�57..��������aS�]Zc���4�t���^?G J�P�Bv]1��m.�Ѿ��P;�)�i�=�0�����މ�U�k��F#����A'���r�:KN$!7�]c�6��7��e����t-ZT�K�Z_���f'�Y�J��"]�`��rՀU�gʩ���6M�S��74*0_��D�T+���L(j�Ө��ʯiޣQEEL
C/l�F2��Q�@N�����g�>�R�r�	�k�MY0Pg���ց��y�|:�j�xs����9�dz��<��Us:2��� l����cL.�XGV�(Z&B|��~׮^O7��m�nȊV�7=����8��#���#�-]7�̲���my%,���p�����х%��2�Z�l�E����?#9=`�;"b#4�q[d�̓�%e�``�ճܷ����VX[cT�X(\I�N's-�{�$ʶ�@l�>E�����H�� KBS<Vd��'):��x�.[bۮ>��s���,@�����l�a�=#�pr6@��6��[+i�4�H��"tP�`뫊�\o#�L2j&X��v�R��5c������3��c����y�&�q��ƽ��������'���#fI�M$����ν[u1?`�U#g�Qi38�H�\ϠqV8�)�R/%\�a�_�t3֓���˷9��1(��fv�s�Mf��������4OՍ�|�+Y}h���a��>��H��q��ǆF��̵�@ i���Ƨ�� ]0�p?ѷ'@��3���w�d�$o��w���㘂h�"PQg�6��is���7��'�V�"�o_Xڏ;��=
��2%Cϰ����9z��6望�l���}�x� I�����M�0�5`,:�0����G�h("� �#R��W;���ª89�5��k���F�t�y���k�����v2�%i���c�#�E�Ion���o��F_*N�pސ�$6��GEi4�Pe�I�஀�U̹~���
�"|�"ցPA���F�eT��&��Nh�󭩰����<U1I���k����+G>l��1"�!�Ah��3T������#Ҝo�F)���5�׌|�xί���]��Y��L�)���1��?�vԻ�����?Fi�@��k�E�.dv�5���B`���n\� �� J�Z�ar�ݣ�D>���A��e��J?8w5����'�M����%IED�iinàg87�F�s�Yx!� ����e��\��f��Fᐽb�v��Qb��|t
�5P��o�萩��̅�;g��<d)��K��\
4�6��������t��a��{��`�9;�1�_�9j�
$`gTg��yYOSd'��pڤ<��d�S'���s�ɧ�I���/�skw��6B^z����uѵ�[il����Z�a۲"�&N\�~U2�p�2IN�F%7��D/e��a�2����Z|G��k��N�ߓ��� /�G��mz]ܽ�T�wpO)�l�s�S�%��6�.Q�#'�e�o�KYQ
֞OC�{R�<l��
@D�0��2������6tZ$�"����X!�ա�dTGG���G���i��0���ΜI_��g贇C��{湧�c�!�nl����? 	��1��L���p2n��%���7=�м?ԣ;9 	����pDM��F�a����5 v��أ�8H=�	GF����.�=x(#tTQ��F�H���Z�8Vmh>��`�s���E#�*aia�!��m�cg�^�i2?=^�aD���i6�qX���րE#:�Qz��� $��G':����˷�׿�z�ޤ��{�<���TV�(6��i�5��yT���}ˌ��f�gE�6�KXӃ7�}؃��R�/�g�pŶ��������S+�9�p-sӀ!
� �"���=�=f'��hH�C����rc�B��$��pf)����Y����`�O�v5��������)G�$�xd�IH������:μZ� C�C�}x�Q�mH]o��vz�̉�Eg���;���}i������IJK��s�E��������t����9������wQd��%?),��{�ҙ����}!�RZ4r"�`�d8|jլ��î�ʩQ���e���>ؾ�T3Q.fT�� �`��9s�V?D�,��yP!�pv������]cɚΕ�fT����0����͙R���&g���wlߥ��%�c��^����l�Me��t���6����:���0L�������%�y����AŪ4S�Ϣh�N���W��J ]GN�f��.�������q!�m�[6E;pH��pga��	� �v{��!j�m�*Q�J�����l�:�$����G��%�e�D@B�6V�*��u(���rt��2��P�9�E�s{�����
l���B��׸�<�ΐ2tB��``����Th�OV7��5�#Z祃{'�E�%ŷ��$�h�5�N^��#@��.I����I�q6"�E[lo�z��	�n�Y��H���/s.�t��&i�������~k{�{�EE�,�vg�3�z�å��*bwY�et�@S<��R���hx��
D=�s;L`-�LqP���ٗI'4�U����#�|���Ci��*5��욮ctZ�RpS�u;m���X�h��U<MH`Dæ�lbЈno,K�4�(�!��/>h�牑\[��l���H���'{�����l�2#VPEW(^7�[0ZϾ�*;�"@�
U70�ۢ�ݑ�1fP�i.�����L���eC��)7ZW��x�x��Ml�4���AT�Yo�c��u�}����䕛�E1B�јf4�?�)sL�2}-j��Q�C�}�`�s�;m
8_�����y��ak�K�D�1��r��T�M��.��C������ʤ�8������ہ��A�~�"��q������V:s�%yi��*s�F	U������q��x����=�n���Di;�y�iQ����Y/��y���ʓ���yN+{�̸���P.�G^_�#Í9L�'#����
G�(H�pX��A3-"T��T�F�F£\�Q��>7c INb��#^�gee-MO��L#d����il���Ji4Wxn#*E</��䕄����N�"Z9�"2t+��e�+�>	�Z�yf�&r��@��>��1�lNC
�B��M{HhD%��{I,��3������53���#�5ʸ���r�c�k8_:%�u�6��!�@2?�y<on٦6:��̇���^J4���-׳�sdu���<���e<�la\�H� _�������d�P�O��z4'�����;�j��N��UJՆ���?q4��
�pi5-ݽ͑� �1&z����W�ɞ������}��q�4)T-�[Tc4p����%ZP70���A�:�����{���X�K�ܑ�tˤ���;w6��!m�:S!AD%���#�"vA��"�9�oCi�����D��cGA`���ϴ��VN�O�qe�V;-�Ay<��;���8Ԓ@�C�i�g�׈�T�[�6q���z�F�a����z�dsI*
C]�$��0�f�.�<r���D�ce:�l����w��c��<T�3~W�ij�kier_3��Dd�D���O��	ej��0G5�\#/�0��f� Gu)���X����>4Cx��G�G���ɹIy��������&��0���ڄ��������yY�6��X�j�������\�K?��/FY�5�+��	
������NT#���F����vUY�޹��Ǵ4��8�-�=_Fb�#�	KQj��zp��$*=p`�k�E$�a�����x��m�����-�A�`�<�񭓗4��S5�I� �C���{�^��4]_�����0��6� �MD��D����fD}�s��8�l��ߡ�����?�Cc�uW^C����n��K\ĉ�r�3�'��Ux2�%��o�D�Bڹ�N9sxaKxx<J�p�h�90 Q�OI<rtf�E�D�qޞ]N'���P<>"׼nco��j�e�t6�9P)�8O��*:���lT]hy-�NB(������ ��:�tU�]_>8#��k�nqw�����ge�9��N�;;��D�pҴ�:���EŇ�9�3�v��QG8xVa�Z�j��HS�����a��5H�-.SB@YC���1 X܇�?�!��Gȣc�<'�85�7D��Z׌��P��n�Lgy6���i��ڕk�2�,�ir�����{w���r�����NZ��[Q�"���땕�?�����!@���5 0-x�*�@P��	Q�:|��_�Vk�d˼s�v����0���.�\l�����T�p ��W�;�1��N*"�R� ������cf��O0��Dԡ/��v�11>Q��f�>���Ҡo՚S+k�}���Pe>[�:����E���W���<��M����E�� �R��2����4F�]B�F1�eآ���:�'?V-0A~�K��~�r��cQ��F��<+c�h�,��xz(����z���� �1���gLc
>�٬ȣ>5�3+>7��4l#��"3� Äa)gkWRV��dd��ђ@���� ff� u�B�6�`�E !�����x.5R
UO�/޻�n_}7��W��g?����O��v2}��oQ|/��Fq���k6��!ˍTl�5d��d�l�ns4���j��Lc��U��:�_�>s�ʟ����R7M��!5�;g?�z�sw�<���n/���z���cG�D���������g��:a�:c����,�����w_���qޜ�L9�{�������uS;Z���-�q��N���"<��:>�^��aP��!����2��!}�L`���#ߊ�&�1�w�k���Cc#�},�X8;""���!N���iແkmX4�5�u�N4a�����=�\�=£�I��W��/�V>�(�㒕���l�,�,�ܴ�W-���o�H'FGP�y/��y�Z8g}�U�@T��۔DYjjgƣsm��{���p���M�����1M5��&4�u"v�!�YG�ΐ竓�S��HX��rÒ@�n�U�"�q�B�K���T�7�*�p8�y�%��xpY�W���V"�π��A�h1K$z��7"E׽;Iڃ��g|��M�f���z�x����B�{�W13����uοwO�|���Z���YF^c���ZD����ʜ�t ��ܗ�oB��@�8��6��x��� ߵ�49s�F��&0�>� ��r��t�pO���/�1F�6^��V�S!�`� ���U���^�E`�3��u��UR7nܦ��IFE?���ƑK�鋿NE@�n���
�O�г
��l�Z{7��h}��*��"�1B���������i�=3l�P�h�����٫G��F*c��OE_'B�y-G��{*+RD�����°�$�ap�F�J�]�s��"����%�P�C�Y��J����w�8 cK|��kƤB�4'����PUŧ�'ndc�Bͬ�l"��W�2����0��0鉟�%�P��:��Ɂ]��9/C8<�(5�<�͐��e`���t�&Ց���XJ����ip����o��^yxv-�D8�L2�k�A.P��KG�Q�\��	���;�>��Td���(Q�:��.��&G�1���0w+�L�D�t��Vׁǝ e����t:u�4Uw�ŋ�D/���n��(��W^K�o�u ���<�z�p�vD��.�I�y���������7��T�g��M�WDvP4X"&���4_4!	�g�@\M�խ���H���d_���?|gT�ʡʁ��L{�o�GtS7�E�G$d�^",���<'�N4�tE8�2�Y���nd�=�jF�:WU���%o
F�����-�6��u'T��� �q(�W� ���ذ)�JB����r�lJ�CPӱ��� ���?Fh�h8�.?��;0���Hf%C�c��(��-�c���6���~��q����Q��q��NE�\�X-+S���`��gu��vj4R�����?tD3���U�岭�Q������<��h���e�w�r��b^`�3p6Xۛ��
i�N�΅k�j��2={�b:}��p��JY��	j�-_�;P-�2�7���|$��?�qy^O�@jE6�=�x�̧?Ǆ��N�$[M*,�\á�"�_�߅顙=S�8�߽A�d� EG<�.��K�M���w�T��e�$7�\�y�	�E�e,�;|"��`lh'w-� >����3K���s;P7�p	�w�r���4;a���֜Ħ"���e�v�W��2�7�'з90�ۀ�H	�0�6PZ?���2�yh����'G�t�q�T�OdN��\��pј���HD�gE/f���B�Fj�9�f��Y�u6�D�*���|��<|�s�|_ޚ�<y'B̥j�F��[j4Qh�~�ƌ���W���ε���+��x�6��dss^������W""������|�F����r�<ec��2�r�&hD��Sa�rͮe;Aze�rǝq�ч�{���pŉUF� N-��Dd�c$Ja�5)��'	%6ҕˌ�\%R��O���0lٽL�z񥏧��f�r�N��ݻw��!�Q�}����/>��Iw��vo>r��D������P��W�i�L}��U��G>Ɍ@�h��Y���k�5�ޚ=�(it�'�(nC�l^��������:f#���u Q��%�L����Rh����C�� ;C�ֹ�0���!�n�Q�hp��k[�1����f���qz18��P2_�H�Lsl��$�q�T��t;$Q잰�i��z���16��Q������2()" ���;_�-�����PQ����r��ƻ�f �vߣ)�XP� �)A�/�>�P殐޾�e��s�9F�ꑺ?�kK�jh�U)6ar"��tg�w��*�>��-P	D��Y.�7!����~L��xw����2�)�En
dD�E����M��5�����G�NS�D�����2��!�/�#�lTQ���$|��ie�&�C�_z����c�bބ��0�i6��̮���jS�۱o��UP��n83��4G4�����"���.����	��ҊAU4�a�K�K9�1;<x �qW��'~p������t6H��疧�A��F�
�v	(n�~�>C4��{�h�5�3���O>1�6�0����,6F�v_�m[N3<��]Bl9�Ȇ��w�;Ct�ikhT��1�Y]�hv»Dȯ6���!�����3th��䓶����.CP�[ιE�|��ʨ�e�@����M�#�H��U��aM�e� KY0��[�<`�Z�k>U6N(#�6
6��,�l&��u�G��er����b��_��g��?����_���v��Ѳ���D��Y2�-RX�����r%�\t�:�HL$��m������0�x���k_��2��K/�B6"���]��KW�����/�,$N���|��?������s��HkcT2�+�o�1�h�A�U�ٹ�l��v������Y��A85�U�#Fá�v	#��B8�9��ע�ݵ�@���|�6(�=��a�c($He�^6�ʓ&�
Ľ����W�N�9K*�eR�9z��viM8����,�N�Y��EW8/��т�˳���]�@�۷ɑ����4�\����M�x��-�'��낌���ӏ��4��9�Eo,L�W�}���D��0����
Χ��\���J[�F�{�y8﹄Ní�|uh�f��}),���;�k�qɎR�ו��8�D�[�������cф�M��ӿ	�2���=�0�PD�T+Ɂ�}�7_	o:��ϟ��� ��L�{���Y��3S{�ۙ1��\��Y�
�4�2�=q�i&��K�CJ���GON���Tk�ԏyu���S��[3���f]mw��9����ѧa�ċ ��VV�MiT8��h���􄜪}9tu5��:Ģ3�����Ԓygg�P$�2������t6H��F}ܤ����k�Gwc�O��"0�d-Y�[��O��"��2�@���4�-�9��ذ˛,��y�Uf(3pbַzYO}��J��d��s�ػ*�0�����z#`{LK�臬e����ݦiR� 筍kb؃\����aȵz��:^쇵�ٻ�=����\ë����T������$�қ��ɺ$�lB�L��y=D,�E��=`�
0�P�o���0�:Zk����~����_�b:ql4�i�n��6�Vl���ϳ�m�mY~�W�"�4���#�U6(O�h�X�@�2�����"7Qȶ������'oÌ�9��$=�[o��Ļ�8Y����4��޻7�/����p���V?��v��|ϳj��1�v�4-�9j���r<�%^][��	�<���]p'Jk�P��)�#1��\7�C8�]n�5�|�����G�0�!F.3P��_��)�����X��Ըw9��K���Ɏ�.��9=�����,k�伾�\�C�y���k�F�J�^g�]�Z��c��@%�zzV��0�T�M�<~&��C��!)����ŉ�tn�������[�[B'/F�nai%���u1��ʍ]�<�;ߑGzg��(kW4��k�+k�����~uv�����{��Rr|v�:�=����9����=)�#"j��g]��Ą�]rZ��C������M�F���ˑ> =Y]�?��~p��$A��I.d�p?G�K��ɱ�z�E��p�o��m󩋗.��t��>�&��:��>.18
��ʭ�����tk�;-m���q6��p^�^��?���U�r��??<'��QD�'�5,s�DuFAW6�(X�9<�C6ػR��MY�\�Cg�iY�����V��>�2{�19�i�R<ٻ4sp|��Z�M;+���G��'���7G	T���E��h�ej�/ߴ�f.l75��ҏ��;����t�Qgݔil.Ru�3ી��?TJ�f-��ّ�|�e�ֵIx�φBD����������+?÷*x�K�O��^{���`n��L4}�r��=��a�|cg�L+�s���7�{�aU<X;"u�1A��P�en�&�_�q�@�{_�e��o�GϜrZ�'��2���߇���:���,cN�H|η;�L�u����2����y�
&��'��[�&r]���	�kR�E��#i�p�V�D,{g�#ojd48t,���7碳�5�ѶW�h!fF�|�sDj簬нg:.&#>�,F��	�"��4���I�2J�\mt2��I�C5�6��Z�Q����dα�h&�M��X����S�\�����f+=\>ټ���;����g�_�ŝ�ee���z^wQ{�gu�N;)�g{�K�����r���H?���x�Qq���3!-��Ȋ������T�A�y��q���i���k��GO�����#�P��IH�7��&2#]NH����85�i��`�����D?6�/�k=������?ŋ���={\��ľuUgc��OŦ�t��D�r����&E�6���k�:!��9,":\:���&�lQ�z�>]���>���?����>�� :fvpB\=�;����56['U�5�ҝF�f�����Ϝ�����{w���M'{~s{�4�z`mb�X��D��ٻ�!�{�2W"�o%�m���z&��6��,�>��,;��fC.k�\n��? 	��M�]Cc�#w�]1��'�79����������`s���收1��)���̍��&��f���X��FGzcl�~���=�}�B�R+��w����!�$�{�!�����t�1Wg��a,z�3��?S��:q#+!<��8K�s�����@�R���3R#�؊�� M�+c"[+�l`E[�V=�5���T��F���� �&hD���I�K���u�6�PQyn:FA�˻�B�C�D�1#���LqdO&�hu���O2����+�捛(��8vXm~�FL��1-�<f����{+�:��lUBz?��P�Y��q���覂�=y.�1��ү��6��L(���2�d�0#}��ߌ�Q]��1����_IS�i,���|,o��۟��s�xuh~2�(ݩ$���	_n0cz�p�ZW�t�f6:}���;0���if��P�w�IT��ghN�Y<__�aCVL��c��F3��߸�c$(���^���]�| �Q�����i��K6�����T�����։��= 2�eS���$�t1�0�E8r<�� v'��p��3��!��XG:9�>��Z���Cц�3"c��
���s���ۘ*�x�l�+bd�����L��ؓ|I�t�'�<qB��8�N������s�n���X#�+GS������3b^�Us0��é��J����t͹��ۙ�^��G~>����G+�TF].J��8��V��bg�J����{|��{-�"q�}��{�ôpLf�Fҧ^�T:|`"���I���-�ۋT�D���)e:4���f��H,�~U��Y��"2 y�<�O����Z���]�[Qgz���Nz�:��X�5�������&��p�\{q�Y_��e��,���C�)�����]�����}��m�q�R�5q�>�1�y`]���hM,o��i�v�KP"�JH:����#4r޿o<���!".�쥜i��;W�����~�r��O�gm��K��`�6$	�[ϋ�Р�r�c���<
CtL65�Ad�hc���J!+QרFШk�����5����6`��CDm��ҏ�"��M�Yn�P�PC�j�m��o��A��QJt�&)G"G�hU��%b�,�p��Y�Dğ�ѱ:�����[EL��}�t6�+�92��\�ӷziqy�s�)��
Ghv>xv�3�ȵ�e�����ێq��,�'Tm�lx>��%t��[����9t ���+�����y��O~���ԯ|>�ݻ����{"Ǎ�F�o
����ƫ߂���p����ә��/�QX�'��?�X���t&à_�|9=��Ir��!�����7^M��(������I��W��P	�*Z��o{)1��M\Ѹu���b:4��f�|&Y�)��l��U��@YG����s`6;}<�#B�p��53�Ϟ�wa�ߠ��GN�C��e^m�J��wa緅o-A�p�1��L)��}?d5�*ျ��`ɔ��=���k�uj�,�&�R�:��b D�goL*���d_E~�g��7%�ѫpD�;��09*��!C���mfv�D
��N�4���al~�@��\q����{wn�A0��:m�E�Z� �9��TX���No�:T@��}��p_�#|Z�7�m��de��LTg�GԠC�!�Z�2�zP�&�f'��s���m�'0�q�8���}���Z�m�H�X�y��^��1�N���m?;�9��?ݳ�P�L(з�(�Xq-y�w����0��Ыݴ)��� �)'����U��|�)cOW����8��2cA��䧲��ԘV�!��I�vA^�^�� �{���OA�%X�4)�?0�Ϟ�Cg��k�=[��Y��*OGz�D�s��0�2�F��L?G��3��o~��Z+Ѡarr8��C��8�@�[q	4�&��Y���J�c��ˀ������$W�ln��jt� �$�h�%2i��r><r�U4jS����bw��&6� u�B��WG1Iޱ)���<�>�m
�r�6��k�kr ˊظ���&�`����&kH��*oXfm�� @��2+����Y��C�xB|�-�3���mn>kZI*��S����];9�0X� ���rL:c�D�#�[y��U<:�q^9Z��q����ϾU���Vz3�:�����0n/<�4p$9��A�/�6���4�$�ur�+���(�S�O��|�s�}HE�%���Nљ����~?Z���N{��SG�q�'�Z�;W���K���0�l��&��ߌ)V���8���o���H\����܁JI�P�x��L:s� }��F�߫�&]���a�v�k�_aJ��Y�_��K�yr�v���u{?MEΤ�Qg�w�{@��K���l�B"d
�k��/��Ȥ6��8ՃY^9v�f�/��lKk�0O��X���<R�=*�����Ǡ�3O��9R뼯S��Z��{���=��$��lr�<Q�E��;�p��M�����c���2���7�E���4���>,�ÈY{�kū^.yz��B��l���^z�����
.3q6�KQ�k�ܸ�O��T�ߓ��>���@A��F��+?�?z����S�D�b���CSp�@u2�C��o$�.m�Jdx#Cަ l%\��q����g�����O���p|T؆~S�h��q�
t(;k>���A��d7���"&[h�����p|NJ�p�C���Q����v<���.H�}���A�� �"4��>�2��$�IY�8��+���� ��$��?�<d�}(�i�n.�)t,��45�(�"�F�KݩZ���^D�P����؎,ʦ��5j,~��"���%Ym�F�vt
�3:y���vvw#s6hg8�Nm��WU��Ҍ�A] i�ƏA0��e�Npo���L��L�"����
�L�k�����AP�",��D�]X�hacx��NBVO��a(Ҽ��R֥�|D�����a���_ߧ���)�M���#}0D���،�H#>��i�� ��A�
�(���5
��Un(���s�թ]h"����W��M�<���*�����L�Pɏm�$��q"�P��nnC�i��#L��3��;�Ӯw��>h�׾�=zso ����󏦓����cy�����g���b�H�	s+KK��|�f/"���Z��� i?�;�u0�#�r��W��g�{6=��@���}#�\�s?vx?���� ��6M>�H�MO��{�ݨ��_�?�������/xe��ԘQ����p�z���`׆�l0��Y���R�~+�'�����m���E?!��`��,�Zc񆬄s���C�p���h��u�|Y�{�jq�ϻk���������GX�t.�b_��N�cD�sG��ßX_�5�#��8`�m��y?��FV���g!�7P����'"�
�p��3��*t����NA6��{���do!z*DE���ڬ+&)
=�&�fY�����N8s�Zg�9L���@T��@�X��<u�C�����y�=W��q��94������Wq��d���%�T�x�ڝ��#��B@)���@��0��I	��s��� @<R�`�S+ {p�Y�SZz�n�̫�T&�6���i�;��6��,�#�S�"�-��9Ň*Bg�t�q~����(w��B���Sȶ�̃�@�كD�ܓ��ai��Ju��R��*�@);[y��l�hroV�yb�~���i�~���;�����IT6�aQjt���p�V�"���bx�z���*#�MSe�X��f��˦��2Y�1}���],��� 5�[{�
Kj}�پ�l�N�p���(�ql_iu]��\�΂�D p��'��gTFA$s�n��+�ȳ�v�!��%�5���W���FF��[�*�_����N��d{�L��Z�P���!!eeyTϗ�m��}�J�v�oM`&��(.��W��{��Eo�6{�e�Ca}�Ԟ�t���t����vz�߇��wd%t�Q��o�}�$�� !a|ǐ�� i�`�m�Fi�O�����\�.��;���o�St|���(�Y��I���`��"=�'=M[کt�� ���hR;<`�܈>ܤ��?{�aK��Q�{>G�x��QYb��̞�J�����H^�|�9�p�ǿ���Ty��A`�A��џ��'�3��ȸVｋ�{�b���q��/��1�'[�p����+ rƳ���ka�#*��8h�v��1x>O̟�$���;?�?�Э���ڳ�K7漚=VnD�<�u�p�@؋b'kP���_�l���N�<�`H�:Ƭ�d2�t��edM�6��и��&c�DT�a�M��+ȸ����<�,��'ݻ���@����iehYÕ}��0�#�u�0�Fy�~:b�0�{Z�/�
�Kmܷ����-]mP��Ŭ�v]E�
?Y��bTW���:7:�2�Ȉ'F�ʠ ����Ed�z��h�@⦑���ׅ�
n���Y������F�F&"���A{ L�0ǲA+�#����	�I������l>��-�Q�ލB����z��P�A�����������.�b��0�@mc�3�-��F]M#0\�y���U���ı�t�:}��! ��?�n�74'HT9{��J���MI{��r���è2�'V*��yؖ�mn,��$��ڦ��D�3�14�Qà�����
ύ =�����#J�hݺжd4Ks`#c�������U(�g����^%,�%�ĭay^@��d�K�3���/�Ґ�R���<:P�:����az��U�9�o_yI�S�E[�BۍzY��k�s���pUA����5��Q\���M�=Ӥ"��[�d�hY:$2��ޤ��n�=���qj#�O۝.�OP�+3���|� �|���xX�Tl"� T�M��2�m�ק�YYZ�8><��.��FI4��K?�Ŵ�z��7K�9�f�&0���w����:��:p.�Ƀ7@	��A������.�� Ֆ�q�w�Thݟ��3��9r�X�ε�i�i:oi�HX2�萐�3�g<�lbd�7�����XVs@��F��.{��Y"as���b�U�W�W�OAZ������5t]v����,�L�|u���gr����8����p�>q}{�#�C�Ĭ:�Y��.,͑�ѐ��aw����9ɭr��"h3�Bגh��x�و�o�uep��67Wu�kF幚!� �!;��8�p�u��^	�<"|��93�!S>�?�1z��
�6�n|����[ A����:e��?�� ��P����kbf3����~by��L��nz�����HW�K#za�@.4��o�uw��]�/�reN�z#��ѾF��z��H������{=�9��-���!Cfɽ�F3�2�n����K�%؆#B������
3h���1Ɔh� �Q&.��_�AgJ������[;��l�L����H��z��b�W[�v��"�i��o��7���{�`'��cG`$o�ӏ�:3Z����E|u�'}�{�h�@4)�4c�a�l��B�@bð�O�ׂ����U����	�L��RU�X҃��:#!s˧��*}�."9qg�)�~�J8	#�*j�e��ǎr ��]�_�#�%��������oGF���ɪ�)�b4��(����jF��䒤�$���i�x�|�ǳ�@&�6���^fԢ c4�iёМ���ܣ����x"�;���w��=LO?�D�Y��V�ַ�G�c8��t�*���{�v��I��p�.Uw��%��{�4��q۠]h�Wei���~�f+��F�Ʌ߾7����8x��>~:�o2Z�֯2�㷿�C8��z�J�}���6h�{c1Dk�:��L�:7zV ���xf�B�]:KDB��KD�A��ܹ� ��]��n`�/�܇.08f��?i��=w!���!����?��QO�"<ʄ�/|�Ӯ `��i�|��<��c�,���w.�7'�=�]C�a��t"!��@'Ѕ�m��c�/�oF���a�"ES��X�F|� �[��p'��������Wk9���a%w��S����v�NI�����=&�]�p��q=���'(C�q6��~;��Dݠ��:N��a�����u�a\�_εߛ�S89w0����-G�}�w`���ՙt]C���-|-�/��:�׍6E�D�L4pny��o�r	�:�NST�A�����H�]&8����gi�t�5�7-�W"�蟜	�r�D�D�b/���Yg�z��U4����U��Pz���u�H@��Zv<"?����E�p�E,�Y<�u(�ևS��R�Mw�+!�	�_����[��ro*:F[[��ܐ*ΩVԃ��2�(�����#�p�U�����?��KQ�:w�,��h:vd����z.�����p|b�N�m�k������ŵt�v3ݞw�'��
1�x�6f�[��t��jqv�I"��� ǵ#l.�\wn����&������(':�<e��=Bl��Xv�<Wgoս*^�\�ZMC��
'��n����8�0�UC�N���6eG��@���%k�&�5c�9UZYA���x�+�ʫ�%��r^�a������6�Չ�܌6�0���y�w\T�11���?�����NG]��O?�^z�t�|�v,.��?�����D[�ҋ�?��;{�'�>!�w��q:�Nw�F�ۿ�?ŀ����C'�.d�y�][�"����0��?=�R�09�3�.��}�t���4��Yy"���� z���-������\��XZhn/p�}�{��$Ұyɱc����x$���^Т���D��S���]8�~p1��Ǳ�nݙ֧���������i�=�y��U&�-��}��P�|�4�i�ɹv�l-M$bB	���O3&lU���Up�En%�M�$���ôLV�n9��Ʈ�3�����F�ZaP:uВ�������\�w�F�:�fFJ��v�15C��ԑH�}p�F8k5��6?vvfo�!3�Ն;`^>�Y�A�זIk�����5�{\���:|�0��~��Aw��{�@$tIuݺ����aC��R�$�^�)B5Gr���1�3�s�D�r�&&��K�p\���w�)��vA�Vl��J����L�	GOlRn���hiIe-�5\�����wx������N���%ջ�$��L��_$g\/YSŏr
��C��.%��|��@"E�gb���W���U�Om�	8,V3�07�Rb������2��f{x��;#8�V�1�yǘ����1���l�������(]��uX�F���PZܐ���������nݣԫmH�gK�-��<WV�y��l�a��#h�S��ˑ�Ng��Cx��|������9��r ��ψZ�Q�-�'�.s}f,lK]�n���*��Mf-��I�B��Zd=���������/�,�GVN��*+��̤��=tx�묈|�oGO�
��$�Y.g-�O��c�c�B鴄��X*M��lb��A� bt�0�w2��z#?z,r�����ӝ[7ҋ�=��"ߋ����-����W�h������O��D���>BW�u�rHJ��p����W��jL_3��2վ��_��U��%���4E���%�t:)!���#F�j�̢�eV����`�׼8܎��uo+��W~/�w�c.��GOГz��=��J?Bx"a@����1��;����?�"���߭��t�&��t��.��$�i��t�@&L�Ds�Y�f#V=B�C�x�DǱ��;
���}�U���Q�r�*�F�� V[�b��*���3h�+��oTgh���1H��Y���eHf�|�޽;��7���3U�׮�� ��A�(�1D�"��1��=H���q�c��G�uF���8��i)sǞY��Ξ'(�;������G&v~h���y0~@=�g;L�
G�ja�m̺0��w�s�ߛ���,�
H����ӧ`��`��.=�#���e�~�x;-o����!����Mp.2��9׏NN<�I^S�f=�s�BNdl����JF=*g2����#=�w� ���49oT/z#��E1x�T\|&�r��nҒd<��b�����ԛ;c�����9��(#ٻG?9�ç��ZIo]&g[3�:��܏��Kts/]��L�r=ͭ�E<�-r������<{��wQ��˟��s��V��2���g<jy�.�朢	K�7��7Dd�r��_1�H���{������N��6ca��=�P���G�֫u�&.�rbSDUYɆ�ז�]�����\^�P����|c�ge��ZF<�S��C �\ͣ�����x�U�2clC�B����su䄉�Ǧ���(�A��w`:}��X��W_al�Uƕ>�N=�(���LG��Д��Ё�fT+ghA���O`�oG��g�|"��|�;���$���215��k4��|�m�{�=�Tc��Q�*9��qmsvuIH�s4��.uP��)��ӽ2�;�;���!�Ћ��(�e?��_��m]N�<'Ym��w�ʍ��k�s��w��3��~�!�1��{dO�z=OP��eX�0�(IE���ɐ�=F0v,S�1�&�ڽ_�{��B��:�r�����A<����Z���u�n���������:��D�NZ���A�;�'OF�!��X��k�15��"��ӧc�mo����jz��+�7���vY�2�}C8�:Y� :Q͜��p��b���\RVE�q�dG<�@�V��E`lܓ}�Q	ע��J'�c�uz��{O�}���@ڂ�"o�뉮{8F��8i;����A�γ��d�-�8��q�M�&�#���YƧ�A��nI5Ys�`��&��<��������{�-�MF��k�ㄇ�����YEϡ2>�O�'��Z����\)>g����?�Az|`ԣ�:3Ғҗ�@�؇�L�c����>�m���������C����0�b������CE�2u�M��`Eұh�n��Ǿ�ɦ1]�FD/b�@$�bstl�wK��Rm���Unz�SE�|�����z�18�����aZ�a7�}72<�܉.��P&����KS���W���;!��/�����99�*��Ȟvg����=��
���k~8>_p�e��>��v������Q��<6 �5�iD$��.F�Un4�N?rA�41���	m����r_x��K��s�1��ߩ�Hw:q�D��'_�П������(�1�3zy�շҟ|�;��Q`1%M��%?7�\Ow6nS�l�=��k]#"'�߻����@�*���W(��E2�\*�D߂p����<9�=�������;2E����O�yL79r����z�c�Pi��q��8����X?7GE�:�~�.e< ȋ�B��AO����e��j6(y�P�����S;rԕs��YH[G���0,������d磏���g���r3>�Z^XqjJ��w�]�r�UI�rb�TFGgϩgN�k��RF�.���:jM"��1}W����4�F���n��j}�pƵv}v��$�lУ�Se�;<��;0��r�[��p��6�;\Qy�X|ǱN7Ea��~�J�����UxX�c���6�����Q��2�\�._��M���K�}�\�U��j8�̛���T�s��^��*C����x�����3*7�/G�!��daf'�k�<�̉�qs�����]XX���0���c	�#��O�Z���`л0��]l�c"td`��z��S�?�)R�X�5f�I���9T�M���a-��N�nE�9JeQP�m8��2;Dh�����=�5pvd,iՈ����Z�����z�����؅����U6|��,���Goǹj)W['+��wB1�"?�sN=��{$�Ă���+w�D��9-s�:��#�9 aeӁO3K�s����U]�����|^�;9��>x� V�e��T�*�0����ʴI����e�ixQ���w�yV�Tٻ����"<�T�A�Wh�ڇ����^���>����Z�I����7ކ47�����}�#v6��r���4�y����W^���PA��O�	 E��5���j��MJ� �շ�`�9l���E��;V���tTp����:�p��T�_��g(�;LT����ۯ��:k�DGP�An|��EW@�VF�ȉNd=}�{����ch�Ҍ�� fņA_� �ʶA���	q܀�JU�sސ=0��p�S�y����S�r��j=U�6�!:���笸3��y�Y��1���mB����3���Ig1b5�μ��b9�ߧ�ߊ	T̌BR<	�!&��0^�}Q����:�����N�� �g��'L�/��N�;��W@1��,�����=�l�G�����`�ee�w�6��3� a�)�B�K�6*�s��7b`�|p�\�ѱ�#8g%]�v�~�4r�D:���c�+kd�VŐ@���Xi"J�>;o���k%�]�*���S��*_x�GF�᧕G�}��W��B��AB�9ɜ�xs|�����s1_�ȡ�8+��vA� zF�*�K7��U�����{�܄������C��y�����Fz؍�#�L�Ƚ�BpI�ǅb��#*��v4"�ګ��,�Ie�����bA��9B5���$6��Lk@�Q��k.������jE	7R�,�݀�9'TO��ig:L�����@z�-�N�f�=��lO�#R)�8��\ܒ�Ā�ܐ���{�9�������&׸h]r�\����]U?e[{f �Y��ʌ�DB�֝�ˮ^Y��>[������85���9d>C)���n\e���7�Ï *�^����O�lS�x.���+� �gYK����(��i�Z��p��\'im|Da�*����fA�~n4(��1���@?�#�����*��೪%��!D�f��W-}�� ��H���3L������R�o����Tjo�%��Q����*��cS�H5i�@k�m���s�' b6Q|"2�:'8>��^wJ� �+��1g���c?i���$�h
aJR�m�o�IÔumg]e�e���R)��?4�Y!w:�uT�e��]�Iվ	�?V�Qn�~}�{͙+݊ ��~�\!�<�z�˙'�Nئ����<�T���^����ٍ9���7ixt;"^�"�̺W�UT-�56y�_*yT�����bLj<���3�7_UE�_9�g����S�q=љ�����`l��Rtb��w��1ཬ9�� s��4��_����Ѿ�N�

�E����r �-�p��,�2Б�"������f�iaD���k���2�A�
LG��"x��sّa�ǀYt^3"�<w��m���ܼ�F�g1H����\�^ӊl�%��^��'E��w`�D�y��D?D�����6�+��<���(6���(E�Xfh̝�4�"Q�e�I��zn�|7� ���š�7W����G�0:��%Nؕ��.C��
jx���Z~�JFff.��j������#����^�$:{R�$�p;-c��$+լ[��+�"_V�0�1ؘΛ��7Pp}||�#���UJ�~�Ыt�v��e��0��&N��]�(��%\��X[[F�[�x/g��OP�.������Y!𐚊D%iŅqa��LO�>�����s9qЌ������Q�(y��~�Ԗ�#/��y�0�E�-��_���.o:*�]deXUu�Mt�˽�EO�:�'�{
�����?�ĉD�����W���w���f��=F{U; jX$�<j	���ko�|��-"�z:��.�=��=�}��W��^c}�ZE�8���h��z�o�!�!&�� d�ē�=���^!�aJ}����%r��0��z�Z�.2�n!�?��O3qk��R����8߽���|�|����a�4@�4���!:ު��Ó�ԇU��L��Z��:��H'���X9�<�NGC���u΃8*vb���"
s��SM?U%�UE�L܇<N�P�mR��C��'_�x:)ν:q�����\���2w�u��W�Z��e��c�����O=`��r�'l���gL�䎇:9��R�A�c�s��Ge�#�w�Ȗ��&a��K�u����z�)�².?a����8��L� ��6�m�{��{���D4���mrYo�/$�Z���MR�C���dnBv���������2��!(�j�N���e���Ι!O�����
I�`���)�84l~P�T��f�	U�,�j0@�1�|�~x}�hܻ{Z4br'|ɇ|�M����u��7/_e|�Q��Kn>IsI��1z�x�uGO������$6�T]p*L��c�.�M�RjU����xWRq06c�қ_�1��9�pO�$&��ػ�m��Oe���>[�0Φ|r��f����K��zoTrT�&~�y;ޯM2r�'�gE���l�_D]�kV�U�@x��<d'ō��������~"�)*
��9��g��]kN�����T�0m���5�}�א{�g��<X���'��C��o��oR~8��i���<s�Ӕ�����iﾙh���_�ٴ��1(f��@|z(���ϒ�勃WW��s��5�����K#=rpo�s�\�����rg��6D5[hv�s�v+�t�γа4�g�<R*��E.���}������@9�c9G�O}�3��'ǁ��0b��̠:0�o��?������1z�?��#UyR���;\Wo�؋�F�L����~��ڃ�DZ�t����[x��Q"�����}Ϝ�xl��P�9����עL�E针��hB>qo�>��������Jp/�1���b}���(h��J?�Qw�屫���uHe:!F�ƛ��N󘈘��N���\f	��1E#��{��S!�e�)c-�2ט���or���0n�Ͼ�zD�y��g�d�v�GE����1�E]�a ��>2r�7��H9�;)�%����v._FF*�M����Rb��i�=��=�#�>�v���V5�IY���W��N���\"��$��9�t�%z}T�x�����M�}��i��+"W�A�m` c3F��t��n
nQD�o=�7X~o��`�	���d=S!�ٽ���2�to��R�5J=oA�=Js�Q��V��w�R�I���!����d+<��L�z �A'���\ۜj��vix�)��n^+o0�R"¦q��Q��n&��m�����=�~�?�<6�C���v�7�=L��##Мc�SU��U�gD���=K/���22��5��5>�V sw�S�;+�e_i!v��ߕv��.���9O�6�hW�b�U�|�{*�:o@�5;��d:�';���4�p���_E,�/vf'2�0��:Vt�2�y"j� z�1E��^��D5�K:�܆�r��vb��;�g4:~yO�x��pxV!�&/nt�3܈�0=�3DgG��ƭk4~���a�v�/�����
t'�	��NPw��ϿH�j:���\(���at8�۾J_�e��u�Ɩ�Q���7�z4r��>��:y�<C~'��Q�H������1��ҥ��������ν�V�'Ϥ=�G]���bf�,���xz��gXd	1rO�\��M�q�f2�~,}�ܫ�3���~�MӐ�"�-���ٗ�L�	��L��A<ξ�A�x}���{�[��׿�o�ЧH��M%�7�u �j�(�[LU˨���Ԙ+ha_ｈ�#�Τ�\�.�$�aV�ѧ��,s�����Q�[�*�ؽ�t9'��X3���Ǟ8��x�D6��äh9�C�҅�OV���"��f4����� ǏReџΞ=O�M�Sj~�j�^��;Nx�q:��p��\ّIpվ���2�ɹ�<��=�EO�)�㾈���\�y˾`m	)w����8c�{pY�8�ΤXY��w�����G�3u�	(�&�<w�6�����i/e�Q�z�Ug���8�a�=�̯��Cu䫏uQy���_�Z��#b{[��z˺!沮O.�Xx��0��>��M7��g���O�+��!��UĔ����v��£���Ҍ�F̬�<V���"q� ��� K'XN�&�ue�\0F�14��25�2��W�8�
���ƊP6BL}�L��S�8CfC?�z���R��F��Ӽ�s���vʛ'� *���Zc�:G�Y��66���q�\�c<sj^�d�^Lw��Oލ�:Ƽ��$d��#�/�떍�4��)=OٵC�5'+��Ӷ�F��(���!���^_��J�J�a�g;E�i�s�������t\3M1��=~�P�E�_�cXI�t���۠��.�@��]"�4`�{(9s�N�����0�ֆ��]�z>���l5m,�M��ۿ�W�2��l����C]�a�F���{��p/�9�#N��S��ؓ}��XB��sr���>_x��������9i殹x���0���|��t������a�k�+i?��Ǟ|T
�HS�����t��Y:�O߄D8	j2̐�	j�u<��>7V���ܽ��9�pEkQﵭEM�X�o�ܞ藞SP�|�<�F�[5�lU�fX�hm�i��a˫4���u�i�KT���h�i�{�aF���Y���pax�(i�ҿ��c2�u;�T�"�#�FbV�
|�\�!$t��ѕ��4��Ng�r̟��'�k�x����-��������Ty�d9o��\G�0��5���ӂ��$�'��@0��}{銈,u�61b6��V�L��ƷM'9;��]��o7���Q����"��R��4"�7��C����\3�BʽXom;?�)�6%���z.�HTܛ�;��<T�B�K�Lv�z&�z Q��^�ϋnMG_����)����T~OF�2A�~��3�� �[b�i�]���q�7�х{�� �n��*%W-���Cd�wz׷j̀{5Sz�n"���hّKғy^K�r����܌ja廜�Ю�
N�Dr����gr��e���4Z��!��&6Xz���������+��+\�L��(8|��l�c�g딬��.e۫FN<�ad��U^mؼ�H\g�#�!d���|�I��"w�W�һ`����1ר9)��~�^��4p��޷o߉}�zn��5�,7����N��L�%*3��ԟ�o�FqF���T�]�M�՛W�+�~�aY��`������n�Ay�մ��,+�q|�ľ��g�A��8���5R�ְ3�3�R8�C���?�v R�c����F׷��qbRTUde���i`t��O�D�^K�����rm���̜t�A��W����?�����E���0��j|���v��W��t�#Np{.=KıB��2��ƨG�vȈ9�l��aZcMi��0���V�^��� ���a^��w�UGe���xUד�x�f.��\���^��N����bY��A�V��%v:z�No#�h�:��$#j�W*�ƿ|]΅ǎnp�1G�9��aSO�@�b� �G����h{;<2��6��=06�D�;�\%ne�F	��H��d$s�;w���1�<cT/]�2�^OҨ��k�+l����Q�X��`������V��A;u�"ts�}C3�I�K����y�Fs�Uk0w��с�B�;@��M�_�Be���M��} .�v��6�ݻ�:����،�>���9���c��*�nm�!)I����ʂ��d��y:9��r:ݔ��oP�Fi�h���_��p�\[�@��^��}d�'�x�5k�u>TU�Ik;��\�:p�|?��)ҡ�!��m��>���C�?:v��3�@Vԕ��%w���aγ�OF?��b:Pp7�p�W0�9_Vh,3^,ܜ�	D�Y�*����VT�BCAt��m,�]lP�U�����2�ݏ�>����q���UN/�E�m��r9��(�.�������o�`^T�~��mY�v�y���-s�*Ԫ����ݎ[ű�$6�p�"�-�f��"��%��g������#�9��:o�v:56=��ݲ�Py��F=�nA�@�lA�o^����׾G�mO4��x�YF�j#.�֏S�"W�L�F����"��)Ubf���d��"����`�����~"��ܩ��[o�{���W������G��Q�1	AU��s5񛪈ҿ��s�YAi���Z�����J����~��`��4|+��o�)��'q���L�1�w��)��u�Ht3�U������1�O�!:����i��;��`y��ōk���Z�=��9�����VV��=�XN��z���(STũ��r��N.!��*gV�1T'��i�Nw4��gGT�-:�5���,5t�i2	M��r&y�-#�����|�e�a�������g��m�o߾��x� x|���x%��x<G��i�$� ���2��*������'�y��tz���A�He@��Y�Zx���2F��wD�Az$�M���B�Rk�0�+�8�D��ip��	s�7q�MMeҠ����u��Ȉ��#Jg����qvGA~N�<IJ��{��Co����bOLl�y�.�hG�,�auD����࿄!6�s�s�N�0|>��R��5�x���1P��`91�j�����Z/Q����B)�>��1�zf�ğL��] Z�Xu ����0ʬ��A}<4����=ֶ,�d+O1"L�ܬ|\���'y��^�s^u<Q�Jt<�Ji�W��>��Ex����A;�r�&ǥ����v�r�F�� 	�!:�5�@#&��aFw�~q���+%kE�<Ɨ�AI�	;������r#�|����!������h��Fj���yɡ�Sn��|�}�g!��2��_�x)ݡ�:9m�k�C��n�i�e�l��^~�&�P��dUO���Ї|�(��.ڵAI�6��'_�z�����)�sD������ݝg��
�|�ȟcحrDaF�J��z���۩���tg~�{���;�+�d5������Ì����#�NyM8V�֨��/���P�\�����t�����@�0��o}�[1(�5o�O}�S�I:�E-2�W�thd�(b���4����=���֭t��Cm{�6���;�������R�iQ���fz��7 %����G�o�
܄W�5��v�����M	�~��)���ʱ����Ga�-�]ű�A�f��鞸�9����p`b��:�EB�Q&���/׍{�cu��e���e� �?oC����[U ��g@9 ����q�y���C����h�kt�T�w�Q˽"J���8u�T����v��`Ȼ�5(Ά�ꢪl�	�#b�,rR��O%�Ÿ�j��%q�������_��ݼy�gv�:�"���>�qtC����-Ċ�X�������@�,�?p(ƞ�q�LL�q����=��R��{8��_#��>����=�!��{4��%���<�.G���r��+~:v9&6O�d�T�5���>�1p��Z��qo��Y�(C���p�n߼�=s�* +�q��Sʺ�A����G4���} �����zsd{�5��޷�|�V�aHd�g8.TQ�����\�QAE�w8��#z�Е
�u@Lya����.`��3ѝq�전>B��\��H61��t~�R��s��;���5�l�ةw�܇!H��(d�f�s�Jиg�2	$"P��弝LV_������%�F8G1Fy���۾��,�~�4�H��6�O,W"���(���Q�K!j^U��ёp�o G���K����(��/s�{����U �{�΍��P�f�,�I=���Ŷ������u��u�r��j�NR(��A����qZ O�&�/~��4��>gڿ��;��D~)�о���G6>2�u�$����r+�[4��mm�
������'N�Z�D�k_��{�6���F^�����*���A����~�k�FIΥ;(y��z�V7�D�<}8������H��_���,�sm]0�q�������O}2}��[����c�ƹ��&�K��3�r�bz��m=��\<s����sl3�r��ͮJ��k����7��#`6�y���T��8P}B�U���a���ltɑ0w�~׶�QD�D��i�+��:�F6�=���N���s|��4��=~�h|pb��2\��;9p���H+ؒx��Gi�j/������e�IwVh,1��W^#�s�>O�� &�  @߿z�%�r�E�<cxWWX���:�4jqo��c��Q<�W4�1�䵍��Q������V _�!_���L�o��0��pY�Ni4�721�1���>;{�lZ�w;}�/��g~�i2�3��@<ۅ῞��!	�[�����:�a�ÜD_W�J�u�Gu��J?�U�&F4�S����Bh��D��^a��>��Y�RNG)�,M]B�����Ξ+�h�O�9U�;�Ý���~P���t�0��z1LyZW^�y��R��Zbmi�ss�
�*��X`�T3��s��s���y[�����To�����a�6� `��h�R͜��ߕqvJ��p_�g���q��Q�^q�$�Ԇ���mw7cH�4c�8��k�P�tB�Bn������b��%�H��R�9J��4�*��(���F�����Wc.Ԯ"�3�N��FG���*�W��U�v3�0m҆U��Qo�?�s!�EJR��]��)5R66�X���ܺP���T��wL�����'�Dc�e��m]� ��l��wD#�Ӈ2�(�-#�1��.�O��L�obh���{<=�{�y�_��o�*���P�Y���0τ��S���Q���K�^cr�ݯd/ۀG�A�f��L�r2R�V����9��ˠ᡼!%:d���b�{h�W��e�*�>������˫�1t�ֽ�t����?�7=��)��D�sN�Wg��O|�}���R&��B�m��a�<k���Z���:<N��9e�?�����/�wY�N�N��d_���[��7r5�y�㸹ǁ�u�c	��6`��TG�q�%܃N^G��#���
���rg�B�|�.�������KW��7�#�� ���k���v����9u���7�*�q������ud����s�3�k8k�������X~������$�p��?�K���͕�쉼u�χ�/���sI���\(�s�8-����8��^p]�~(�]G`��;�1r���Pj���Y!�S�|�Bb����Wz@�~V>Sv�ׅ�="�7Dֽվ��f�����W�B�ބ�rCx`0n=�J��=T���8	�;oE:Y!=���Ơs�v[u!��nN�d{�s���UD�`L�A� h��1�ܼF�z���_8x*��Sv�l��u6]�����X�kHr��:�4���d�p386`�L��	X�����ߟ�B:�Tb�x:�6ŀq����R���t�#sڈ��`��W��f��@�疙9��EW]E�ѣ>�Ϡ(�G�d/��.@�$4{�ˆ^ �Q�h���c�����yB���-���]�m�n�7ڐql�5�FLAH2B�����;i�!�^��D�^�~.a��M��oI���F�J�KKx��a"�IF�.m8"���瘔5Չƛ�+igdb�i|��E����N�,�:�=ޭ���T��}��f����(��R�v��8"k˞j[s����0"�hʽ|��q����v�zI���_}����uF���ޤLO��#����Z�^���ι���}7R��ƶx�A
�,#TW�G��n`�q�~��E΅��{��a6s$�ݢ�o���ƽ��^h"̽���1V=����Mk ��W�/П�繺CC�w����- Q��0$��L����@f��2G��GNEU�0��~�m��o}땪�RU������]H���Q�Đ��K���L�N�n��R�E����;T[�u�%�����Z�b歍�={���7���J�"tZM�,c��B��w� )�)��H佽�؛샚�hN�!u;˶�8��:D��$龱W�U$"��Ȝ�N�!t�"r0��c*B�hG��Bg��3�r-l�ZR+��mЦ�_�~:��I�H{�y��.`'���;���[�hdu��ߟS#��*8���s��\��0��������&;��p ��|�Y��誟*m�P M��|ti�5��Q���z��0H.}�~J�6�����ͭ�16!61{�>bL%"�Xe.*����Z�MP�D�l)�c�C;w�#�[�6�ϡLʙ��t��F+����&����b�Z�eF�1N3�����N���'�/_J��*j#��P�vF�F�Swʦ6'��ly��1Ց�$�P�Q�A���	D'�$a�rI�Fh%21�l�YX�C����U�[o.t��{d�˼�4�1�nr�d!	J���Їu�4c�s,��m)�{��t��T�'�wӣ'�{���/<e7�w6]���g?�I�?�z'����&��� �>r0����+o�M\	��nh-��/�җ���@�z��(�:�b4E�a,<,�1�]�k@h4�7�K��VwHq�KU|*������_���@�1������|��my.�X��'N�"�M�Xk$]8w�c�� ��v��(1�m��SGN2`7Xn�]J��o�Q�j�s����15��8�z2%��,�}���t#Ƞ��>������r�i�k��� H�����_������d��&�[L����!+Z��,p#kj�W��_�W�b��K/dh�{���o���?�/"���Fp_f?�Q�(#l1}�3R���7߁}~!]ۼ{�9�O����K���^���������	62�.Bg�"~ s�k�*�o���y�����1.��"���7�*�f;3�]�̙�w��x}F�����}�����{�W�/Goź�=�@���[}�S�;oaۙ��zq��H)�][���bE����r�}���>�_���;�O�O�g/�eV���mP��`F�L�I���r�W�{':��[Q���C��S����e�<� �Fu��-��:D����>����οh]�K��*����{�4J�U0R0"#��A�F'Ӟ�T􊸄�������t6a�&����F3s/�IwX���4lq��ш��N��J7W�?Ls��\T�N�yf(��+c6�cpUFl&�f#P�������-ꞷP�}���N�G�,��+*RHo� �|d�#��pݢfya�u6�i�U�g�"-qst�g��7�-�w4d�Ǿ%oY���������㘟q��(d/�9?�۷`�Z[-\xY���cR�
�s��(�Y��;�k��F��Q��J���{�3z׸�6��Ds�(�1"뀾Q>W�m�t����%�3ju�f)F���[0��hr�\�w�|�hMp.��ޚ��i�r��ݺql.=v��������=��Y�S%Z���L�j�b��sS�,׌���H(uv��U-:\M����D�C(�}����}�u3�޿L� �e�Gg���~`Rr�������T,Ҥ����sms9zD�`^[V �J���A�K��k��;>�D�4�	'�{0 )O�Ns5��7"�?�ǁ����8�g��뷙5�à�aCU�&�ڒÉ�	�O ���#���w���������N���sW��>s�t�C�C����~�Y7�����}M{2��n3,giy;���p�W)a޿E��.�>��6i��6dɨ��Xc��_A��$E-�k�r8�h	x� 2C�*���"`�k#Ĝ�nw�t�-�M���+Y�nv�<���]�Y{F�~�id��������0�w�6����kئlԡ4�� ��O��i��8�i��7�x�4��4J��C��`�qFYU	�|N�T���42�ѹ*2�x~.;"�b���&4�C���c�Q����N��o�L.�X<>��!��^��cjѲz9n<�Q�Cc��J�t����7�n���$���m������hT��H*o2�d	:�����qF	�1�10/�XX������S;0u�BnӃ
��^�*���DL�I<6��nu��jy67��;d���d�8���sΞ��N{%L�n�sf��,�$b8=r_y�Z�[��A�lAL3����;G���Q�؅c��ߛ�]cn�a>3V���!�k`��ڐQ���(�c��Z�񝷧'�ϫ��v�1$��K^�ƍ����(x�M�%ʙ�B��IG0����K�>�,p�X�G�<�V(͙�&ơ"�H ���"���ppT�ܛ��B^�I�h"��0���^Φ;�<Ɍr�A�qm�R��֮�(>�;�Ǡ���+�џ��1�ͨq��>��t�Ң���:z�<�8�����*�D7(Q#eC��Q�QyW�t|ns�4��q��>x -��$-ɗ$�__�&�2nL��������ԏ37�3H��;LΛk��ܐ���a�9���Dz��' ꑣ�fr�鐺�K�	�a��l����Gy2���O��Y�|��)�D��Zԋ��@F���e�?�L���G���VFM��Ҭܝ�}��q^�Y����O�_]�@�FS�^�1��=�h� e|���XA�5ʜ���}�W��b�򟥙.�y{��D��1?�@�H��%pի^A'>:ʹ���#��c'���#��Y�m����D�~б�wJ�&d}�Ϩ#N�㻧��9Ώ��EΣ���[��\��BW��Bz'P�wp��|�����A��9�� ez^7�Μ!ec�"����"jw���eԐ�4�}% ^�$���Iv���k�N�Є�φ>TḎ�Y�<��-�M,�3���*<��a￞�N�4=�Dd"�+�Wu����N����RK�jiwIQ\�
):Ё�Б�CA��`��[�r8;~�̴7U]�]�<
Hd"3����~�7��F���PY��g~�5�����^'(�%���|\f>r�;��F��ٵ�؃������ƍ啙0(�3��E�tT��|p��܄�j�Z�����欢@k�>��K�dAF7�97�Y�%:�9�s^\ղU��4�~UvIzs#�J�\�Ŝ%ȩ���N.C8��Q^��n�H�!�y�T��T����>�\�ש`2<�O��p�NaF5<gP˜���Bx��YB҆5bfW(Ց|�2������JqԘ�G9(�+X���q�on��v���@8j��h��Y���D9����K�n�5<��� ��=���KQw�~�g�P���>���_�J�w�ys�C���������¾q�9��thң�BZJ�а���Es�3O?=��Ю9�������v���!7X�4��g�@f�q�
Up��۔�T�$�f+~��ÛG��E�ԟ�|rx���az����е�����ps�
uʴ����`�݂��|/�_�[�=�n�9L־�R�y���e{A��4�
��p��eD���@�kX	�\O��6 �u��x�eK��g�}p���I�ީ�S� ]��ͺd�.�v�L$*�|�6 �S����q��~�i/R&�U*\���(�]�ڰ�Q�EzWQ�a��XU斲9x����<f�~�;ޓ��k�4W�;
}��Q�@ćcM�0���q�.0E�d����x�{ɉ��X�W��M'�lT&|����bIS�F�@���B�{��n	�{;����~�j��:��QP(g�ؖ1^�����?I�q���B�������(�Mj�I!<��/R޹�F<�{7��34��FV=zγm{�`_�_��T(�y4�'�)-��Vc`�<��(h��||�<J�v���}ָd�+���V�|��y6M��12���K��t���D�6�Ñ�.�w�&٫B�������2���k�~��7O?s���Ք2vS8��N�Z�g1օQe������ʱ�g<XZ�|�H��o�Za�딭U��.�,,bU��ϋ�b=T��˾-�r�xZ�S�/�e�����9�LP�!�� 5�=z����r7W'���&Q2Z��w%��c0���~@���+�|�w�����؊Q�m�ok��a��5�0LyC�E*C�~ӭ���J
��r�)��2�$�����<<|�k_~����#�h����9:��e3���|>��zj�m�{��E t�w#�9h�u���9B�6���z�ס����h
� n�+�B�۷|���JD�1iZ��q��>�8YB}��z�ں�p>aK�ȏ�ﴷ�k��'>1<��8�d�N��7�
�[30�i��)�bv��	��	����g�6�D�0��+��`6n.�lf��Ƞ��ʶX�6�0/N3�z��N�
a�
�u���m;��h����3Dv lK�4�&�g��^��^�!s�*�� �������_|�TD�!M�#��/рR
~AǫT�z���&߭g�:����Ɉ��`�1�e��	�O�M�zJ����P���g����Шb�뢸�:�]���
�������ծ~�rk9�d4|�J�l��#�n�|�֍�)��"R1E�,PsI:c
j��B���(���T�Q��q4
<�3�w��wϺ�Iń��J�A�_�n_�o�li���x�ﱦMH�� �J��t�̲>w 8���dD�`#4�%���d�_���lG��dUqD���!9�d3�%������-�P]�+�5:u�2?xe��q��b�,�Y2��9��7��;�J�Q�������Y-���������}`�+G�x�܅���&��'T���� a\�Tt�����Xҵ���"X�
Z^�m�,2?k��Ŕ���Rj3&;��n�FS�k���y���B��@s�jcT��[�j�Tv�Λ����b��&
�v�n�y��Y�:	 �p�
^�2���o#x��K(n�d�~ X�鵌�H�1^�D n2.�
��m��qL�&���sl���Lk	b��SbrЗಥ��zVU��w�p4�=�y;^(FBp�põ�'��z�R�f�eeW;��D��gO=5�c`��]�]n��C�J�x��3\���ԗ�:��y�?�2��dZ�1�kF�w�ߨ���Tw��@@^<�@�&Bt�8k`e�@NOe�U�ч���[i~2	�ε9�J�1�)�E���]{����6�}f�XR#�E�hH����$(�mÆ�;�q��Ls�m�6��O�g���V�f��wNCT2_���:�����~�����v�\8��;�8��ȁJ��8)�-���Fֱ-P]ɩ��x��Ž`�9���v�LԮ����?�O������o��E��VX�R��u�^��8	㐙��~m�b;�8ѵ��N�6�^:���?{J%N��8ƇD.*�ԥ�`7�Uk5k�cAl4�����x�+�c*�x̍�)�����"-_���Ո�������c��:
@C[�R�����n���K~�d��D�M�)־O���W�'�s�N ڻ��ä����{]�������?�'����I�i��<z8)�*M� i�^X"Rr�H�%���FC "Ax��·���D���^�k��#���5�S�څdX��*.M׌ �̴�ёwV�po1#J����t��-Ґ����Ż�ш	~��`b8�	��c���ZF`E��}!W����*��y����������O~a��]E��vZn�ƑTy�8��c��c�LO5�.�Zd.L�F��|�,?�>�A��֭G� !ͬ���:������hZ�wPp�Ϋ�����-���9����L\{u���]�y�V�u��%S�� ,���<�==�
����رɌf,���&;u���2=���\��m�нvcs�����;0��6�Q�·��XכһË�[|ۮ�����B�0<�����*8S��<t�=A�����-��tj�7���Q���
����'�R�n�E��_�o��,!4�i��e���8��[�p�O����}��%4�O�g��M	�"��֕rk;e7dp�@�X��V�y3���xف�2C�;�N2�;b',#2���-��
��1^�.����E>I���G�f�3�{`���<�p���R�=i�����&�._�1�2�f�E�!���m�F�8sb�v�h�}�3,<�
����'-� E�$��%���S���H�yZ�J�>]R�w��,�w�<���c�7�G�W4����0~�$�~h�%9"�mi��3�#��g�J]{�f;�	�k4k���C�|���'2�I��ly���\�Q��m �M�1^8�:���@Hyq��To�%����v���2fU�c��_y���F:F��@8#d��w�U�8�DFDƔW�:�ڊQ�)�Liio�4FUƞុ��ٞ��ַ�4L!{dA���:c�\d�8�z�Dl:�N���=ua8��%�^��i�p|�u�wX �֜ ����\���I�C��5���`��a ���}�y�x�&޵W^QNX�Wk�c U�� c<��%}���T�<6��7��'�Rb:%�FX��`E��52'n!�
�x�>�V)t��#��c��g����8O�r���V ���ڮ�B�buǕm�p�Y��a�W�]B�[����r�2 �M��B��@�ZJ��.Ű_NW�8�(�p\]@Y��XRѸ`Y�Z�IQ�5t�Z���I2�y*aTr��1&$�H��ROE��PEzji7��c�	�����LT���*���ɥһ�n(U�{H�β�bh�\$�w�Y%���$��ң��;�����{ �J̑�'<��@덳�6Jx���/>��':���p@��L��c����<�[(�1=w�<�gsk޹á��Z�Ks'�o�O����P&W@�K���$gj�F&؂dM~x�K̽mu9*��fm��Lx�e�nBO�9A(�����Q�;i��O=1>�;�N� @��78\<wq���A��a��.�'�~{���� �x��&���?�������+.��P�� �׮��wT�����`�\�K�w�����.�bVb��]��9/�C?�r�!��Է���~+F^M���Qk��Ͻ/�}�	���n�\�^\&2a��1@��ɯ�5C���X\��W���x��'�O��F�ʯ���5$���2^�aۊU><K��Ǣ�w�1�r���Ly�}�:\Kw4D��h�pLꕪ����k����zԦL)�r����6l����%r�D%���s*<���#�t�����E�d �XP����%�>�����I;����s�u�ԃQ�-��q�F�0��1�R{"M�"x��0?T^,
�����لe��.�k��Zv0앫�e�c�{��ks\L���p~�f�G#?i�ȍ��yQ'٤T�~�B_��JGȵ�D��}���0�/��6�lɫWn([H"��nc�Nccl��[���y�%��Ƕ�3�_y�����~����]����O��-�լv7K靮CK1�:����G�g����%�W=��j)3܈�2g&zSkv	��X�z,*-��<
��+E^f��׫+�5��@	~����0���*-<צ*����}q+��-�w��+7lj�Oᚐ}ج�5��1zPe!+Nʤ�-�9�#,�}�;�U�� ~�0��M�bO�ڋ�* �27����{z߆�7n!�ņ��L�$��'��%�%�(9p{��@hNH�Bn�p��'�[��o�]�����fix����f�5��-��׹��P�T�8&H��&��~d�ZH�� 6��F��ܨ��Ry�kϽV��)���]#=�RƜ�E��8�Ǹ�0�D>�^�&=�ُ=2���X~�:��ɻc\|�+_��<�Z��?}8�i7ф�u��cPt�#��ɑ�|v� Q��\��ћ�����o}�ۑ�W�x�1I.�0j����S���!�'�}��j�I�$6�W_�FO�I�I�dSP�
��D���]��)(t��rҘ ]$� \ �\�r/ZFI���������[O�"s��x�����R0#�(]��6�%�*%���$��0��mp��a~(�Z&���m����L�Գ��c�i����Ch�{�0|�j#�]��Vx��m�)3E�`l��a:�:ߔ�73.�p҅��Iz�d�Mk�Y�}���+_��p�=D.\+J���FGa�)��x��)X����f���f���!�7�r�̕Ke5�{v���Ҵ*�W�qIu�i����!J�(��x�A�`q\�?y���+SLڢq)J�7�`��S�~t��_x�5�;�OS�_��
�{�H�q���A�J��ߢ����<t����_�����N����GLI�D�R+���Va�BC\��Bw�ּ���]	�߁)����V�H�\e(�u�P�z�-�%��6j������k��P��0P��!u^D�h;v����<�ތ��^��b�x�mg��o[ϓ�U�Z �p�\|�i��<�PP�}��A��,��Wv���q%zj�7xm�0,�}�ӟz���ގ���n������ �!�v��e=��-йN"ף�n��Zw�2���(�D��?��'��Ƶ!�BӒ�I��D�O�?I{�9�������c�/�s���f0�(�J�͒� z��5��;w���g?q�����c��L�hT>y5A�y�5��$�C2�|ψ�mČ�	'5A�o����3��N)�Jғ�������a�N�M��p���-�����(i��۷��ӱ'��m�6��l':aG6��pϮ�i.C���Umt���Ȯ~خ����p��ùc�������e�W�����D�KD����Fm���Yd�^��4��Nb�XC���x�x�[�a��m]�L��rr�s��w�v�&��m�u�p��2!b�ph�+�q�d1)Wm�l�a�2���B���N�m;�O<���ڊvZ~<iA���1��
\ov(u�w�X8��	��V��Pm���T*��> ���<W1,�s����hqJ[_ז�O��jW��Z�B�Z�[\���[ ���։bg��pΞL�9��5YND���^dYK�i�濍8����0��geLg�3u�J�ƾ��-��,/�(�
�Rk�jP�b�l����ޠ�dR9�翎����t��0֯��p�����c��.̽{շ��p��f�Qj�f	C۰���[�зl����w��k�w_~���$N��l�U���%˺<�0"��V�	aC����V�YU�1d�<�N�Ŵ�XQ����0��&w�P�D���Y]��,�p$ǳU	��뮞Q0h���X�c�k6���_ee�0W۾�H�(�2�.h�RD�x����u��M���~R���yE��uF6t�a�Q�	!O�2F�(EXM�W�����a�4t�/���V���=����?�j�
�OB|xI�7oC�/S:�)eb�jl�4k�1\�%����G<Be�2�q�W)�Zo�6vٻ�0���gO��0��8�P���?s��u8��:ӿ��"��9b�IGx����:����?L��4���u���9T��f4E��;,O�&�J�>5S�ݔ�P�.�͠�"%��o�'h�Ǟ>����/�J���TG�ݯ}�K���\��7a����Dr�S��.y�s���:�w�(���v;~�V�G��<����꼝�!r�OS����[#:�^�u؄C�_<�q\��=l���wE��!h�2[	��zܖ�i��� ��>i��:D Ԭ�� �ÆV����@�u�dp�`z�l����p׽���?:�ѷ^"C���f��nlD��(=uC�2ѻ7�S�,��,���TK|�}�a��WJ�0����N�MˈD�&UL��P��x��{���"�g�QD/fm��~���S���Q�c�#ytx�����������I����B ʠ�d�>f��+�%.��E�q��2�?�Iq�E�V$�A�L�)��.�D�b�G�3S����?]�k�EG��<��M$A�կ�9&�x�r�����YG���K��4Q�H��%�������=G)��ĝ�O���w�и����EW��w4K�3�R�{���x�{�|���G��� �InZe��ٽ��5Ž�s��y�wֲǨ�U_�U*��
�o�R�ň�*KH
ei
GJ�D���X�k�O���/�����ԮL��S�{��5u��nk3�͚�4��U����_6��\�2o��x��c������q]R�������{e���+�&-��9��q�ׄ��"*k����F�v�4��$�|彄�S�Ns׎�����?��%C~v�j�������h8r�����(�q)<���F��/������<�|�&$SX��U����CI���7��h�-v��>�9��%r�o�x������?{f��W??�s�]����3m�̋��?���{�Mr���m*«E5���F��<i����>�&m�a+�b��ukC�RBB�g��~��/��}����cg��|c����[�;�ޢ�����W py �>�����W_(o^��n1 rw_@�|���"U ۩8x���<j�(&s�7{!mI���xſ%;O�9�!(-+��)n�u��%5q���VR0�8�aX���gO �˽tB۽�s�Ϟ��"E#�����4�y��=l=��%h)��"0�I|��6�a��l�pN/�J �.�3Ģ"&à� s������Sy�t�.�|�*��0ȯ��H׼�(%"oi�J�A���?�2�3@�%�{����Ç 7�X��p���˴Q��P�����B���V��R��
{(���J�X�1����#�-M�W":������҅k2�7j�g��&��Y����;y�"��e�2���Bq���q����uu�5YX��B�wR1�W�YƉ�B���֩4��$ұ�$sc�@இ��ި�u�r�Qƹ��po��3�k�Þ��U�{wm9���?�������;R$�ۍ�̏W~���jG+,�{_�e�zy�	�6����j�r�}Y�1ݬ7Uv�����	(��[H���:)p
<g�iҚ$���Gf57C�k^S�#��0x���!G���1�sݖ	
��M<��w�G�K�Q/z�3�M?��K ��s�3�`a#�3�����R:��!#��g~��_���XƽlD��s��!�;���c�B*��`F�z�ό�}�ci}zLj[!ZٶmԔ/�` P��a~^y����{� ~�S�/r���QH�ڥ�=w�B����e���,�kMX>2\:׳^'c��/~ƶϣ$ls�n8����Os�i�f�9_��?�좘��⪬�{���m�7"���'�D���V6�]��)
~�o�wf8z���*���^#n�&#�҅m^�������/e�����9X�^�zI7���������;qb8��4as�l>v��������K��z��$��e	͆mZ2N��3��,��
}��<9U{ �~�V)�5d��z����CQ=���o��o�?�di�{�^�#"��h��q=Jr��q���p��� �����KKj�~?��ہ�4�,�0��I���oL.�ߊـ���(3��NT(3S+�V�W�֬�:�k�&]���#n�WSf��{�H@�и=����/y��̺`�v����/�w�F(�]#L����w��%�5�c0r��,�*�5J�%E�]k�Y����-T$$����)�O���;�W��5Gc�	o6�jL?)O=?qz����_o
=NA��0���{�y��1Z��]���%�)P��a��ņ���c5O^CZ,�<^��������ڰ�ͮ��1�x�#%:A��߁�2�w�㱇�g�x��g����I9U<���s���p���5�Y�a�Ҋo���D(�n�D��k��c-���dE�w-A��J�N��1�7c���OJ�������]&e9�)˙��[���4�n��zфI�,m���4�1) �qC�l�����[u��C�}<�$Q���<%B��]���ᓟ�ܰ�/�ia�(�ؓ��m��wJ!k谾Ma� x'a�250C�Q�b:��Q���h`9��۷w �߆�� ��V����7�%�l�T���xQ��̅^ ?|  �^ji׏�Y3[���nS+~c;��_L����K�W�f��"͘=���A���Ͻ@TPʒ�%Qė.�^z���9�O~�b�,��$�n����a����Ry�z+ˤ�Zܤl7?Í^�(4��Q��3y�UD��_��%���w �}XU��n�p���p�<쮝	�26���/e
]�"FM����?:a�}��í7iȂR���Y���O���V����.,�N����6��OS븧P؋\�d9r�/��fHl�&��1���o��'��U���W/�?>9��֫ÛP��Zw=`3p$   IDAT ��sg�W@L\���שHI����GR�=�(q�e�`]�f�ӻvS�G�|����%j�W��H� <�&�c3F�QV+{�4\lz�r2�y�.\EIHH���Ű�J/_��h_h��C���-Q�D����s�6
�:|h_�yS����ktE\�f��zɇ�������p�,� ��n�<���N?���kF}�$ʽC�h�"v���E\E����Q(<wu�U���uu�a1�WO��,��~N� �}����!�}#�E��T��	qT���~���!�Ns�]$�˂��֭���~!��됏S�O>{���1���Dy��`Xo�`o��L����رuәO=y���_�z��.�!��M�#��4��^�9*:J��p��5�\u-�����%���Եqr����"����a�u��z+�o;1L��p�g4��k�߷�f���-]��2��ɵ&/�񻐚�C�O�y����� ;��#��	"�)�w�>IXj�*���>�R(���X��'�dNQ����o��ɒ���N���ƾup�I2�	J�P@v���[zQ��L���.f��P$S!�XG�}3 .�Ֆ��x��@D:G3����{(���Ո9�iǦL��s�]��~�>,���_��㝆8��u�'��ƅ�����2���w89P�E�^<:�-� d����C�_���c� d���7�S���E�4x[�z^JŁB5kb�e��hS	�9Q����zs�+�G���-�3�#�-s��= �1<�1�jv�}�5��1@;��N�B�(�����e8z�I��g>�����4�X�i��.�X��g�NtK��.�t�ˆ��v������7|�k_L�ȵ�X�D��(����}ï}�K)ۊp��ˍ�,aI�3�x�u�FB4��W>W���L�<p�R�Y�SD{6�ʄ�%@?��7���^��v�wΞ$�����o�9n�zy�:�r����/
C9Yb%��{F�]��F��Vߔ���м��i���>o��=f��b�S��r^:OKң�R�~6��K��$G|S�ԩ3�(cؐ�غ�ѫk���]�DK� ����LYY����)y�#������@Ύ͕5�S��5P
�=�w pS�~4>�m��y0ߡ��s�Oc�})!��}s�^�ޔ��9�������e"(�]t�څ�2GqF��LR\`�X!�*J<ӚXc�	�vK՛C�!Me�v
�[�/Wqn�
vv�3�s���M�J���u^�;����gXf+�֑��=w���o��KO3�����.�{X�gnҸ+�rU�ٔp�[��n�}}1�3�e��Ϧ�!%[��RSC�y�Y 5�D��S7)*�M�a�B�V`�5���$A1��U��Psj^��z��	��Pg�!a�(�Q	]�Ra�s�E&)��kž�\��a��|�S�L��	���g6�?��%����5�^sjfʜ��b�n�粘Y�q��w3j
~�I��aa-o�x%l�=�^�u�� �}O����E��^�
��;�E �Ea	tQ�o�]��Ӥe���xtR��g���ߖ��Ǐ#�~Iu�e�C=0a���}P�.�+�3������a���a�P�8�&���.��>�3 �g�tv�4���p�R���j���kU�W���/��ʩ7�o��!]C��q� �	� ���D�e4�"BO�G�<$�˩`@^~�C� ˗��Z��zJw2����w(���A"�|�u�*,p׮<�;%Y�� �nP5p�p��y� z�(3���݈�߶g˰��^<�}H�5=4�{��ݤCLsT�9덥��B�S��gݱ\E� �S��;�4v 㬰V}t�f�T�Ft,s����MM��=�=�%�ћuo�r(ίwm�Pǆz�1�܂��_!��@����$�	W�%�(�%���3�g�\�S^�v{=�G6o @�r���m���ڿ��3���0����t���*��|��!�q�L�[6���h��S^KU�p|tye�j�-9��+�ޝ�ȟ�%-�V��U)8���X��w�=����������Ż�h)��$�M���X�R `S���L�'0�&Ѩ�qN���X��A�}׃�Ҏ��bL�MCvc��N���S�S4�_!�b.�ֳ�_�^�^>j*���=OdpE��sy����y�����f��q�,��&����@�+���"$��e���������K�}a~��tr��D���圜�!P�pܧ�\�Mq����QZ�Vv&����Z}��t3զ���B^�ҵ���Q����5�n�W���lFØf[��	[ī͢�+��r(�(v�=>7)�Ǧ4��
�i��(�4��#xƳt)CH�=�k7�bl�M�N����>�ȣåk��}`-�C�[ o�^PP�Bɰ_Rd�^��Ԯ�s[��קj��
l�jyF�-(_o���Fw/{������\��z��Ȍ>�ƶ���ˌ'������ߊ�sp��t���������!�R��?}щ��aɟ�y����>?������3������C����jQ�C�UJ�n�'��8ky����k��x��w��� tS2�]��%�QV�����MWs��i��g����)B�A�kt��o΂!=�e~0RTl
s�3�߲�������w�G�/3^��F]�g!I�a��O�1���&Dy�����w�	���!L��庶�-MX�ߵ-k�P���}ix���׿��a���Q�B�v#,),�~	ı����qu�J����q�4M�,ˤ'+�y#&��W�g�̏�����5��^M��p�ܠ���w��4�n(︩:�M>{։Խ�B�y+9ߔ�aL�/ʧN�IҟbR�s���xQR"��h�}Ɬ�N�$��=��m{��)<ދ쩭܇��}�ꆅ��so�Э��쥌����Pi�5y�z��H9A�+�%@EdD�Q��v��.��&K.���,H�y.I���*4ܛ���'�޿���ZJ%����!�Iw9&�.&� �OR�'���H�T�:�K�j�rxb �4�Jvi�o�Ny��?���1_�B0I��"'�UvIQ=�a9�v.^G��&G⸭��������:y�FiН���:�� ��,�u B7Q���kM0�����dB����+� D����/�f����Ͼ����჻�ڶe���k����|�Y�Y�|1¬��K-��b������ب%Y?���:(��� Q5 �lY��Zzx��&W�V#_%�&+5��ZB������ZZ�*�7L�MKī�׸������*-QAx	>��3C��~�)�0��g�ҙ��~�7~}��'?3�M���?�%߷��������JjcJE�D�δIHVȣj�+�h4�'�rB�MIHf7��G�=\V�r�9�/�vlx�$%*ze�ъ� �=�����*m�w?m Q�����
'u��[�m5w��-��?��?E!��瓠��s�F�ʹ�\�Ar��J��V�[�.G���K��g#@�c����pe�S-�IP�y��Q8(W9�7m߭X�ב��G*@C�x 8m�⨨8�"��fg�ۆ-c`�*�OJy����U��u�~���a֓En���s|v�I#E�k��/�>�w���O=	z{wJ�ާ�t�70�j�v&����t[�V��}d��Pqz��yǍk�*aRk�mt��·���h��}O�a���s�'IL/�4�SY�G�ʬ��84U��X���]�z�f����w^SI�$�o%��G]宁gT�p�5"H�C��Q,s�c���)����¥�wm�wH�=GD�hɲ�!]a�K�G��rͨ�
x�fOڹ�u;Ѕ�^/?.Cɢ.��L<�R�Պ�=�_JFm���w~�H�|���F���N�:����L}P�R*H��%]!�`�E{V�FS�Yl	����j�UT��=�h���Q=�F��%���á8��Ð�<0m���^���%o���I���*�C�)��͒�g����ȣ����~]����ggΜ9���G��w�;��0���[A�'���2�^��K��O�����B��ҁ����7���uǮ}����z��g��^��JE^�Qy�U��|�ۮ��s��*�Z�Q��FmSb�TyQF�Ik��
�z/a�&L�'Ne�{��Q���d�T����"�L�eI��9���T�CKڒk�> ������"��V��!*�x��	��+�_����-�YM^}����?J���h��y/��-��Q�������ס ��]��6�1�d����9���}�<)0�9~��9(IסP���?��0�n�<���	�ʾ�Si�zk�Z&��EU0�P�i�r���pZ?��(z�P����������ީ��׶�'��硿�x��mx��8��MԺZe�o��@޴��-���XBG���ـr���
��J9�ETt��4����+p�V����e6��D��M-���eD),���M������TET�W�[Ě(�ϜuX�4�l\=��:���(QQ�z��p,�����~j��ٿ��9؆kW�%�:0L�x�_�b��q����DE-�E%������L.�֏�[�KC���3q�~bx
�)��\g�T
�5���������fW!������*�5n��?��Ea���q�:��Q�����^��d���*j7�n��+�y��S�� ��`P��|;������4����5�*��!KX�w �`����FH��f
$*�~��5���ipV�ըb��x�h$��M@a�A������8�.]:�:�+���g�Rr
 �c��O�%2v  _��0)�2�zym�%�#s_t��=ȝ�G�4�w��?���vqn�I�H�5m~��M��cvX�YX98��!qg?�H�2��o����O������M�lCf���ʱHxK�P���&�5?~bx�w��w��K����������^=1�B��ށ�a-��)�Z*Z��a�����^eg��?��|���6���\ˢ:�94=|Q%�O+�𼻕��Y����
���h��i���q���"�=�0*h�ɍ��k�(�<��@�u���\�}0�݆bs���[g��t��3i5-p9�}��7�W`esL��'$��1��иz5�p	�4˝y��l�QR�6��1��=�Ǣ^�l�����s_���Ly���)�E��� ol�4�����x&֏?�t��{���zX�.&�.��yʵ.#D�?9��fx�╋x�(h��' SQ ���+�ߢ��p�#�u����y��e:�� hs
��4h�M�\_�Z�.�i�L	Hm���lԧv7+p���x����5I� ���1s�G��*�W"6��XVS�<�&�r��v��t�T�(`1����=8C��0s�u�BL��Hs##��ٍ�l� pr�|pRx����N����u`�v��`=;OZ�����gZZ:&�M[��;aw5Uc%^��DՃ˘�xd�a=�Z7�Ʃ�� #�i��{ډ�d4�j	����S�yH�����ϕ���A������:ɕl�Xe�7b�x�brR�ǜz�@����#�]Z����C��F,����AX�~����X�{Ħ*0ĭ���M{$F�n*:�C�y⢦�ϖ�o���eZ]q�#�zİ��+G��%V��҈Q�z��ƹi}x�H�87����V`��#�脚��]�V�()������O�E>�qSUE���p�)���[�Uhf�t#6���w�t�4�j.a8�h���q�5M#{�Ƹ��F��y���qw��H��$N���˟�Kߓ0e�Ͳa����`���8�m�9�1��իsc����?��//8rd�ʆ7�����%�'j�Fb*�lH^�Xÿ.�"7���
�<(���КMu��X����aǛ��G�'��煐�Nu%>�@4o$�X�IՁ
݋�]��}�@d�ғ)O.����rb��K��i*����9?=<3Ӈ�SL㍢;�%:�i���کKo�{�@���}��a=1���ئ����3W��|����
$#�=fd�KƘc/�/�kq�5�����|��+�P2����I��N��)�Z0��G����pmx���ၻ��m�$jq�w��'��m�zʓ�06�K?���������[�3��w8��α�c��BJ�^}���_���߰$��U?`Z�{�K��?2����õö}���H�_���w2,���7�d׳�Ab�	�rME��g���6{|�0��+��(�|�<k��݆��`�`|�"ѕ�aˆ�Y�z{��	�TҘ|;��;{)���h������g �%-�yB�7�X&0���ݧ��vq}�v�Q������瀢���(^���r7�n��u眧v<�Fj]��.�x��&��S
?u�*Q[`�	(�s)��1����Cc"���@�4)����^�͂�gM�g�R#ʗ��� F������MR����i�k�Gc4��8�6j�ǝK�
�v�(6s�+�Z1�&0� ^Z9Ri�n�t9e>ηQ�	��@	n���y5ũ�X�f����u oL�D���c�TT������\C���M�D�8��K�Vj)<(�q��,F��=����OzcF��w��8K:�{��S�v�؅��X���?�1�	쿆���7�:B�[!��6Ǚ��@�h#r`'�4n�y�ell�BX1��:�ە��#�ޑ
�|��+W�����Fk�u%�7S�g�k�;�e�*���� 	�]�����7�?�%8T�0E��WCI[~��S!ބA̾Ֆ��a��vQ�6��@������+x|7�ӕxb'<ͩc��*j�i��v��c\�7*� ��ZK���r��-����٧ W9S�f�i�T�����)���QɋEl���v���k4do����/,�0�����-���K����^��PSl����K�\AP��K%J����>4R�6Jƭ]C$v��\���K�;��<�0��9�W��?ǂS`���\`.��֓��G#���
�/_��'oE�l ʰ9\C���6�w������@���Ȟ8y�\�g��g��ǟ��ߠ��������<ш�B�d�̟�Ռ.g_��g�3s?�N`<Qs���%m+V�-�6?v7��6R�Gͮw&�����dK�k0�8�m�����9kՈ��@ ��7�P�J����W>�E�4��R�r�{�H>r���[�AD� �8��:x/=�w�N���c�""s�����^j���KxY���R�!	ھ��1<zs�̉{,���3o;�4��GaSa��p�����)e����*|u�"@*{�k<��V� �|WJ�*/<@�9a�I2њ2�Y*oհX-Em�<8� �v�u��=])�� ����o&q{����}�Mj�E)���-\���D�d�xp��H�m��|(��ua�o$"b�}�X��˓��T��.����īL��z��v����k�y-2
�@���w�h]_ZEg�W�?^�W,��{vo�[��ƞ/�k97��7���p1{v#�� �i������x��?ל�er=�Y���\�r��D0����{v�[7|���sL���~���W�&�^� $�ug?�H�~�ԩ#'O�|�H	Z�g�}�k�\�n�s�K�IJȓk�6�6��<����+ִ���ʭ�{�&- Il�EBD�(�śsxy�@\'$R�&
��XS=��[���%c�;�E��$��4p�������Z�s4���5OKp�x)��WAf��\��2��xM��n�̳�F�e�bU'�[�\n��Jql7�����J��S���KM`� �������b�����
Ԧs4�0�+�ױ�4̰�5�цʧ��yB���T��Rꞡs��Z�]���F�	9�Ζ\��*�m;���_^y��S?�MZ6 �[��(3�&ϼg��?98xdx��W��������tl��?�6ㇵ/�6^��
䓟�7T�������_O?�<as��o��0�#�>1<�'i��8y��a;(�6Rw����a�#wSK|	0�ld֒@E�!;q*�Xza���[���0{~�Da3uT���0��4Ѡ�z�T��A��r�m���f=���qHtf@J��:���������$o�>�Y�BD��W_�P;9���Cۜ(��}[��3��/���0|�;�a��°�mx��	��a�!ް�3_��D�l����w�f ���xSU
֍��\E)��P�p�bK��Rajy��i���h�0��|V��2"��*R{�4���u=K�E9�Vl$Ǡ p����{7ǟ4� ���@���gs0�V���-�#�jS�4�߫&+�����C������f�=�j�ltG^�TwW���N��:�:޺���&��#�+�z)�b�@)p�aq"�`�h�YQ^�L�t�\U��C��~§|��$��6�zj�@�D��b���F)�ܽ�����lX�:<��Z�!Z�x-"gM�1:u�-ڙ�;{8<�1rɮxa��K��O}���U��t�A:�8��ݘ�ٹ#��������I+��O�}�cOgE�)�Z��0���J��^�Y�r,���az�aRy��� +ih��VN/�I�h^,����"�3�ۻy�N�3
������R.D�,�V��Z�a��0y����}I�����uLM��ܼ%��dֹ�mEY��1��8�}��{�2���d*��e�I,/���?<>~/����1/�cv��"u'���x}w�;�H��l����*�1��o��2<��e�ȥ����+Ϧn �[�y��+��� ����1x�7 �D����Bk	��m�l�R��r�E޿�k�@�ior}[�������={@�~Э�
vD ڿy���ã�?>9�o�s��e�;�?�$u�0�!�o���۱��Or�7�_v���������!D:#rnu��AY��-AZ�^f��1�)VÖM�v1�i̼9�����q�(�~�K�n����7o�����H��F��9�3' *�t��E�V�` �9Ble{��n7���/��E~�����X�4<���ý�>8��|��&
�j{��U�SC��S^���U�rd?VɢUU3o�Jo�P}�k�ʍf��C,½W������(I!�et�Q)�2���kz�r�e-
�2����x�B�=L���R�֪�M}z����[Qyxe�Z���g��c���g�Lm�5�%H5��>+N�D%�3�-�]�'�v���-���G1W�M��y���0������.J�v#��,�������h֚����U�2�6�W���z�y�Y���*'� �`�H��{�6�� �(s�M3���t�#�~��0	6F#6��ѱ�TZ�N�Bރ���r��q���C��Ko��2|�3������9�L:�$2�f����8�n�o}�[��A�_^��X��(�<�z��E��z�*$�Hy�.P���Sh{�fO�AY� ]���p�����V��`^���������˽B=	�!X�B�)�E�P�T1�L&����k�
d��L�*2�AJ���O��|����P����+�����������p����ٓ�-x]��W����_{��h��H�^��vj���z�8��`	oE=��iȴo �6�N����}�;�^���8V˝�97��R�FTz��8�����\)1���P���z��P�2���%	ḗ6��Y�v�x���C��#��M���`���u�@z��!��/�K�,?F�$?�n��'?����o|*�Y��]��3��=���{`�]8�#Q���?(_���(��n&���YG�b���%X<#��#mL�5E��%������4�'�ӷY��>V���w_}���9|��?�`r�(�R Nӡk����
-�|����oE%h��,|��vh{�8�~#8B�{ȋ�ݵ���ѩ�T=l�0(^�����u1AM�}�e� ��جE���T�,'R����*hhS� Ī�-u{��+��27�?Rѝ~��ձ�J�E	������f3:����X~�?z�^#@iS�x�[���|��gYثƇ׬7��ZU���O'R5�an%�a�u	 �����5��,Է��������:�L��H����R�f$�Vz�f�^]s9�e|�,f�IZ���?P�>͞�c{B=�����i}G��|ט��|-)PC�R�{������O�����wŎi�@-6�5��/��c�� HSeas�%��H����s���N0<S�dY'���8F�E��]���q
���an��.��Օ�����X-ބ�0�W�2�c���7gABzq�&�{�����^�E�j��ўoʂ^^�:���K-��!��Mc���Z�|$H�\��t&,����Vw��b�1S�{���)B��Kt�EX1NE6��K՘(�H:�����A��n�@�w��+�Gu#I����w���g>���y��~���D���&����B�*u=����e�T�8C>d��K�'��	,L��j�R���o�)$���a77�|�O����#�d3�]�}�ʟ�ٟ������2��K���>����j�5潯���M���µkW�9���!�Y��h��2
A:;Pdy� ����Sǆ�}�Gx��0���W.۶n8����ǿ ��hޛ��q�TX.�H��C���D�G��Q�+��9��� ��f�Vk�Qҹ��%�#�b+�I;�ɰ%"�҅�Ʌˌ���ު�����t�z��qx��'� �w�J_n���ٽ{���{�)L��fTqæ��&hUJ��Ш�DK�Y:��Z+�כ��@���_<|�Q:f��JPy"����p�K6�_)��0�5���������%؉<p6o��%����׹���!�p�3KM0�
��k7:���5�P�i�,c��uվ�7)*����J*+8��Kz����M��S���oʥ���rhL�.�
/z�ɨ����tS����Ys��ʊJ��/��U������X���rn�^���Y9���m���6�/�sߛL��4 ����-��m�L�D�؍1���dL�/sź��E�i��%��sϾ0\C�ݼ��)t�f��p��W�N��N�_�6�z�v�ǲ�m�RT%8F��d1
@Z���N@�C��<��
*��+ ��Ʋ+�,s8�Fe��u��֠��{���oi-������ ���cK�e�s0;�U%r��Y~�c���wNʞ�/��]��>�$�,Z)jK7�����!��%d���B���=Zk!2� {��
�K}^��#�w��1�ع��!�	��M0�i[}�����M�]�=�֞3ɷek��\��yqL�k�֏{�1s6�X/��(=)����T�?�;~��� �.�^sk<�����k����o���5����4���8\<w6�Y9����lۼ5���#o����֛o�}�I�~^�Y��s���j���O��?pee��7��~w���ߢ3���e�jo�;O����ې�,P�n¾I�t㪍����B�>s�Fi$9��(@ْ���Y(ry��D) Tѐ��*V	N�>}��ik���9@�=utx���Y3c���q�rܟ��'ׇg�{
��/�u���}e�C��}򙆹w���ߑ������F@u�]GH�Ѓe����
Wp�X�~��D>V�,���V�.�=�V)o#h��ve�Asz�v��;.#���VO^!�R��5�*�ev���s�*�|��#Q���s.��7!	�\B�ݨ(@^u?sYW)��H��}����*��[C�;^�?`(;2�Ej�ZY�)����Zk`3�cٚ _SEa�[uh<�^y��̀Lz�jR_	���l�x����ｵcf+^4�b�T��x��Jw6E�j�)"�!��I���H���%�[M!��A����tu�PQ�p�P��"�_:2���@�ۺ��-�jkc�'�}FD�M4��Ϩ��1��硳�& )8�l�rΆn4�2#�P9�� +����f���N|�A�����Z����5�/����c�G��[�3*�l(�"�<�c�Q��Z��
�y���'y,ȐW@y�����}gq�x�89�5̃Z c��+��j�+�'�h9�E7u���&��J�S��&�R�\�B�?s��qΛ�H�
;a�e�c�Q<����rs�Q�H�����Q&��L��N���K����*��&L��#,j.���n�S;�l޼���թ����+y��dx���1<d�CQH�b�����!1c�I%`�E�X����N��B�C䌽��Z�������{÷��� ��_�,�:����_f>��O������n�Ќ.M��frFx&�	9�,L���I}�JV(����*:�.c`w��>;�I[����E*�;
�G�`6`�,Q
D=8�w��i �����[a�ӈڈ�mH��Gxax�����H�M$������/h�r����ch�K���q��hﺧ�ʹ��;�M���C���<����:aޏ�ջ'T/7�)�
o��,�z��)k��O/��V�r÷���8���{��&/95�A����;��W�t�[�=|K#Ğp,�2�3�E�����lޏ�װ(��I2����$q,�0��≶��;��퐳�Vz6{�sf})�HU�Q��i�����;VT�)���zV�r_�m�5�|�xД{��\�9Y�;�-��5�qͦ����;�&]͘�Ik��X;wFO=��:	5��Ҡ��3���m���b�)\	���II�������|������#�.qx,��{`��B�����KȆ;����:�mP�=�ܬج�Z�k��B(�4���\f���i�g�i1Sn3��>�^�z@tn<��aF�{Nar���u�.��/ٸAʰW+'gs�F��1&��C�TaC�n�p6:��3.���L���~�B�s�Bh�ܪD1��$O�aC�J*f���Sm�״���	N�����`�������-'H�h�H�Q��ڴe;�Q6䖝��\;6�d�����9�$'���(�|����"d��$5�����e<���Y���s�s�����}������ӄ�(���tnnx��W	�����?��&�.ԯ��?~ix�w�	O������ �J�|�`��!�|��������ȼ�2������o/F�Eh���	<ѷQ���|���a?!�'{hx	p޷��x���x}�k_^��������!�g�PP_�i/TJD�lx��Ѵ��A��<(�D�<���f7�Z�y�҄U�;�����`>�z���+�0?����kg0�v ,���޿�����-�?Ex��a=�7o�J�����׿}lx��3����IJ��1���t#��2|��-��CJv� �{�!j��ʺ����l�z/�*0��.�i��h^���+҄�y�g]���\F��>�e*]�����U�w�v���qy��m��=�����_���0��ɽ��!��iŔX��*�g�L�I�|T�:��ngDo��*��,���cO(7LA ����L�-����
�7���2�43Ҡa�do5�X9���*>����.��1�#�w*�����c�Δ�
���(��(y�x�S�����u#/�H���;1u'�U@�6ne,6���}̋��$goy���D�\"�IO{֛�8�K:v1�����l	`�[C�����0;�%%��|N���VB���q
n#�"|�ee��T��s��n�o�4N��}�(,d�BA��B��7�?�gΖ�h���.��$Jgލi�**�S�;fH>��*QQI���JS����W�6�һ�s�� �;6Ӱ�~��� ��t�O�}�� ��S���5"B���{��d�����e1�6�/�{9�
T�?���҇��`Y����G���I8�}(˴���]�	y]�4����6}Y���~��5R��y�gZ�][�O�gi7��I�5��e����zp���'O�<�}��D�~�� ~aN����hs�h|��:��y����W>�	�{�ϟ~*|��P��C�z�_Ʃo~����3�������׿J��j��×�u�t���OS�n��[i�"���+��'ՠ�oC��v#\�n�����*S�V��a)�F%oEr;�i11ů��j���[i�J
��U�C����p��4�/,��8�>>ǜ\w�P<��~�3��=BNCQ��&�o��:q����/_^{��1;���'>9L������<|���&�����;��u\
�E#��ඡ
�B�F}k��؁m	Is/��C�*����[Ei刏B�WT*Qb�%f�h�4��Ϻ���<Vg��A��s>��5�G��{�}��lͻMN8�2؋;��ι~�f� 4��g�P�h��K>W��*(�t���7i�Sv��M��F���N�<Vs��f�M۽.�ȋ�߲���@v]���`��C���QR^�X������|�S䵷��x�Ց��YS���4�@�f�HsD�^y�d�-�����L�����h�w�>�޿�)xD�� Yv�ȡ#�,)7���J�-r0k���N��4沝��TJ�7��!c1ޗX��Ww�_�<�͔*�*K��E�%����OV�ц��#
�l#��� T�#��ɔ�n�H+(���n�e.�+������ G�T
� @1dS)�)������>���r��/ek���@����sj&o���j��-/�+��f(�Rи`��=�^�S�1�W��|��7J�f����8�T�#$~�6���D� ��qi�� �&����l�#�����(#�
^�)MKhl�1��!���o=;\#ל|j�w�xyç8fRֹ��'G�k�]X�[�>�uj6�ܰs���O>1|	������?��!���DAI�aLۗ�/������~��p󔶐���&�ٳ{/����>7�_��=�Cy	P�b�����q��˛f���n<���&�vָ���;����Nb�RY�~�#@��2r��a����G�R��'��/��
Į\h~FzW��G#'Dl4H+�A8rÖ|r�6S9����OcpyXtDS�x5���g]v���9�{�$nM�.��⇯s�*�'�)��uHe�Q�{��k��U1XX��x<ɋ�'#�(J�r��i.�[\��*$^{�{�U;^��]ڌ|:mu�m�T5D�S�֍Võ�=��yG�w��=���=g��yM#eP=T_)����~-Ui*K�vUBW�#?����9�ԭY0 �{����M���B/���D�zrƽ����7*��������7e��bP�0�qf���B�B�!�,-á��4���Lc�-��C�	\
�<4�����}��
��K�c���apY�D�^���w��Y�^m>36�9u�ʹ?~�RFJqSx��o"%6�!2������;����f��~�s7Zk[�j���4�,���8F�7:v'�/Ys��8]@JyS��<�Q�,H�ۿ�\����YңY���&r�	����#
���|�£�}��*��*@DJk!ZRȤd,Q�*�����"�'}�4MHT�+��ޒ�Mo�����: �;Գ��%0Ap����m�o���g|���BWc�R2r��?�5����ʖ�J��F�)ޣ���Ux<�8�G˻��}
�Ǉ�߆}o��"�ۻq���?5��'p��/��^y�h��\Ǥ��`� g-����5������_�M��p��O<����3/����3̓�Dy�dӪ8=���'?	(�������?��H4�x!`$n��/|���D��=��*_�	M��pFs����/�a����K0I���W^O��M;Q�S}���g��k�` vC�b�{�3�=��%��5� 4Ȱ}b|��]���r�c^���KYPи�`�\��B�"@� �m���z��.5c���??{��̰�0u�m��EVKM��FoX� ��
^�x�唧}�49������%l�;%�$��t"p�Kaj����Z�5�Df�hzs�����uݮ庽�^:V��jD�y��1���d�,�����X�ʯW��iT�=z�Q�1�/e_���纛U ]k�2���y}�d��yN��x�8˒�P޾{@�Jq4vY�8fW��j'�˪E��;x]���^?+���U��)�f@���Hd�7�(wٝ��3��������1��ˤ����CN�〔�km��,RW�� ���k 8�,�vd�:��r�W�4�#����W��)�$���� �F�ڏa�)p3�8V�6�x�-	p<��`F6���#ֲ�&��r�0rk¹���|�Q
�M��G?��,V�����V������hÅ���L�^,P�`��[���e�*`��L�Yeq��ꐕ\Yl=�[�7�Z>���d��]�]�v��+��9W����dfj��Ά�����+^�m���zhOm����%�o���{Q�����E�{}��a��yJƮ\�?4�`�l��U W�k*48�V:��M\������������_�2�.e���M	́X�n[�n׻+����<C�nF1S p;������O}�zqx���	�/��~����ç7a�+ઑ��6 d�]�0���!ex� �Js������n���3���dO����I��v��4���/����{��<���O�����!B�[	G?��G�9Q�O���[���7Ŕ/I��Z�f�J@ #Q[��Py�bD��۴�
bY0d��.g]��׻��-�}���[�����rO�5{�G��q�r�p��Aal��M�T�N�e2!�Jr$�IL�z�0�����9TZ�,��d�3��V�(�W!������cG��1c�q��{di�3����{޻ל�ptO�i���,t]9�Z �|נ͌T()��{�}?�Q�v���[}��GB���u��~n��̬ܽ^2�o�T;��%ru�a���e��5I���ܱ�h5*B�f�ٟ��ȇ82��Onwɓ�1e�t�\T�)�j���N(as{k�ȫ�p�}�O��g��_��p>�����0$V����0��j!{�X�l������ѵ4��l�Ȳ4���D���HS~��|��oڴ%�OβOg!O�M��F�w�$ߟ+.���H6���c���W�PɞCc�CcD�����������O6�8���LW�[��^��Rh%>|��|�Mn��6�����,�Iȭ�a�V*2�t��j�$����vd��^�Ql��h���]K'�ڣ�G�l����YU�����{n��[��p:d��*^Zh�����ߞ�����Kn�����S�~�l,�m�9�P6���L�?�ϦәD�o �d*ہ}��Ki�x/dQ(\��>K����DT�D��C�x'�5������}L�j?I����?�]� ��A�g�9��w�����Hd��2�Ԡ���2˲L�m��ݽ�����y>��!����!����r6�������N����	�x�)�H8�p�e괏2{���� h��Ƒ������0 'FJ�4R!�ܭ�w�a|(f�"^$�0K� [)�R���R%�#�L�b�p�"Q�׋���K/?p���y-��R�o+�����m�bZ~ @rT�����@�8;3I���x��`/��s�ɿ�]V�)�*]�4Ft����,&�b/C�{��Z+=��7Z�֑𣯅��s5�|������Y�^��D� �w�=�<�����n���8J��TB�_3Ҙ�nxS@�K�A� U[ Mf�H��	1)�,�P���c��M���W��F�E�P��H�e��oFs�[i�9�U�ՅLˑGV4i��r%���#�6�tM���/�f
f��4ڀ@i���_�Ѽ-�YZ��(�#d{��B`��d7�S��b��j�{��H�á|-�/FZ��rz��=�E�;���ߊ�p�Tur���HlAm).����;�q�y���>��F(�� d�<�nE�NK�Fk
=��'Xko���,e*r�Z�m��"����Je�w�����nm�x��{��L��4�&a��ΑQ�k+�_ @���,���r��3�	>�X��pC�Z�uWX~U���إ���W��A���,��a@��S�w~�\��q+=�������:!Ϋ�$b�Bmۻm�����@���8�>��SO��ng�(y�8\#�o�7g��T���WX��l�}Ζ��_&��kJ�1P�\�����F\��:(d�%�sM����kxBzG��������S����y3s��~���(�z�P3�5��o�Σ�o��������}�5�(p�+c�o bq�<HN��T��z	��e+FK�֣c3߆��θ����'�u�R�f*E�*ذs��fH"T��д�sK���V��9Zs�\]�^IB�K���~���Хh4����6���y-�N��A�G��h�7BT@�y��M�����4���AџV�Tŉж�ӛ�Q�Q��k�k͌���1��Z��w�(���W��AM��y���8V3 z���1G[�f�DqW� �y���M��g��k-������F/4g!�Z�q>}R���k��M��Wࠨ5]�-ͷ��w�D��0���.ӡL�Vg�B���n3���7۾�d�h�G�zW_�]�-i����/� ����\�e�bD& �MY�H٫&�F��^�c4�{�5�J���
H����JX�q�$�XL�F�ăhlIh�ꭽ���h�w�c�|�F����E1�n�W�IVI���r�<�����Չ�kz�g���V7�/
�5�*�qU�>��,!Q�����^���Œ1�����`��Z(�V�1�b/AW®tp=W�������P�7���W��v�,�n`�����u,Z�)�j:Q- �����t*�z�y�no=Y���V��B�668J�J�{�@�������yrŷ�w_��8�y�°o�V:��;��ß�8<���Æ7OR�}a�"%G���)��_*��AUT����#���$
}o�uq��+U`��{�@]7\N�8�1� _$��"����OϿ���6%p�xG���A=w��}-/��a��}���[�>�n�I����c������tx���4*Am��K)����t�7�����P��I�?׭"R΁�`v��׬���鑴2���/��EDs��R�ոEF�.&#9l��\i?��2f��1�k[�>l|�w3�o(�+����uޤ�d�&>��P�e���I��+ݨ�2��~p-��Y�]�n��+�5"�bZS���^6���Bm�*��Z	Z��U%�k�r׵_k�:�=��=�C��T����f;_|��xӉ��q�v���ȃc#;�	�(1XP�6x
q����T����T4��4X3n倗��tq��p٠�0<'0(g)oF���07Q_,�.=�U�s��}�Q
�	��t%�Y�s�*W#FP`䏴ՙS�42=V���-{~ɴ8�k����B�iRVz��z�[Eb�A��A���:���=̽	Pv���#�|��F�4b%��m��Z']�_K\�y�`D{|h�?�(�A�p�¾����J(����U�וe�hZ��nĳrsIo�7ls�ڂo�0�$��)�ڐz�E=�����WBYmA7�]�YRH��R^��C	��
p0�FEF���]`}������k��[j9��W��(󤫛�}��ckxK.z:��:�����@�z�Y�c+����sP���?�~�F��oP�{�wO>CD�<@:��#/��e�Ǵ>{^�u��A�H�R� �����0� o) ���,�FF>��:���0�K���5�}�.���s熟��-j��&m
��G �|����<|�;?޿���H�Ǭ~�����=�������䖆{���w�O;^|��A�+x���kdJ77mH���?=&<�m[��Iى�fl���&c�1��1�N���"�+ox����ɡkTVT`TL9�1�;���?;�ri5�ˋ����ֻ �_���3�o��ǳY�q'� $/ꞱQ�� Qj�uv�F� Mq����*5�5sՌq��c�� ��"���hSކB�Zc\b��y�M�3�Fo�(��騇������
�P]Ft�A��!:�Nb@��0���Q����+�����;�-�v�n��D&�b���c��x�7C|A�8&_�+�w��Cw-��߰�ְ�>�Da�k��_����4P_Uy����پ�+B�oZ�����^���Li��Lo�����,)Q���5b�'"7��E�卶r��br�_^_�����`.�!�S��9"Fc7���q�xЩ[̚:+���~��>��Z�B(��p�{`���b�]�eQ�ps����7�0OSB����S�mPJ�0su�*v-�n~�o�^NS sh"V�����r���{�̬��u��� X��skzkB�E.?`x���t+h�ս�
�l6�OE_���"�"�ۜ& -B�Q�[�Hoī=��Y��}��n�(y��7m�3����xi[���<���e����O�1?�Gw3�����Z�|h����.���Ru��H���X ?���K#�5!9м{{A�O�5�U��_���8����u�S���L8X�vmx���C�������ej�	0�a���?����6P�/Ѧu�?.�6���\�"s�l�P���Њ�6C}���č�6�g	�������3���-��F.HJ�m���0��1�.F�9H6�$�qb�R�i%�rM�#��՚�
&�chi^>��'�o|����֤o�y���i>��/�)8;�ɀ��P*x���۸k�(@r����ֱ�6m�B�:NK�-�=�qK"T
�x�}�y�zkͰ� r�}��>|�{�#K� �H�댏�.�{J�����Z7��
�%OAH��7��4�Ka��]�F��89^�	�3u ��7;��*�����t�6c��~�Ţ��;*_L�I�k?t+;D�+�4		Us���m0�h)m��&�`�J�d>8����������jAJE�`i�(j�O�)�N"�H���QĒ��{�7I�#(8�)�fd�as��%��TZ�����d&z�r�#������NOɵ:w��|2�Ӹ�Us��>�{����WW{��O��L�И�p�g"7ȡ��|Y�|�?�(�����w�^"jջ�/緹��[ُu5����ݤW4�PS�<�G4k:�Cڦ�=�Z�������
ǜ3j����\�.μ��)�%�)��P��(a��H7k�r��ꑚ;�L��c4De�ɱ)��y6E��|�k6�(�M�ӕ�L�	*��5�?��φ�|���w�X�tk�p+�q�\�o�{.�BnY�eYS�WDK�D������M �I�Ys=A�BW_+p� Ebz]9�-�f���Ǜ�J������Gh��5J�"��-j�W(��K�O~��c�.��[�(6����O=>��Ɖ�,�>�����̟��O鋾}x�����)5���Jr�Ǉ�jr� t��Y�7����	P��'{;�B��Ĺ���>�ܳe�����C�+��0�<vt8~��a���^hi�E�zvM��0L�p����*ty-�ZE*�Z����a��-D6q����箜N�x{�|��a0�-���D��wu��ؽ�S�ڷ��),q:Hv`c��Xi܆11{U�^(n��
/ 0=��ᦜ�k�M'O�L8W�R?}�T�M���|����Qڮ�"g�x���?�I¿<� ��s���pp�sϽ�0�QR�wD�믿��nݺ5���h�����p׍�k�-�U^�7kY3�{DN�g����O^���T��Y'��������"�Y�� �hr!	�+7�\���HY�8?��ui,�=����x�T�Ƅ�[E��v[��M
%
���,�&�j�c���\����Z�m��d��;!��u�[sN�������v��s=�o���r9�F����>����Ez�;f��I��m���3��Q
���|�H���,�&��̳��k륈*�X��QE�A���&˛��訁�5�o�x,�ֳǩ�#[Z����@��D��l)甴�+�yچݕw��&�=J�" �P��®m�{�N�مO�x����:
$Ta6�iE<ե���+KL����
�1��S'aJ{B��@����!��ߦVy�ҩ�F���ѐ�������oa��ڼ�w<��m�D��eYz���+�tF�ڔ��x�.02R��x�O�����&�G��Y����EǾx��o���J6��Ǐ'�y;���ԑ�0����dmMM6".�;��WQ
;BV��<>|鳟`�@��]B��޻cx�8�;ߝ���mU7��^�u�R����������D�.s=�9���Y�k����3?�i���=�P�׸S�����u=/��Y�H#fC�����g�n�Y_}��ч�J�s�>.�՞=}�����X�>��0	(K�ۀ CzR	��^	Zy�6�֡����8�d���]�az3�t�Wٛz�-�j��������E'q�w_�;��RN�V�c��2��u�.�s�N��e<�t��[W�
���n��C䣑,�׈R�������th$��)�s��w����5Ǣ����n�d�k�l@�[����u/�YN�c���4~3d�|�HP�5.sa�,ƹ8�>k]<	 ��q)��7O���NP`�]=ٙ��ФB�M;.Q_,1��;�b.|�9?A���E�u׉�ۗ�"or+_-�#"
����7�y���m5�E�y�R�	�s}�ō:Ǣ7���������)�ߌ������b�{u�yO���f[�G�G�"-�̄�*�R�]��?����-�PqLJ�E����b�sk�6�w�m�,��!G��hf@��E�x��He����;�vi�֕z��=G��5�ۯ�[�]��r�CzG���a{ CQ%ږ��Q��Lo�7���K����X�1�l3��%0v	$���[ J9t�p��֣L�ʑ���OT@a��nº��Z�56�w6�f��κ	n�v���@�V��!�P��[rd�:щ2F�'ᮢ������w߻��Z��G��v#H�3����G�G!��Ƌ�H��g��0Ϟ� �qc(�O|�I��_�X>9���?�yܲ}3����ȁ�a��㞓���4�x�����&�������{�� ~/�~�\�|��utػ�� �u\�E:D]&Up2i4���WV���R���\��7�.�����v@ͻ�Qy�'1�0��>gc!C�*o@�!�HJ�K���>�������d
L�������7m��22�,
}�*VE �U��M	(ح��*^��h�}MaV�qC�O<N��S�վ\�ߋ�+u�`|��ƙ���>�����;�9k������a������~�ϩ�ϝ;/^%�7B��o�K�����k�Nq�`bTX#Fzɯ
�&K:um셖W~X+}�y�?¸��`r�(�h=�uܖz�*6Z��rH4,��hY��)��')#[G�xU��O(����4�m�j�lU�d�w@/����xOw��b����u�8e#�F<����\~�Y��^��R�e�{���:_��r\?�f�7���@7�˾�~P���b�5���<��&�1E�%F�-Ѣy҇F��N~~�(t��A�����C�`o�23�_)��������-?�-�t:`�OdϗE6�A�BUڝ9�+��~o7���X�t����[�\�fh��.��j�����G<u�Ӆ[`Q����Y�e�S롗�\��uޢ���cu���R��R3�M��X�����*����ϧ����3�����n�ӛPN*_r�7�H'�/me��3wo�ܚQ���ث"���|<����]E*T�=ק������X�Ȉ�9k�y���G?�E��c�ޖ������5��o|�f-W��	?h���O<pװ�<�>j�=������H�����?HJ`#B�����	Ť�FB̀t4��[]�rz�z��p���BV�-_���	�TLw�&�?	�����j�f1n��矘Vi ��^�0!Wю	<�� �륺E`	��)��P�\���(����]����"`@�W`�KȚs^����>7��?�ï�G�,v�����l
������k�,4�[�(�+b#%l�W��j9ZX!N�x��jM�h��o��/�˽���z<�*����D>����Hw��um�u�}���������<J��~뷆�{��5���=�\�̿�G�1u�Y;eT9^�D7N>�[h�Q�牆Q��׈�l"Jt��=7���`+��HMzz�&%ʙ�����^ެ�짢�6���\��S>_sQ?��R������
sת)'c$"�h�^�~�sJ�Ǹ���_���Q�5e��i9������`oND��k=W��{.>��J���%�<��C:��l�Į���Y��O#���1��"w�BG�����K��e�,�n�L�h�Η����N9�A����hH��7y�7�z<�B����⡶ܕ�7���zۅ�A@?_)��L��(�����{��|�Ub���J�F[s�6�\�޽{�ε��9(�N�2�GE�G�ExՄ�IU�Q����O�a�!�^��׭ �Q"�c4���h�U[�҈}�r��hQ��]�|Kr���n��j��X���P(�Z�ʖ�©zo��?IL�f3���ն��ݸe����?�~��p��{���vv�P��Aj���u�	�k�b��رe��8m��:���Ƭ�׳J>Snup�[�D`vflطs˰o�f������O%�`��+���a��)��
�NB�I�����@t@�#�m�r0�bL_d� B=|�
�4�m\�ᚖ���5ap�5||��}ۇ9ش�	�?��/�0�{�]�wP���p����UfZ�Mo�l��1�!����o�*8�C�Ғ��ٸ=�n���es�0r��b��5o2
Y��t�o��o���
炈�n�t�rޖ͙G7'���`���o��o�*ٵ���?�����?�T�a~=��Q0:0���[��%T�;����[��U �*���v(c:���%�l��:t0-|Oѫ�ƕ����$�U��dHV�.���&{]㹸�E��{"�R�떉h�����1�k��g\h�)�M��7W���9+�E�O��<R�˿Tx�^_�)c�>��wߥ��,�Q��-]�ܑ�^@l�܂����¹T�K�Vi��{�E��ږ��MD�<�x���8r�k�q'>�c:��Bbw��)������n�(,חs3��Qd���@�6!��(�f�^���	�7?� 5��\�:���u�fH�FF7��*�\�n�[��d� l�Xs�������������C�>	���m�;�+�*���Ϝ�w�guғ�vh�T
���~���'A�ޤ�ZZ��Dy߲Fk�l�[xL�+�&���8����ǌ���� ��:V(��,���Av^��f��{�}��-�#J��-��*��E���ί�Xfvf?Cx{nx��w��(�x��C4��v� �
����1_�{�-+�w��&*s�#`��K���]��jt��� �e
C��m�Ƕ��nڻ~�Ệ};T���/P����7��4���)_�F���(X��߂���D1�W���q|�!bDJ�_&��2O�h�Gț������͖?��<�;��&"�v;�A�s�P�����l���l���VCv��102�����4
�̈��s_ۣ�tv6�{�n�s��\� @��5�mKW���p(%��8M�َk�4��w�}�N���[���{�{«�?
�Ν;#+zw8C�K���.�F�Y��?���i,}0��(^ߟ=��>
(�s�1�F�~��50T����A������ʐ���"/·�S��(c���Y��g��M��ɦu�T�>�3�7���,�ri^w*���_��x�m�� *bX��jV5Wt_�۔��ټ�;4����=(��d<�eqe�z]��G�s��_E���˟�RZ�c��M��P��j�@��k���+�j<��C����Z�����(�UWmu�nҮ�no
��z�j�`S�0����o�Q��?������=?߅A���[�Џ;*$Fa?F7t��)4քb	I��
�E��+]"�4���l�?�Nݻc�p�&%�+�l����T��p��p���6Qص}�p� yG6�['N��C#�'�v��ݥid�5�= �>K�Q;��Ү�iK���3�"n�f��m⡇ڻ���Y�	��Q,�9E���H
�����?����fw�!�p}8rx�p�й�����I�[��u<C��i��ѷ	S_B�V7�!���Z�	[5� �	�z߈
��K�9�V�o-O�s`����y�Y�֍�$>S(���w�������h�s�:Áh�ٍJ�gO=;����*�-n���]KNr{~8�o�h�V)����R���hN�q;Ƚ�o��<h#�P^�B5C[�M ����nb45�Ԓ�7H��A�T��9�Q���}�����]�T�ɏ�Z��5:�#���jѺ����U�7h���p��)�	|=��6�ƹ��5Q�ʖ.�R��?y������G��tע�9j�e�uv��0j�����Q��R�DalK@��t������������.>�{�	�d�e��l���c�(?J;K��Yq�s ^���2�Q���V�S��R§-1*ڢ-����P��{��Q���ɾ̚)o=�ʳ22Jn�����7�F>;5yss�`}֑4NZ$4��KK��~�:��FD����M5�e�o��T	P�:��:���Awd��Nnl�P[J�>(����f��bM�M�׶�*���2эW�j�u�}5��2J�t��c�V3 |>z]=?���2����qG��hnԋ��O������W���%D���
�`������,ex��������J���ײ�������˿���w~���� l2=��~{��o=�]���KU8��Q��Vm��Sl"Ѹ�2���u�g��R�+�2�e�!lJ$�$}Y�e�7��&2j]��O�y��̰�u�R�g^<6������ �]'�2���a���U�<l#��H�۳-�����7#`,����\C��S�fl���5���MYP�w�OOu���Mݲ�ĺ�nnӖ���
���;��T��47L��4|����7�7�^�N?:��ҋ��I`��q�,:���j�eв���MflU�����O~�>��)�C�.���#�:Rh�_>���s����Q��_��Gk/vƶ5�u��{4rE��NCjd(մA�����d4�N�@�����U������|���'w�a�
�P{7��LH9*�ei��h��}ͰY��O9��%� jE�a�8���=4$� S��S�yLgC޳\O<O��k}���>c?a�1*T���S�ҫ=��R��3|:֞K�����q�K�b��V$A���K��h��8$�d�ƃ����g���Ջ�,2^��@DO��i
��Ƚ��R��d���ߺ��z��0Y��qݻ/m���w��_���;��W)��_����C���L�R�n�[�]Q�z��F��׭ U���J_�i7\�!�������������z��������]P�U!�l��F=�n��ޛ�x�_�����֊h�f����7���~�f&o�?�c�y-�pѐ-�mt�?�����������~틠�g��{�G�Y��K��rnzۅl����zЅ���0�n�Ox�����"5TQ؊��n	�dZ[}V��۱j�Z���;Ǉ�����S�%�?��q������B/G�F�eI�U��%� ��s~��ru���DX�&�]�(��0Sy�#��m��=ÉS硚}���	�n�p��$��Mx�� eYi]���ؘ����ר�>2|ꓟv��7��޻��edx-���]x�@�Mn�h��ER"0��ّm��i<�bP�%|�s��\�
�����Djv��5|�����/��] �9�� �u�q�GgyT�}�;U�s{29��k�㬳.���`8�!�3\Iʱn5jԍ����L�ݣG�����T�e�B[�6���~�%�Ͼ՛cz�/[�4O�����p��<��0���v�}o�W4|������0o�1�u�U�ݵl��q��y܃g��Z�Y������:|	x��c���V�o��&T��S�T��Ζ�aٮ�ͫ0�t��7��=g՘e~,]c���2p�|��j��viʚ�&8���2��`+�:��o8�(\��/�<ɽQ����i;;��v�Yw��W�{*X�`�}1@[YH�K�z�,�K���[E�D6�aKl/�7�Ք��z�j��D��|���FI�T.#�&'�n2oW�����
<�+}�����66��h����G�ص!��e�<i�[ϑu��n���\{x������u�н�Qo9ۢy>�!����u�r4��?߿�?3������y,�;���>:< %�|��ָ��7!��I��Y��4�_��}cQ+�(�ϧ��A��A������g��9rǗL�aL37E�^gдQ��Jd�t��x[n{�h�Bj��#X�Ӷ��筀!�܎������/\{�rϗ�^@#��]���G}����3x��gO��6d=9��1�vQ��q�x* .]�Fkǭ4����>���G���0 �zr���_��_�{�[���l��ȯ�n}�|������5v���/V.#�P�x��	��^v/�)*�)��~�4��8�,\ ��ֽ���wx�����Fʤ7�x	e!�(z5�Rd"�-{��-����������`�_g�N�-0��ݲ�~LĲ���!�[�W��<�����YC�b2�77��R��&J$X�2���Ͼg�am:]7���={�D�-A'|��6JU�7��{s�/��O~�c<����U����Z�����h�L���{��dS�9��FJ�D�[�nOo�/�6��r*[\g(m���c�ZY���!�j!�!S�1�A �Mz!\��L4a� ����.���>֣t�`���q��8�[�}�S�(�µ�b�����W���0�;%�ڸ�fƎ%о��{>y���{��'�
�b��$B#Xͮj��=�W�N��p2��T�{D'}��g�y^)��}L�J0j�Q�u�C�lE�-n�*��s�Z(�K#V`�b�/I��O�$`\��K81���nxY����e���W�%�u}G(tۦ�����)i(�`X�G�3d���p��mH�q#�k�)��q-��J��(b�U�������!�
�U\�{��~��*Pםm�wME�4�+��Χ�{�l4"0���itO��u�~?�u�
y�g��� �����4j��};�6kmA_o$7ڕg��k1�/�?��	�mg�Y�0�-<�}j|K�Wc�r��k�f-��u衏�ٞ��Q-�^��R.����̡�b�\}B+k�}��gs'���_p�J~Ae�W�P��Ye4~�^J����C�!���}N�7���� l*���ܗ�����-�6�x�
����ϜZ�z�9x�Y��?��? Ran�B�Ρ��x������K/��f	O��h�������3燧�r��q�|v�ҳI�#Nuy��I;�N�7}��(=t�$����~�l����r� �T��������0�M&�z��^"Mq�:w��BC�Ϟk7H����W]ʲB1T���	o��.���7��K/z~~nx���
{۶�	���1�~5��~����)s٘��U�~�*ts�c�4��E�\�.�B_�1�s������J���eª��F�Ч�;ʯ[�GTN����P�>������˯�!��ڸ��&���	/���L�A�u�^5�S�1S"��+G��[�i�Ҕ��<v6I�t��������c�����Ki�깍�X��PІ���(t�m�l�����95�7p�(e��C0C�IbR�s�wf�C����vu�u&#�^�F��Zf�<��g�o९g�\.3f�Sx�IePwʫ��
�
<�����9~���ϟߨ��W)�:�5�����ە�h.�a}�?�P�h���g�
�!��P>k;��Yx�y�	�y"�JД ����Q�|�����Vs~�/��[YJ�H4zz�$��$f1̥�+�3��Ր���n����.��n۾u�qe���Lʦ�)�m�"�6�%��%��"�eU�G��_�R�.4�35�\�p3筷" ���3�
���}��/������o�XZێ}��׋�d�#�!
>���.<�i`�1�۟ky�8�xN�t��7��<��ؐǈx��L�2�L�����U�����+�Ϝ{�p�L�4�
${���\�vO�R�#=����÷����ЃSQd��W�-�ҵE�f��\�K 	�- )>���&A-"#�8��+ MF��\��@�� fn��	x���o�8;��{�~�Y�^ZAK�ת�|�y�-��x�`=e\���Py�Z�G�X"(F��[��]�"���{4*�\��[�p�H�ji�� �����0���zr����o{I"���/�"�z��1 F���{�ˈ9���fa�#���:���>j�/�e^r��ި��� S�f]C��a_u����7��ؓT�\�L�����:�'��� �Z�U΁�[G�r��|U Ďu�TY+�3U��s����cgiժw��hߖS�G҂��F?���-Nf�m`G�Kl���<N�b�A��9��t׺ڻ�tuH�0<�o��P��x6*bT�e��F@����i~��կ�Ɨ�O��S`}ڍ��w�9� Cy4¨H�6.cD�n�4RH4��'Bb�"�X�������kyF]������:g�'���M-� "W��kn�
�S��H��g�w䆫�N)뎦�������9�������tEdv)�B��
ܩE�r)~�gz�����[5� �'B�m��=7���ٗ�W���|��# �����h���$U�;���c��8�Y�Gp�q?�!j�F��"F�X��n����-� ��Ƚ%�g�K��X	���E���6kg����S�4%�ؑG^���N/�OaE�M�VC�K��ϡlqu�Z!��,
\����4�Y���5�w�|���뷇̈́z�Onx ��ÃG?��χ��.��we��{_��'���C����e^�c�Bs��q��<�Y�C��Q%f8���&Ü+�k��p���$��s�
��̪���5�m����Fhĺ����FV��S��UE&�󺥝���Z�Q�%�/Ɣ���\r���4���6"J{U���1b�=��=�M[*Iic�y�2�z�E�\���ź��H?��b>�A��^�ىiV�U�K�m8����#G���q���s�o�k��~�����);���� ���AJwV`�MZ����1p?��G�@gv#@8A_l������@E��-�@�#b�ޔ�:+ݬ�D۲t�����{8���$R���/%��������n8�u:+J�s�Ȝ���r�*��0 p2�eK_�A�ԛ�"��DO\���s���%�$g2u���Έ�ն8�~��ᕗ^.\<Gl��я�����9�{y��+�n!@f>eD,?�#��A��PC����x�:��>�;Fi�y�,��iQx�uZ+)�BGi���&,�x�=��Ӈ�o����[�a����5�[m�(�4�(��[��t/�pV	ʘ~��F" �e�5���g~�_�j��ЮA���m�K�ݕ7%p��z_��X��{/Jo'!M�va�i�B���h��W��f�d���
�*�� �s�P�5끱�R>R@!ˢ�VƉ�R��z���������1>ڕ��X�e�!AS���>�я �"׆!���/j#���u�� ��x���ُ>B,<�y��:Ы[��	ᎍBlbry8t׮᭷^O>w�P�ۇ�ss���9̢h�y���"�˒�,"X��?@�pWB��6�nϽ���U_{�V���r꺩B�u�R��88o奲��b�s�r5*`O���4� ���jc�w�][�s�<���Lx梢XkzA漛Kx^(��2iq*𫕒i����(�n
��"�[��*�[��]!�G��M[�q\]�=�$��6ڞHڠ�ٟ�Ǽ�N �T9�� _Ŝ8$����a��k1*/{$��w��.��[5�c,U4n��&��c���Ű9���b���H�l�Yˆ�3�w��1�sx���a����ṗ_.B�,�KQQ����h�u���������2����pP�e��[���#��]�"E,
r�����3��.^=���f�y�sMkh] �r	�}9�O�:�{�N4`�u`EMR��e���s	�s��ft�"N�k�6���d��w��sx�q����k��Q���X C�n���އy�%�o9�Ir+����" J�s�$���#��#��s6֮��>��? ț ��Qm�+�nߊ����mu�eE�T�������2�f'kg���s�)��ZM�T{�s=�f����f��hRX9���w�C/�G�lZ]l_���`�z��)���]��N�"̇Ww��S�}�P��m8�Ojbϱ)i\!��_i��uz$��m�w�Ǻ�j_� ��|Z���Sc�T��<�֌"�o�aT`¹*C,�临s�2T�;9~�A�y��(���T��76�g�n����<;<	����=4D�~d?�����˶m;#��1_����������7�7���ςt�}��hn��j��n�lټ�\9�0xЏ?~������6�˞@���`��W�ܕ2�J�Nzz']�ҧ�J,�r��kߑq��Z�QGO $�)�Є⽄���4ү<���j�-�g��|`��S�	��.n�ǐmt=KD����mD2����������2�cIQz4�\�%��'/\Q��T?O��O��ؕc�p���MŰm��TYx�}Ҵ�����/�@�6�`�Ɯ�4�*c1'��� �^P�*}���R|�׹�{w����~ޭ��HKk�RX������z�}��5xMFcV?��3�e�]!�}��9s������!R7FgX��bd�}����P����#=�Q�PK�V�T帷���I�"j�G���������0�)��m�bӤ�Rk������笖G�B�e1��+�רܸ|�"J�<ǆ����({@��V�H*�5���U�P,eX j��Y���,��")�i�?�#�����"7xq+�RX6:�����Snq?D��%��kb�Zl��N�uG(�3g�<�BO���+�����z�iS��6⡛�r+&�Y��*�X��+���9�icu!��fߕ�6��c���s���Lj#զ�{���;�4��{�B�!�<��z��Mx�?J3���B���`���Xʆ�@�^Z��� ��g7lb���>	��1Pۻ��n�]-����t�76�̆1:�m�x�}V�8%<����j��eNeP��7� ��5�F7�F��品)��Q݋��Nݓ�ס@�GP?���^Ν;3�w�����'N�&���]Ò�I�Ɵ}����[��O�n���$�~�zB����p��"����'��>|/��pE�;}�8��ΟG��$��j��'������������"�ERQZ��Ly��1�w*ʤ'cX���
zh�y^��}��s2��642.
�r������n��H�R�Q�#�L  ׬�_On}3�Ķm;�Ӕ�A�*P�9ī#^ߖWh���:sN���(`�����|��.i��uDy!�ס�r�
��`���a��O�� ���} �>ɹn���3�=֌Q�������W^ɱ��և�MYT�2��L�YI���=��B�Y��+�h�NX-Ӎ��ze���.v�,��9���,l-w������NA&$���mɟ�h*��>����6��������SI�ŕ�
['"�ܽS2$��Wբ2Ճ�ܠ7�R��:a�ײ4s~�,�n��>�T��l��c��2�������w�?���`"(�q��u��
Q�MD��Ll�>���?}���J"u��@���J�	4���A�,�X��LDjy��Z|�9� ;��&;R7��R�"���
�f,��_�˻��|U��M�W��G|���"��;Z�Z�Z��_�Th���Clk��&t�'\@���� "@ݿ�6��iJJ�VK�l9MYp�������[��ZN��H�.��������^}�J	��sӊp�w��Ʊ�o_%4��{�j|���sj8v�,�׭��]0�ɾ�&�j-��]z`�|�:���p��C!����r���gtUEZ!��t@�E!��ߚ�^5�F���Uom��ֆ��`UI2V�Q΄w��a�޻�m�ۆ?����e��D��$>t� ���{|����\,��#�5���mG�T�voR�2S9**s�zW��%���T�m���9"�����3���֕F��X��EB��[��x�έ�h/�r.}�υ�Ӛer�1gT���w�x�25N��c���i�#+[^���3ˏT 7m8�o�q�hog=�{�ܮ�q7�*���LM�[e�rDs�^\v���Q���C��*�E��8[ޫƶ�c�N�I��(�E�]o[e�O��=�r(t{֠;F}�o9�=��g?[�|�zT�6e�����!�M��j��e^�zu��!2���Ip�U��~�a���I�b��2I�<��"(|���x�W�ȉ�B����4�=},J�,�5���ƧX�V���$� ��S�Q�� �Z��i��0R!�q����
���-��#wz*����T���62�<�D5cD�1;IYޖ����w�� w�p���ͷ���b����ڹ;�����4.+��!geEpB�Ş���T2��NX�Ls�� �R����H9.r���k���<P�S�3ރ Ks��J@�EZ�s�W���\�!�p�v�U�����T��S��p�:�E)X��	���������?�R�ցy�]q��v/~.LX-�չ��ZW1'�Y�OO�ŞZ���.G=��Ʃ�o�p�I-ߚGIlH�j�Q�P�r�����OH��
���m�=KxT�Q$2�ݦ��p���]�B��j�8B�{HZ��RA/}\����\�%4���!�Ǫ��{+߷�ښѓ�ݷ�9Of�a��C�G��|�r������e��SAn_��֕݋x	�	��MO�p߹D'�˷��4O�>B������w�'�Ͻ'���V���5t�|T
ȉ25�D)oU��"ԩ5|e�c�f�_�����.�w�����w�Ee 9jR�_�.zzZ�=�6󻛶�2�۶��Hv�|�k7�����w���
k#T�՛ẁ�Q1w�������?�P���u �RV�[���M�Q�_�җ��=?����~Ơ�4�/�9����>|�p�ǽ����tf;x�`�D�خ�͛[�.�1<�q�FdMS��=�X**rRh}��B�:�A�Q�������	�)�8K>)�Ҡ�-�-�#�|�=*Q�'Ξ��Q� Ϊ¡yԆ֙v#oF�R�b/��G�?E��<)�E��b�~���ĳ s�DU�H�sF2�m�3��2zȻ��dcM{)���~���(w90h^�yv���C�'N�����~�I6��(H�(�m�Ml�_
�N����)���%ݓh�t�|���d6��	@��k�~Y�Ub�s���{�֠�����]X����M��4d��js����J���>���-g���u^�|���Ek{�cv
��q6���Z���%\`Z˱��܅�����GN�*�	���b���Q�w�y+��'��cTN�SNzIn��`�?/�{7��� �*�����ق�ۏ�|=J`7V��,K����+g�#�n��y��"��*��P�lS�b��5���ꡊM���/��z8׹�z�l�h�.+x��H�iSr�0=z���g?�	�k�W��5�x��g�W�=?� t�G��ko�z��p���{�`k����t�b����x�g�_z�<��tM�Rr4C�6y�n�jX�s���6�R��������E}Ҕz�K�oW��QЈM;��s�Ʃ�1k�v�X��2���:��N�J	�]�S.��u>���}���Í �(9�[O�\�PS �����Q�=e��K��<���<W�T���1 O�	B�c�NA �kV��P��+�����%j���y�Uu�4?A��iM��H�ֽ˦<��?��ᩧ��5\�ç>���պA�z!���hL�^^�u�΅����a����^KeI�,�3�l�����N���9�V��S��%4Gj̞ ���l.�����������s��"SOz���sou�խ�4~���';����3,ş�531��͉�S!�l{?�:�G����4JR'Kz�Bn%�������)Р���|2\�0g��L�X�
嬍Y:�>���wh��j�@�9
ގ�\�ԯ�������3_���Q���L�y�kJv��tp�K���7��%]����Q����2����1�k�rh=̷F@SԅO�jJ��(j�`?�r��s�uW�w��\q]W�C���̾���&�^��l��ּ�|�+Jx��a�u*�q�P��7<{�w��ل��|d����?�DاކDe^�V��%������/㼜<���l��cg����.�R�J�"�f����@�������.��rk��5���RM(s#@:��gl&�2?�2�ַ~2��HD��������>w�(E�ɻ����S�����a�7�z�?x�p`��E9\%���5�	#����s����mÏir�}a~p(tǡ�=z��p�<@'�����H�2�����DzJ�V����?uo}���+�[�~M��sX��G)FaS6��1�Z2�Ud#�'���[�����Uۇ	������a<���!��#��5��ZR��/���`ޗ�(u����hz���l�F�D��D9��Vqv,L�Q��7����}��P��ӷ��}�N�{=�֍��Y��Z7J���~4�ѽ��.���2�O/k���p���|yf3�݁~�z[N�oi��@b(��jD�d2dD2�m���G0'gUWA���V��-E�<Y���JmY9!�����U�1J1�E�}e�16*���f �����LJ���X�_|��U�֣�+��\UfDC�� M]W��?�U2�j�Ү��q�05YkVT�ڒ��r�D)��"2�1q̲8�kʥ�C
����%���1" �_~u�:s�{k���4���Rv���x{�΍����B1��{μ�����Bq5�ߔa?��@��m�c���7a�l�2`�r�.�)��'�7?eN� ��eyf�g����-Q[���e\ʡ{�i��Z�Bp�!@��\si���;Gy�g���������3}���w�����?����g�C�JJr3�M�lm�I)'�����o��mO�|�������αТ����FěWQGn� ^ۘ%l�l¯{D}�z�aU�	����|;f̬��lt��E>���ڸ�p��~�0A[��k7�M��ax 2Y|��q�����;H�ov�����(��D*���P�|�^��%�!������a�{�O�3��#��y�ҕ��#`�� ������M���C��t*]�z�5�N)�R�k���|�s�:C�d�B�ѕj���gZ�b�lhpp�S �'	�&="�&�=�z�!;�ځO��2(rrג
͐�zz����i5)3��l���Rr�%��='ajäajc�̑�z�5C��My�֋w������W� ��a��n��+��݇rè]�&-`w<��xe����R-"�>K�u}�G����&L�x~��Mi�B	I����Y�&�{ɩpP�7q.I9��Xq2����3i����8��FA��|��� ʕ����6\�Y�ab�=�r�4�̌M�4o���Zn�Βk����S��=���P��X���
4Jf ����Mos�+�{����>M����|hЅ�^
�nql��`��0�}�m�tם�l�,��$ę���'�vX]���o�B��c`�MZ��������/S�<�R����J�B�6r卺�ݰNg��G��g���͔������&A7á�[9�`�����л���aʛ�`p3&Z���T_{��J�Ɖ�w�6M/�®�:W'�螺���Z
���w�4c��P����_�����������=>|�?�\dr؎�����j	��畅��̮�����aw�:�����Q
��Q�S�Ү=����5OsT��6��hj�CeT�y��U,�\=�Z+FSd�ByM"<�Pq��e�wx��O�tt�D�r�z�1�x��i��w���"B�'?{a�v�2�y�>x�o���#�w����e��+����|�QhUOsN���<��ZO��}D�����T_Ö%�Ǩ�^स-YJ՛y�<b�A__�%��fx緓"���K-��#���	�p��В���Si�{^��4+��y�*k�G��ʡ���1��쑶=���(��U�A�Ⱦ���s��#�9Rk��!�,���wc�˓��F���B�G�=�vT��T������'(���xW��37�!;�C���b�B��?�1�/~k��_���p�VV�+��m�R��:�*W/��]阤ɍ��5�������FZ#@2�+�A�e8�H78��
Y��5ra���o���Qn��D�lq�8����F�d���H������4�����9m�i�|r�e~OM�&�1�4��9ڬ�f^���0�:=9}}���DP~exܝ���
e>��:!�C�yB�YL�lkU#�_�X.��̟�O��B�k�. ���7��A[�ϒ~=t7z�\����~U}v1m����ũ�f��"J=�t��P�
��W��r�����x/��&XFQ�U�ܬ!~Yb�P[��區��|s��?q�������+Ã�߃��cSA*�y���G��Ͼ���ir�z2vW��(�'�9�#_�|����kx�����}�P�lKK��tn��ix�]�����G�B�Ѧ�� ��Yb�MJ�e�s�?Ԗ͛�d�w�����A�� H��x�s���_��_����Q��>�7Ets�"���ӝ��Y�ǆ��憓��"�0v8�5���Lo;b��A���|fEՍ����u��o4\���w[Qh#z�q�أj}mEV��0#5n~�~�)+���D��>�:_?W�f�W1���s�����Q��ڃ�Ǩ��s5e\�R�JԆ{L�Q~w�܍�j������xu�=A��``��J>���*`���.8�{2J�Bc�K4�Y�N_��
�<�x��u��*����Q����\���$��k*��eO,�[��0��<�g)��~��P=	L��d��r���.�yE�:t'�����a��&92���&�����+
ԁ���/1?�5��SsD���O���C��Y��>�(�]>�k ����=`�1X0S$".��O�y��*+34x
�D����إ�2cB-�T֍��+�:5��6���y,*:�Oڕ��W�K�B/^�*�"Y����	��ԡ6y����jFC����\3&�<���,%t��6r���Wy�������ǝ�SǪ�e�{�J)���+d֭i�k���6�߽:/,��D5�p,�1�h�в�G} ����
ݟ �	�:t��a��Y��o�V��h4�%o���������α������^ĳ�D��B�(:�����w���|h�tZ�>�m����{,��ͨ��4�J���LِR0�~�k�~;y�4΀|�N��������ʅ��RΡ��"�,��kO�v�5�H�iD;l�=��sk��m�<u�*y�R������6K���z���Rxױ��ڐD�`1�T�� U�5�1��)���T�.LyFx��(�}��#����"�%V�@��:��.�hĪ<슆%E�wM��>�����hV)�5,@E�T�������wϹ{�l&���D���kc�#{�{�m
3�>�a5kꑀ(�6c)!m�be�+��5KT뽢�'���-O�I�����>�;~���ʔ�a]z{��M)\�5��	'��x�z���`��yd����j2F٤�d*3s\Q��COz=�����b��{����s5��<s}������*״]�i��9�U�)sl�<�/]Μ� ���p�'Z2V:�#+E6��+e'@�h���z��8��}��Np4�Q�Sj{���9��^��˝���x�n��iEq�t�*I���Vo�O˥��9e@n|>iɚ���R������*���??�������y'e)�.��F$k)�ch�f	��{k�i	l_QTA '�)y����%)�>���zt�����P
b��
\����b�,ky����Ob�9��ޠ��n�P�`�+;}�t��NQʶ�4�y��%�X3��07"�� �>j8F�>D��=F*`�UJ��=�]Uޣ�է�r轼�MY��T<	W�sm��n I��6֓yS�Ҩ�UFEnb���ю�.ӣٶ�-L��z:��h^B����*%��=�F���t�����Ի��^m�_OuYԾߌ��F#k�"Z.�>>�H`�%Kr�w�Do�K�(��<���h���HS��Q�az|�h��K0�k�w�olM��e�c�T���b�O��t�X�{�Ae��Ux�GBۮ$�K�޶�✶�(�`�ۢ����ާ��{����!�ƷzZ�_�&!�Am�"����?��9����
�������Mb�t����hY����5���3g����F5�VQ)SqQmkժ	�JG��3:�	��Gj)_ݏ䶎�bo�1R����V]E�z0m�۞���H�^k4K�p�f���@�V�kx�ļ��M�7=&��Zr�L�\�``߀��=\�z����.ڤH����Fjh�T�����o�B�r��y�ڟ��i��.&�֖z�i|���bv;s��Y�-$������.8������~yM�Dh�Φh�7�p��>���)!ַI���ؾ[a�zV��UY��e����QF�E�W�~�1�u�q��b���1��w?����~E.��5���m�ַ�v.K�9�?NC��I�S@U[6A�I.+�AE�f#�E�P��@@��(3 z���5��:>#-��������f<y�2�����;k{oFa5χk�h����H0�P��@��WB�z�M�I��egT�el\�u��=�Tv�J�ܐ{u�?&��T 7��+���y[3��B�z�.�&l�zZ�Vk�4��¡|�cN
cQM^<τh`��1��5���m*m�6�I;;c~ݨԜ��6;��S
��H3>�;����^݃	�Σ{��*m+��P1���]%\��|u��XZ��?�Ԅ��	����)�B����	�O�������
�I�*���zծ�%<r��_#�B����^7��:��m<*���)'t�Z�Жr}�9��w��-��.��B�1� ��K��\L�u�q",R-��^q�'�@e�"_*_���a�X��,�+�a����^���WC�d�bn�P;�1oB�{��9N�H)��a�^��%d
�G�;M=9Y]v�>*�	]Y?�IOl05��b�!(}o��톗���Nw�A)�p!��۸@���L�R���
�Eu���ѣ�=��#�v�%�-K���^8�'�Sea*����j�Py5��l�2˴=��%dz(�^[n��[vUx&�[���E4���j0DpU�U���m(Y��R��$���u�Ⱥ�ٮJ�U=p]S�ڇÐu�Eh☨���_^���\d����,M*u�^�C�bG%�)��^}���|�M&$@�R`��{;J����	��̦�k��Μ;�/�yj�}P�NTh�<��S.����",9�"�Uw]���ސȩ6h^o�n���d�&8Q:�!�Lad����g���K8��)�*"o��pl��W�Q�"z5����A�./�6�h�7�h�ʻ���O�Ys?m�eR�km��(�����ϭ�mK[\��Y?͐qB^��ܯ�$*L<t�Ή�78�!�Y<F8��K��/�YI@��f��$��2�{>����;��<���nh���K����{��v?f���ki�"s_��<�2��x���9�EO������ն1����iH���R�#�5n? ��k���C�޽��s*��+Dk�����'��K0⥏���m]ז4���� (lFf��Pk�)*CNe�m�v*O ����3�z�<�7���j^Rk,K�-��e{���4P&�Ȼzm�tq�J���o/B�;sȆ9�k�g���9p���x�<QRx�a��]#���q��Q����iC|.�c�ųW���&�u5y��̉{LB"C�v���!��3�\�ק!��s���D)�hJ�����I�%,:J�I~���j����. ���޾}�y�Q^���WA^�-�x�ݹzoL�
OB�X�.Feg�^)6y�K��քf)��~rj��Z�Uy���V.�_��J���%�ʫi���T(
��!���C�B��6[)�R>�g7_��X��������F�<��M*��?;�ִd�)��˦��'�@�{MH��3�۶��{�ߤ>���,��T�7K_�^��u��
P6��@�Z�@v�R�ʏR��Gگݼ#�Z�PRy���ѨK�Om�* �c���lZ����W�s��{��a³�'#�6��&�<����Jr��~T����/��.���`��gT�/���}h�;�QcR�q��￴n��w�W��<f�Wj��J�����<�0ev��u����̺?4�g��)ˮ4�Q27�qZf��M�]e�����s2��v)L@�k���5����X��8 A���2�;kZ�r�
����F���c.o<���_5�뚺������fhTX�;}���r�+}��w}/�9~Vw[��zP��A!7��N�UqKh!k��׾�ȷ��&MaҔ�2FE�܆���Ŷ85�-�z�=����� �LЪ![����p���-�YO��fY�LJa���(ps�!���K7�ٴL;9�?q@�>�E���W��G��dm�����)�6���H[����d+��睂��7U�e��xV ����FoH���ۉ~�=���j!�]�:�؛/���E�_?v�'�U{����UٔZ6�ĄMF0�vSx��v��\t���_^y���th���U�>
P��l�'U&����y(Z�10*�ݏ��S�j�\��%j��m�z��Qǭ�o��n����cc4gY�uab	� ��A�ڰb�^Hb؀�傈.�c�M���CW������ȩ�7�S����=6?��z2���F;x��
��Bz��+]�ڍ���{ }"�Z�l�B);���S�4�����c͛�^A��B�"{�oC2��0��ǉg�G��q���4��R��L'V9�7\���*V �o�{R��/�~5=���z�i�#���[e�Ե��e��(���
r-z�2m�U�YEq�P�T�i�'W�{-|ֺk��5�Z�)c����r޺�j_<���j�3�BʵY#{;��Ws�μ\@n���`��x�Kq�5��汃$;m�,c=Џ�g�r��d���-K,�n����Q�F��+�ןj���^>L�;��W�n��[6��KM���	ʫnB�R���%�������҂��#���&3e��m�yx�Y*�m��s6b4y�%�4�z�\zO��et�,��7�~���;ÿ��?����ȅ����x"5��?��&A�Oo�gh�D��,q�݊r��30�M@_;�ޛ�^~�,kCp�DL��m�k��	��d����q�J�D��g�Ƙo�R�5Cwc�4��_nz	��"�^1߹�My�M�_em�J���>��+t/���CG?����>��G�6%X�E�4kcv[݄V����&�`r�Γ�
AB}#V��݁
�*p�KU��4)�ڿ�߫�s�.�VC�K�ӂ�X9b��{[S�=4�OX�#&ESh֌w�VB��R�ȚR�p*!���ߍQ��w���}���n�������y8|�a8��9�;A;���*���i6�`8��oË�lF�t�Nf ���)��<*��Q�y�yTR\��cZ7����v������3N�kc/��-��!��X'�ە��Ä$׳��P��'J�NP�FAX�[��Խ�&p[�fdI���S��mf�a���J�u���rƨw��F�:F��wM�B�R��R�ˆ��AY�/�/ ����V�š�5��~����s��(�j#�c���ɨ�l7�_�^�ųF��a�ʜ�~�O��z��$��:�F���q��t��^K��t55V��bX*��+�>U��y|O�6bX��wc��^�㔜{���cu�ܿ�e�����e�6D���X�\�+�*gL�AnkX= &!��>�1�-T�CC��`��K�?;���2�ub��*�uQ��x%�aD�h�/j����N��6�n?{k���M��Y�SP������o��_C�&O/=�S��<���;  � vk�7�%͞��nn�A�r�4w�n�ȟF�4��8��<�8������X�ʍU����w"�M��U#ZC�K�#{�{ǨY!2�����Fd��7��=��n�S_�#���;����?��z��=y��}e�ڮ0k���pvE��	@��(��5r6��<�EQH�� =B	=����Z݊��̇@6v��k�W����B���c�s���n���	�g����,WJ2��#^���4ή��M�F�.7�@aQo����5���ۄ��<m���_�:]������#�
|賳�C�)��B��nH<�T��f'����Z�BF/21����.�T��K�l^�jv���~j�k�x�M��C��i�;��7�:>���2��+�ʣ��Oמf(��Nb����$��Dq�[gw*�+�޽��t���HJ��+�c=��$��,�I�
j�����%�]�\��E2{�QT
"8�'[�YE��z��.e��d^�:�*�*���bj�� 3Ӎ���b�FU�v���2/]%Iŋ� ����K�����\�,��U�dH��hZS�}-�*G�"
��\�H׀��^�TT0����m�w�0G��j��?4fF�p{Wv݃U���y��2��L�w�^��52�'��S���q�0�:X�1�Z!�c�_�QEW��3(���W�:I�@�E�1Y='H�Fi3���ӛK�E��r�9z��4<�{��ڍV��5���!u������[!�Qyʵ��z�z�vPGi
,��S3#(��.~%|E?�ʆ�|Fj��ŨK�
q����ˮI
�4�RX]{Ԭ���>�#�;&,߹�Ǯ�$z��8ձn������C��#�c{�С��|��?Y��e�p݁�e�/����!�B2�w2^��C}sv�9f��@W����
��|��n�_���B�a~k�ƨU_.�W�TB1��w{��V���}ЈX��KH��I<<�t6t/-��xS�3' ��*X/|��D���t��Job�-�w�᎕l9���ۆ{��3�w쨭��?K���;�Ev%!_�=��B��ă��J��W�:FJ	S�Gypx��#�������O~���"%s�-Mn�y�y_�M����e��	�"$��5VB�<5�����T�^�uK�� ���j-���-3����۵�r�Q��b�1�mA���o6��'�y�(�DE�U8z�*2<�fl�Ll��"_O6�B��ʹX��C�UZYG�U�M���:j�����8�����.��¶v��._c�R"�xg�u�鞴M�s��(Z�Ѭ˵����m����{�0��g������7�A+��XU�^\ka�sKeh��51x�qk����:#���i��Wb�pv:<G$=����(�/i�J��hv�)0[��Wg��W�k�|1D|��ܐ7@5�0��t���t�#��
�����Kjʰu�ߍ���;�W�]�b).�P%,�®����V��d��Z�σN�awK�TO:)�H��}g�ȈT9W����PTk d��+�g��9���9<�dSR��35���^ܼi����ް��Ũ�y�����4��,���?��]������] k��Rmֲ"�wt��EZJ@uϢ��`x�6k�F���9z^~-?/Ɇ�
���̡G�����zL�_u�����댣�Y���{�ĭ�B�>�Q��=Gk���l^�<U�P��k�`ޣ%����������vV�1�Zл�>D9��a���({�l
P�l�KW/�l� �6C���'e.\�ݐJ������|u�N��饾m��i��D?{;%A�;#��&:rYs���В���Oȶ����]%΋ ���'|��޲hh)��j�:k�c��f��<Z�)�!��8�8���m�r��u�%�o!�4�����%�j�����4ae.Ѷ��6[I�av�UpH��F2��F+^�%��j���Y���TI�_�*�)��������fR�C�e��HE����"�5���zԥ)��e����#���IW���ݦ%�M�W��IG�U	36��>���Q����y�NI[{G��:)�yt�|������*�A��=`��P܆g���r�]�b���DO�*:׸��b�2ec�=ZC-�8�3w_�̽R�G�ɫ�W�[`Π� r�ȅt�t��G��[���J�VK�O�uj�+m�cV�X^s��
`Oe�.�A���k/@Jed�8�!��ލ�T��J�D&�y[���]�r�����U��u�[9��l�M3p���yҶ�R,q��;�C�bi�����~�.^��Qf���P�׼������]�zJ�X���t5TX����c|0�6�ɏ��G�A��"A��^������V=� .��߫�B����2WY�
��l岎�CI�b��x��ݴ
�>1��-�������{���.j��?{:�}{�K��
g��=á��Jٚ�]��#n���e8�4y�rB����	��^�
�=V�%�2�
*(~����7��|���a~� ��=�W�Ͽ���/}���{����E"Ԕㅌ�Ӗ���8��lл0-�� '7�"ׄ
�Tȱ�v�p��U��2���Ƶ���`����q�2�eIR��4�D'���
 #��z�7�'Ә�oh���oܓ�Y+Y]�	���nƳ3R�s<����[_��D�f@*#��j���dnу���L@i:��x�Q�^97F���������(k��1P����K>�E�������jF���\��Wv�}׼lE�*ZT{�Ǩ1�)�W#Zm�z�<�� �|W�V���u���YJ�Sk���5$ś�W�?�,W�=��<�1�9n�x�*� �r/u��u����]q�j|��Oh�y5�2%��Ek�����Iv|�$��ک4���u���b�����@ȑ�Izs̧�ep���-31#��! �͏���R��V�uQH~�Qr��ַ�H��-�)��{K.��@��Z�R���㱂Ar�肱�M���������m��y����Q
�����y�Ϗ�w��/����K���Z�K�W$eTi[��.����~/�h4�֟w�V�>B Ѽ�x�V�SI�.jw:Ey�׌c@?nZ6Gg٪�e�0Z3.�N�W�ݐ=��kҋn�<=��x�
�ΘWQ���a{J7d?��к�w�=>�������'A�1K��$��=�n�V��u�Nj��ފ��8,=w�MenQ�ý�����HR]��WYm -23La\L��,��%��MH$��3�����O|lx�{�	B0�m�����P�ax�/�� !�t@l3F)ڵ�j�x;z��n�2$��x\�^�� ���߳"!���(�b�Wͻ�y�m+�}g�����US��\@���:���J�֋^�V��@	xv��2�*)�Ne�3�l>����
N!hl���7^YS~/ec�q�P0�èxg��MMiQ Q���Nn&҂����^�K�YuM�窀����[�)+���j�J�;k��o�.���+S��ז{r����=�l����VYiy�Ω�[ՔݸU�������Elb��66��B�IM1����E)��a���SbxM�fK���A[""S1^�Hw�a���7��0��(�Ҁ�h[�iL���#v���W��rx*'�@X\{תUMO�g�ZQ��X5�W��
JZ�ܴ��ٷnc�D�N@ش� 7M��ē��֔EmϘr}jb���)��=Z�g��ޫ���j���Kn�@����r�	����p�X���8�k�ڿˡ����ۯ{��G~��o���'��ϔU�� G7q�Ȳ�w�':����S��,����Pt��.��<��9�JW��ʼJ}v�Z��ݒ�����楤�(���m�\rX�>��CV���<q���(��u�Lϧ�6*1IHS�\�~�1YO�x�^�����7}��|Fp�ŋ�$U�	~9�+�Q���:&��B2U/x#a�l@@
)_� ��鱨#VKj�j��-�tFJ	8o���M��]���E������	�y�y��O~�Ӕ�m^}�ᩧ�f0��&0�rO��q��-���T膱+�Hge��7���q*T�9�x�h4���_R0�KB������s��R�׬�@�[�,�v9�z�Ƭ�o��wc�tLq�e�nb4�jVeC֓�!<v�7�w֫�+���c��ެ��I�t\n�n֓��+��<���n|�=�=��yo��e77i�+�3^S�����GԸ:FO
]B����W�\�cm/f���n��%#
��A����B��Q4|R V�s��)���U�P�0��
bI��j�M�����0Ÿ��@�9
�F?R[�����9*2_�������%Rs2�z�o�O�u2
<`���Z�;E�8�m�\��kF�
8+��ll�o�p����G�40*�P��Nm�y:kc�h��e�)�kQ���k��9�~t$A�Ǽ�fER�g./��������ܦf�u���n�%~�?�(��Ɠ���o��O~����εw�
�mM��O�K!���n���&\v����=,>������r���ѫyLSAjn�z7�S�h� y��D�aK0G�E���jy�,��N��j�7=��5�^w��%�J!�ICZ��$�p���s͎9}�\@*ָ��>O�tۢj�Oר��f<�^�8U��e�w�<��)�cJ����ޞ�VaƉ����Q��W�x��p��iBㄉ)?9:i8��+
�+��u0�{�9�Co��Y 
�e�����KW��g�l��:k�>Fu`���=�ha�H���$ż�B�:�fg�����&-��Y0b��3>�ɉ�]θ�<�z�`��I�2��LI$j�D0����;�@�}>��5g��)8}����S�8������K ���L�b�U� �8�\]Wr�^7�3*�������`��)k]�6��O�p�S�Ѱ��2�F#i�8v�b�����V�W�T��徎����;�jc��*��h�����^���ⶣ�y�l�^��,O��*%F�>3��ܯ�o�3ctdl�0�deT�'��r�P��!�=�$+C�s���|?i(17��ƍi���:p"L	K�U]m��Ϥ[7�X�ф�yp �)j[>n���^l�`�#�m���^�p���]7&�]�ʯ@K���*�3�\��9͚�TH����&�Z��I�*��xk���7���ٗe�u�wj�5O=w��#A� 	��Hɑ,ڎ�ر�(�Z�W����%oN^����!��Ȗ5��(J�8�	�����y�y���|>{�SU���$f�]`��{������w��8�~�?S�a��7Pָ�MGLL�v�'{�;8Ws���_8�.��.=v��O<��^�I�r�iC+Nc������gs��{UH]�In�X>��Ra�`���eБq�ߏ*���ռ���11�AxP��ī��JoR��5D�H���n��Nh	���	�<�!�:UH��t��aN5	AG�t?1N,��_uPlf����֙�����|t= ��M{��(��o}zz�����(t����x�ާ9�������`�" ���qOӄ�O��b��&d5r���	�,	oI�e�5��͓�C!7������dx�E�t��s�}9:�eD��
��e-]�2��z-r���t �a�<K�B=���~T&��ғ��zD�v�pI��=nz9b ���ǈ'�/#&�Z�'l�����
�\y��K!��3R���Cm�;�>��6I�Mf�x��Di�h��8K������ @�%!�#�.�>P�]N��^��=�w�2���	�vjl׹��$����iNg|w���~"SIATi���9�N����?YϞ�^�=�)o��3M����|�^ON���&n������om�9�y�J\E)��h�x9������{��l�׾�$�ͣI�/���
��Ԅ���=�1B��h�#fp�!�f<��D���(��c�mD<2�������*�#	{D����� EZ��=D'H�"*�L)h\YZ��Kܞcq�b�rL�mD����8ׂ	YȵiL����ަ5����w�R9�FI� hRcZʎN{ �ďr�I!�ւ���=w|��B*t�������w��ݿK�����z��<�N�hݛ�R�_g�wT�S]G�7�^���oGO�E:^���*��b��ӷ̹��[�Cc:A�G���BID�7`��M��m����� -�0P2^vH�SQ��^��K-��c�x^
B�#߾�n�GMٽ�����[�6[�k��ff�bn����m�0�ܻ)n}�fl�a�B����/ޖ�o~�s.��i��4߼�$�5<�ȹ������g�����m����7���w�ſi�,Fx�����[X^��:}�/##�51�NR�*���R&?�gM��5������_��*�4>�/��W1,|�Q��Q+N|m<��*<��Fl���]�G�ߵ8��C/x~&L�قYld�#�����̅�"Sچ�����4��^��|vP%�k4K��z�B���I�"��������w��tC�f��b�>�X�_�܈�5�=��)��}��#L����k�e��+a�1��s�~�s�]ĵEt ���;�	����{��Q�g�|6Q���y��O@�%,���\v����D���W|�Y\�on��sf��YE�A�摪�#��ܼw�=�1Ҵ%�-k#E�ͣ�H��d���M����!���:rī%`��`��p���O|�FK��
=B	���@�}@ӢlqluG�~z��s��*W�Ja�V �o��i�\�F,�tn���F�%r����ҍ���m�p����p��zpW�D�
��4k�p��l�\;���R����_�̧?��_|���k͘j
F�q+�:�"�ruq�� �E��S~?���Xy�.����R��Qk�;g'�қ,)��@P�����p����E�r��k9����w�d���8Ɣ�P�{X��O|2����nld%sv��h0i#	B� ?���;�34�ѪwF�!x�D�s�3��ͽU����ݏb��m!�ז�>=�wwP�F�<c4Pio#�`�����������e��fh�SF^�F��������y�=J�h�y���S�>�<���{��a�S6G=��[K�����f��x�/�I�Hң34m+�"������3:�Jo��P8P1:҆QYg��e|�Y�����mg;�"I���m�S�a0{kgiZ����2�c=�.�N}�R�ʳr̤�0E��������A3�ۆ�U��"�h��$�\��k�	��Ur��Y�$4������iC���Q{�3&�ah�y0,�*m�w��\�^z-�P�i�vFa�{��J���!�H[D�?�;���z?�9k�� ��<K��|�:c����6��:�9�Uʫ<��ʇ��MQ����Ƕ��Pj�?��盿���As���w~�f���!��|�f���g�ɕ���7����4	.D����U�q�{�E�u���>װ�g��OC����͘q*��j�l,�I�ݧG{C鵻�$�EU{~8�����q�<�����"�(�Ѿ�9.�=ƿ������T�t��r�������C����6�Cw�9ʚ0�GF���L�c����Q�������޹�Η)�z6-eQZ� �X(��ܝ�3��b�M�  :O�g����zj���G�~4��{�ߏ��'?6*�I��3o������Z/�56�^[��Q!9X#�z���� �������z�,r4j �������ߧ޲�<��#��_jVP��^~�ы���w�!Źs����6|�@��K|�M�'���b�k}����-��Q��?�'�L�4���Av������wx�4A*��ƕ���7�n�^�_��fk��/|�����o7�;�,o��L���~���?�v<[7�ʧ�e��yq�z*�܍��}��ƂҊjy��9�p���X��7��w)nOj\i�v�IU;�$���G�l�
+j�go���ni��K�>�]�a�D>X>�$�/\OˈI*9�~��n�$3�u�S��D5�H<�	�����>
ì�Y~��i׻ޤü�óm��#�z���o1��Wǌ�k�N���E�'1-�B�p�Qw$Y�%��}ֱY���f3݊W^G����|w�+hSU�W�!��f�6��ڴ�!�k	c��"#}���C9��V�ȝ�Q�L��n�|oǶ�e�V�s��G�n�.R-2��GJ*�0i܊Ib��8��탧�@�L��*cֹg�!¬�Ñx�c��b�H�tI�4ܝ��\1��p14㕩^��Zq�� �M�E:#y)��E7�s�^�����ǲ����]�/GbfDF*��d$G������B��|�"�N��k������7�L�\~�М�����<��u�5Q
�`�����j��͛W�����������,��\��W���*�����b�g_K�4�8��1:��z�H1.�nPDw�N�t�Bl��u�������M�ކ/����γ���S��Q"��Vtk�dC�ױ}Ӓ>,�jC�Zˎ���6�G}N����n)���ԙ�a+�G.>�<F}�Y���k�gt��SgC@=X�n��v��H֭��lDH/�1!�z�a��/\8�����͝[6��4�y��aA>>JN������w�S_v5���B��޿����1emO7���'�'��c�P�2B�
+��a�C�J�P0o#W� ����9�
�}��-��!L���x.
#�:�|�B3��:'~e�6Nw�0�{�s�#qy��x�o�8�����1#<1U��P���u����q��p^c�-���vJ�I�==,יU �B�㤰F>S~0jԡ����#��W$!��Tg�Do����фH�ۥϞ���7�RD��i<��u!`�U�������du[B7�z���;�u{;r��B�������E��Ѽy�=L�������q�vv˞���x���"?g�(�ߧ�g"��xQ�WK���g۬�m,��ք^���n�V]Z_l���+�{�7�i�Y���"�z����Vי�
rr�`�
�XnYFe4"$���yn$ͽ��*�`���q���xSWØ{�^	m	�4�����n��`��H%���(�רlG�O&"��Qޚ�6��=}Z���%Ⱥ�H/D�Q���#a$�����5<Ԝ\ȱ�+�c�H��I'�8����с^o���J�\�����ԩ[���g��G����>�~��]غ�LB@�J��=�\}��&鄥Ū,�)�±��b�U�'�CO��ֈ���?�u���+G��]K����#%�?#X(�<#�IC}w�kO�5�2�^KE豣�*����襴�?�GX�=��[���%�p>sU*�ȡ�8y�Ts�q�
�S�<�,�>ǆ�5F����杫7���o�e��ɨg6��W7ќ<s�cΠ�7�w߹�b_aR�B�����:�uȆG��$��������.9�7�4��/7����?�̟:ռ}��8���y֎��
;1�, �h\k�M��4� �О�����'k��4��)L��,+�^�k(t��my;J=��(��V�����l*�\j��x��3���ꈃ�u�����K/k���!	I-�:(��7���i����0�l�bL�G#��X��kǝ�P�~�5l2,�sJ#4�D&�(��ni
.K�_7l:��}�����l\��慳�B�b�HI�V�����_�ͱ��[�/�.�q7׼��G��`m�oɆC^��k�kP˥M�gɱ3�`�adb�Z&{�J�������o�ܻC_vHj�]��
ē7JC�gs�~c����z3C�e�����(�h�yWW�ھyg����f����� L(�rd�^��lf���}��"<����>�� =�>	��6%�q%C>d�F�'øK�Q�j�x���0�N�e������B�{�T����Jz��T���%�HDo�g��C�9N	��T��|�4��[4�Ʊ��Z������x�S���G�x
B9�G
�&G�y�Ԃ��w�1��/؟�	��ӵ�׺�kחZq�%z���ɯ���Ʌ�}����s���x~�ŭ7� �����*i��¢C�
E�Ǉ��\b~���BG�4B���������V�l�}XcnyH�F;�P!�h����rRkz�ȟ�?�k��g�u�_�淛7��l��2���̏����^�����Rs�)n��a��_~�����C(���:P���ϝk��o�6-gO7������?�I��dS{� ��{-<�1�(�Uo�� X�#4y�� B-V�THj2��>��%�>�T�)��d<�x̆+�#ސJc�TũS'�ڲ�W;����r���9C�wQO�^|�;C�[?�)�%_j�@�lݿ�A�x9��}u7"��]�B�1v�#��g�G�x�<G�s ���  v��s'¨[�q#�6�"�>��J4R	��P�vޱ���;6�!���-�3�����9�8�֜��~��Ј�[hD9b�m��kg�DH��Bm��S.]W�a~\�=�����`�5I�������ޛ?{����:d�:�ha� T:�z@Z�އ 	F!�LS��co8�O`��i�Djc7Z�F8-�/U`|.T#���s�w�hʴ��ua�Cb���о�=�H��k�p&�so�h�`��V�����b�raa��S��{�0z�ʹ��0N:^�21�g�fHB�xA)sM��]��ht��6�Q�^�������}�1�K�:�B��1(�u�J�a"�`���pB��.^y�����"�{��_�6�?��k�~�������]�l���>3��!�T��3�jC��wܒ�R<�B<��2����w��5<z+����l޽����vm.P��EڒI����G/<��>ͰZ�b�}v{c ��� �dhSoh��h����~��<8�Q��>�C�PzI��l�"'ڇ��&�8���8��Ge��<x@o������揿�fMB�^o`��)���j�Y�q/f�!�c��U������	šQ�-���O����5�2B�Cd&��d���5jӱ�	��mHv#��� w�ݯ�"7ji�ރ�D�f�;s���KHC)]�C��]O(T�Y�U�&�T��4���83�5(Reg����&N�a)U��a�!r\Sg��|W+�r�&q(�P��j�[$�E
�(�� �m�%�S>�K�K��YcLPo������f�u'�}vx>�[�N��ʅ}�-<�;����5
x�sv|�h\����B�����(0���@C KO��:�{Z���B��O�e�G�]���:��U���t$Q*J4S*?�Cq�U�;��hg�$��OC�&���Wa�߈5�VF�Qe���u��#�;�Ht��}Q���a�o�N��:��G�&Fnlȣ1���my���*� ^{�`��j�^��9�{G%�1u���s�F�H�3�uGe��&�7׉�i � 7��	+����^:�O�� ��'�ӈA8)V"P���:���S��P�g)������qF�P1z8�B��gѓ�)�B:#X���q��,t��/���	�_��^�r�%��]���2��x�D.=@Wwn�g�nT��RmI'0:X0��U�#.�x-?ߪ����ɼ���uJ�!uX���IH䷺\q�)z�FO��5_����^�\�jdW+-��|���l��?j�ܹ�ܼAv����L���<����m`1����M��k��\�4dv�]r�!��O�FA��n�o����|������uE%��A4 sz����;�|x�\�n3G�vgt���;ͭ{�x�vY�>ˣ�޻�^m���ퟆ���(�K�����;��_��P���9�����g���g����}ʯ�7�^G��	G�����2[+�՛��k/2���^�b�(�g���@�4�O���)��}��(� ��屍 d�?O�^G�)rMź���tJ,�8nx��HA��L��F2U�"	U>���m�=�����u����l�t@�7�t�{�����G�g?�k��T���aj�gK���	q��:���ll�JD+r��_�(���d7���gG�Ď�����dx��|��c�I~��6��� ���f�y��m�7�0IY|>���L��U�*i���H;6}'[܃]��h���p�I9aX����2*��D/u�ϝ�5�o���9���1��������s	4�~���W�������Ҡ�%63��|Ny�F*L1J2�y�vfA�T�4�k��2)�2��4]w��Ix2�E0��
V���K��*���&�D��{��{<�0���uי���b���N��i[5L�f�>�T�L`0j ������¹��'�z�&R�1�2�p�=;�L_��c%ω�C���Ɍ�#���,��m���˱P�M=x��7��k��������y
@i4ei�󈨻�)�?�uif�]*��Rb�l����pQx@��b�J+[+��t�o:噬���$�a�'f��^&(����{��6?iX]�#kWCXi���l ����L`�z*_ϣr��娤�̑�ם����A��y����8�ę(g��
Jr��,k�C�������^�.������懯�I�o�}� s�J��L��g�p͌��XgN7���f�HǹՕ��������!B��v��=[kd��\�cey�y��+�_���n�CڻuoeI�����C��B|�f��1��1�>��Q�-�7��<�(����͋W����9r�Y~�W���s�$��m*+{�'	�7e�ut�J�,�:H�2�e�s-�S��NC�F$z?]4I��)T�ڏ�e����1:֫1��"τG�jTH�:s��fm����KЮ��LH��e���V�?���^��#z�����5w�>��k���������0i��w~��f��^ZZ�}e�ڻ�ܠaJ��w���j�S?��#AB��ԑ%f�*M�s�qϸ�:R��]��5��g��?{��5����f���WY���	l~�8��'��x�\L{��p�z�5B�o�%N��_�00�������D�a���p�^�לY1�֘JْJ;����gg�rQ�΄)�|p���������Kqh�z_��4�n��e�ӧ�6��?����=������i8�ϟ�K���v�OK���x�x�^Í�Q�K\[�jr��I�����M��ɺ_�T��{8)D
&g��i�T3C���g�O�;s�Tsc�k�����	h�2��n��2��([;v_�B��T._���/��7>����<xx6C�.��=�p�1�<��Oi�f�N.�͎�SX��:e�לy��m�;B�~�ͭu��2��q��F�cR��P��zZ�Z�6����^�~�T�%S\�z:vO2g�ʜ��dBieu-z�v��h�pax
US)��?w�酱�5��y��K<ћҫX��jum��x�=���Rs�@(����F��!��qz��d��$��� [83�d3M�{����I�+�<N�׏��>z3ؿ�Ԑڅ.zr���̟C��Pbޥǟhnߺ�ܿw�&�o��+��Լ��_n����Z�n���%/��ֱ���E�Y�te|�ĮP��1��i=̃��2�>�f댍�I]�#�RqxHԷ/���A@����ٍR�w�y��6Q��a���(]#��w�}�XV�|�\����d�HG*�n�)���i	��>3��9P��	p(����jDo��9��<�B��
��e�U��Jɘl�0�r����r���Ϝ{Kv4�3��<q�D*#PAZ��W�i	��R�<�%�,E�{�V���~q��ѣnB��;���;�M�"okԣ�/ǈ0|��7ud����Wx�m�,��R)g(7Yb��ez�ɺv���+��c�l��KD�%ԙ>ED&�[C�w��r:��yD:�VUY!G8a�a��Q�x���ᣑ:��VXx��v�k<Rg�y�1.���d���>�>���+ݐ�U"\�H��&Mj\�aH�~���z���ݨ�Q�q�;��p��L�<��M̳/�U ����BD�B�[��
��������K#�M� �/s��9"Xܛ2��F�~�Ȯ�P.R\���S����C�7����� ��[�Bu=��\�����<���Sa�u��a�4mشP;�̕���m^8_3\G�Q0F��uu:F�cG�;�}j 
l�˭G����~�f�����)�]�6���V��I��b�Jx�9ElOp�\�3O?��C����u��z����*ђ��@�4'��W�D-�<�;`P�*����+���[�����?|=�h��]{�5S!$�Cs=lę�y�n'���#�t��50�18��ﾌR��&]������`���A����Y�;��
V��o��5�׿�����|���@����y���w߿׼sa2D�{��5����(�9���fԟlk6�<+�(r�>���!O���G��4�j���k1��0r|j���Ț^hz�9���O�A���b����8^�]��٪�<���p�^�2]�T
��7z�%"��hg4 	R�%� 	-��Q��Z�t�g�Q0���}�{��#ͅ˟h�=�l���?͜���'Ϲ�46�5Ԇ�e�o�[�pm���� �E�kX�~��ݸ�u��p7�\Lb�84���C^3Jś_Y������@�ͧ�����z ��2Jѱ�;%Fl4pɰ��%���a`���G�Bt-����:�Z���.�֥	BF$cr]>փ�����fWF�,i�Gh\��>��@�U�ǕJ*�x�i�E�O���;ʓ�Bf�|��}�s}v�z��4Gߦ��|�aı��дL��9����tc�� 7�v�<,�nu��<FZGtd,������h`-p�K��V	��qQ�%)�S]���e��F��0����ĵ�^��V�3$�R:E��)I�C��SA<��d���~C6�>L�}�e�ܧ|l<to��ŋ��~��~��_�Z<�8�lx6�;��Ps�-��"��B$�L��.��,H���>��[!����IO�:!�5$r�V
.[wZ�)�� ��W~�|�s��1=^3Y�d����M�Q�x����{X����_~�2F����;������fS�v�^�ܴ��fJˉT*���*pC��~��#��ؼ�d�oSC��z�ܬN\�%to���ר5�<nn�c�Ż��^Bl4'榸�G��r���*�lj� K�����=��3͕w�mΝ=�s�^����{�o��5�8H�e.?J�ރ�F�ʞC��%����+b����WX�5����_d^�B�7y�C	�$��ģO0��"���Tx�
l�y���De���yd���l�3����g���n���L�c
�%BZ��7u�A%q�4Ó�2��������mv���-y*�+:�+:�2\�M��z�������Dֿ��Ƹ&0P�R�{�TP�<����xt�
�4@�gT!��S�������R��׽�Cś*��a�λ�4���ꗰ|p��s�M�!��?e��+ �x,���WǛ	���Vct�t�h�t��e����}�?Ԗ���i~���"��r.2]l�ċ�l�2�3ܧ�Cy�z(�}�ʠ�@n#��������2U�Ai@���5B	e����G7�Svz�"i9;E��v`�X>i�M#F��&?}�1�V��ȁ��.\� �'$@��oY�*�SPF-��*�`�aǽ<|�u�����PNd����Y��싈���x�� ۩nxx࿟�{��t�:�m��q�'����WSo��7=�����d\�*�С��J6��V���v�ux	*��g��usG����J�dj����z1Q��.�6�/�oWu�BE���[��zv8�#BV��	)�}S(�	6�ֿ�H�q� a��^��g�m~�!�0�/.�n�U��LY"�72���dS�QdG0-e�7���3��M���V��«�ԃKg�s�ᙛ�X���U(]-x=G����Z��f��Vs���4׮��\��Ǧ"�֯�V<Ke6׷��$��=�pq%�1�}�3��O?Ƈe-'����[5���]�C����pvi�s5�N|,�'�m��6L9�2�����N�����X<i��?	>=��L���qbclj�9wz~��X��g=V���;B�5�^�8u��J�{�;����''�)��D=p�lF�3֖�\r��M8��7n���й旞{��9��߰r�.`D3Z/�[k��[���u�K�X���K��εJ4��?�l?�.%�Z72�Fv{�v������a^����&�f�8��!�{��y�q��zޡ{!�vI����;e�ʾ��7�Pm�U^~�[7��=sv[Ø�F<1�s�˸\�q��MິL�j�K��(Jk ��1�$�QV9e��DK0z���{�ܠ���<I7�F�v��Up:��c��9��JA�t��_{���0m��tEK��g�g�<��3���&����SZ�a�M�0"�٣unF`���1~�������Cw޹F����}Hwɓ�bX���  �I�1 v�$�=�G�!J}-��8ǡ5�>����X)tD��/����޹����=>;�q,�֒K?pi�����R�.sS�rm=����Q���!�k919���:F�	��Ó�i��9rz�i)j��nQ! �[
��)7!���G7��v��<TԽ���;F/�GR�,�M�a?�$��J���tu{��w����:����}ɦ"��� ��\���"tsS�}��5��&�-1eM�������r�+^�fQF���ԓ�4/>����1�2���W_��N^>�O�[O��l�;�V����|��Q�x��K�����ʗ_ʦ74�09��z���W�`hc�)]>2��6B/�A��yB pQ��B��SA�:D?�2�%� ���)��I����`=L�6�?~�R��(��òw`�^^�
��O�z��G��g�'5���x7mM���T�l�ȋ��_��F�����x��k�B������O=E��ts��"��&7	%�`RC{�-��]��0V��(u�9���1��v��*�Nٶ��S�b۫��?��[�|8�ۧ���(��?gX��y�qE*��g�7��"�B�]��gv��$��?4<~��ɳ��bDmӼrx*��T��5��=n��T2�Y�7pa�u`~~��Xo*F+7\�A���ޛ�$���`�1�'�6kr)B~�b�=)���12�b������H�$J��1>9D��0������$G���z\���i�|�:\�&[=�,䤄R۷���u�~�a�G(��u#��ǝ����`��q㔌ҋ�	k6��=��Ĝc�u�:^��իW��~���X�_�9�y܆)%Z��	fy*��n[/$���e쯻��⏥�v��nY!"�Y�VTt:>Cr*�l�ϼp�k���gb�e�z�a�g�~��C�|��]�ܧK�|,�Y�鲟͓����UX����-���S |�l��~ȆԚ=�dB��6�2��R׋��V(�$
z͹�N��{W k��;W��5���G����wjDq-*!�q�(|�<���&����Õfx�Q�\�]��3ǟ���bJ�|yy����#?��o�Ҽ~��T�j��_iN/�i�]��b��UrJ�lQú�@5W�Ad6ro<?���l���<d�g�>�H\3
�V@)��w:%r�H�P�fs��у�p�')���eY]�յ�ם^ZF�|�3fb"�zy=��������R������!��^����w����/�����K`u�����J_>��
��O]���//�u��ur��r��YD�O��`���&�>��,�>�A��x�u�@(i��ID=���Ͽyd�S��;�����ȏ>���M(Ep���"�5w���5��!.�h��k�����ll�ޱ��s�-��Jn��GK���ƥX�pA�8at�e�.�=r�`;Ȅ���r9�{��T��d(���!�q�^v�-��<q�L3-�ޒ� ����!Ah;��C�є��K��e�|�K�n���u���r��ȑ�,/Dއ�U��<�I���{"���0�|��gX�}~_#�O�܍��"�v��^%�؃O�\��#5�5;���8�7u���W��/�����g6��';�\&q�&n���G!OR��`�=�r�a�Oi�ƶK���T��26Y����w��<�DZ�q���fX��
�ŮG�z&q]�����s�����i�q�����瞍\���uk��{�)N��ajx��o[�v���t	��>����GH7�Ru�VO6s���P ĿTT�d%�HV��`����L�a�u�@�����/��4�hhX�Iәw�C��z��m����(���?l6Q��u�p��vg��à%g��t�ù�����fh�^�D��;w���u�I28�Լ��¹-��")�1lM�����|L�B��Y2h�,C�v����;����ľ�A$rB�`>!N��<������4�7�8Ƣ���ǰ�9n�F���$I�kc�)��Mmvv��=u�9�~�d�"�L�����2Z��>C�^*B�>��\ �#���|�`D�Z'��_a��T�"�z���kD:iU:3����OC B�]��#��`�yu��܅�;�h�������M~��G�]���l��������z�t�uQ8��ѿu��)�X&�%��իH��,��n� �����|(Cd�GJ�Tp �_tW�?��w�fɛQ�7����������$��p�����8��zO ���'��GY�VHl�������4���}+64��c"���Q(�_͡��]p	>͚S�dv A9?�|{�K@�;5r*�Y�����G�6鸧w�	���.5��§��g.`���,S\c���&��0�#�M�1ׁ�J��1#'m���?�������[o���7���������G_�vwz�~��vdX�Ji7R�M�OJ���(�|w*��ׅ���R�'9UEg������nkSUzZ��o���N��>m�Q7��,����G?mN�3�܋�b����h��v��Azb�tĩ ����c7�?A�°w��1Bɩ��v�2���|t���q���k�L�<u:Y�[���#�^��<��q�Q=K7�����|^k���^�*��k[�ܳ!���y6�F�����벱���G8|}e�z7l�E~��[;\����c��$�-�J^�Q�`G���x�He�]�8�)��#�w����\���JE�W7����!�%�s��Ǔ��j�4���d��g������o�x���O~�q�@�EHv��=��pNC�>'��(,���n��m����\�Ao���7���g�ˏ_�S���o."�ei���9~r�m�!�G~��m�v|�*�a�ƙۻL����M0M���Ge]�r�Ր�Ǿn�����so�������+���h�'��{0�v��%F�/��G�w��Q������G޽�{=<�xV��������N4��$�m�0�YEA��0�c�˨Lx��%.<y�Z���4J1A�������tOtf�c�8~o�tK]�T�7Fk�W��M�������.uhl���`s��4jb*�r�ՙ�8OCsxġ497b��Z1�4�nkVz7�u�c��vpxtbj�ejl�-�d��ټN���g�w6����4����^��j������0��b�l��Ϭ�_�_����Cy����k��O�x�3����c�A��r�k(�옵C�h�j:7Y(:7d�@���h��ôb�l�����6�B��:1&�K��[�Ӑ��KS���(��gRK]'{]�<��6�֛��A7�w�4�.]���s�Vay��nR?��՛��Ս����ۥZ  HUIDAT�]KچCs E��ƹm$C���6�a�g��i�)���'QGJ�v���åuڪ���;����v�G�a�b0�������^]�)�3j�ǨR%X2���[G:Ӝ=�u�����8�@#�.u}��J�c8�k�)o�(s�Y�gas�*	���n
�s���G��e�*N�N�Q����K�)�i*��	@��eʆ�	�0~����`��S��������,�O��g���\|�R�s�!sb�1^a����
&��5�W\��g8��zΊ�x=S��kع�F�N�7kͳ7=��f�Ju�F2��=h���5�L�"���Ŭ�e�w�4s��{܊���`��rnR�/j�s�v2��*ǣB3��ҋ�m(,l*��R���7�$�U�g���{}��������	G�L�w{��Н�{��U����z�aZFz'Y�9�������vWf*/'��?FYbx�F�|W�F�"�qzvz�Ү{��d����F��N�M��E�����he�;91��n�H�͕OQ�Q��k� ����=��<�ϣg���5�ǭ��'k̓+D�Q���������%/��t�SO?�l�
��I���^�~��$�v�}�`r���w��${f��2gf���~����B�+��o���W~�W��������(�q��a\E
D?&��G������q#�s��ݒubr��0d�anM��XLU�Z_��[OU��e%t
9��ءl���"��µ�a�|���Wv����{��w�����c4�җ�D���[��х.�Ʈ;��H��IbO�X�2Iݘ�a8�G�R��Y���2�C�/>�x��~�y���j��g��^�&�,�y���u���lR'J� %�XC��1��k�������v�2�l��2�9��BIwc�Y��w��H�FmXh���c�q6a��:vi�3���/��1I���Q���|tTNvW�Y:ųرL(�xX�U>�K�)Y��+N��v��`R�����8?�vn�k�k�u�`��>����Qϫ�Z���{���U�P�a9�Ŧ�Vb�_Fc�ퟎ1��������Jz�b��t��:�W��lךs�(7%2��8,a����T�rLI���ڟ5�}S6��s����-¤��#Y�1"n�1b	v��4��mj���q|��c����o�1�����|6y��{Z�m�����������ͣ�L�V�`aF����n�%�BN��B�9��� ��8=���ud��q6�r��>.q��=��x�s��S��)��ӡ{��2��J�,Isg���)����V~��"�#;�g�-y:���%7'K	^7��mSNe�ۻ���Pf��ȥ+��,-^M��5�,=�ه��P����q��%���dD�8n�N�7o�n>�y����2�떽i�sO\���n��I��5�FPE	ɱ�:�
�'u�ɧ�����o�ӥ����/���כ����6t!��UٹI�D���Ʌ��f��Hc��ް��4&!p�N���.��b��<q��Y���e��d����܃R.�PZ�jT���%C�2�������9m����4�Ce�h?�*����ߣ����L���"��%l�0J��B ���G�"7o�Bq,E�n{�u��)��d��4��ܿ���� �G�J2��KO�Y>�\�v�9�7��M�g�w��3of_k矽�w���X!Ң��� ��p��L#xْf��ϜXEvor���k�lO쟊����)>$����>�`�}l����¢]G���Q�J_3�s ���!?ϧ(1Ϟchu�ڔ���Tv�`�~�l�=�V#�����U� c�ǀ�qs������~2	�zi��-+��w��j��=*$"�ӯ�����Mw ���K�A\D8��C�� �~��t��ˡ��k�\�:]��Xt#���ꆸ���t#�_��:ls;F1) x�ܷ}�!�]�+>�9�_�|8:�U��NH5�s��r�=����:��l�%�ށsX(y�~.���EW%�$hp�H㮍C��{pww����� �!H���ڸ$�;�7�������թ�=���s�V�����Y����E]׎�@b�׊�]���xog5J���ߔ.��!��x��������<=�&�Ȕ���˅�u�MҘt�I���Į��_���n���n�\��)~�p�~:��2o_��w��s�<��"a�iv<E��kO*:^NoE�w��⾸g�F�`ҭ�
����U�a;I9aճ�G Kl�}M�S�5��ou�g�= �I4b�e�Mv��%���#�<�ȭ�
Q㺞}hQ�ԩT�0��f�Zn�x=��5�T��� v}ZǍ=~a'�<;�F �ɂ��7���� �*�`���Roj�NJW�Iz�W�x+�V:t�S��Nlj����⪝ ͚�m���ڙ��B�hL�.�儊PK܋���G�9{v~4�&{�3�ݸ4�:W��*�+�o��8ӋR����q6{�L��J���)Ͷ1B6��!���I��e[u�g�v�p	�J0�`��0E�JF�B梠��n�O�ȷ�o��"q����*�H����m�/*]֔����8$�u�j�=-��Ƈ��w��`���ˏ��q]b��I}yΩK�pJ[���<�/�$��_��E$;�aKN�-aKN��&��Drrrh�=�P���Nĺ�U$O�G+��Poq(PCŭ����Ϥ\6)#>n�K�0��1b%e/BW��U�4B�#��k"��e���+�.^�E���T����ާة?�6MZ�������㢶�I��3�m��'�;=N_���8?+����%���t�jcK���A�-��
IDC�]K��(7b�?�����~-��M�r8Hز�E�?�^O�ǹ�H��:w���y��S�Kн�5w_��W��H<E�g�=�x|����S����t�v[��şQ*/_K��D��(�~~�u0�����u�
�LFȰ"i��l��p����k�p��<�Eq"��;4�
nI�=,�(�qm��|$�L��!㽒� ��E���=��~t 9C*F�{�nOcCs%��L��\��|��h��2�(��J��g�J��mE��ց��h@g��;b�Jy <����-W���6�y5��A_殾�/�'-/n��������/��?-�a>,��H��X�����Z�5�	��c�w�fhkw�R_O��2�6�$���mʲ)�]�>���6�����]'���\����/�D=����Q�LD�&�����8��mG9މ{ަ�/��B~���|�f�
���uSc��w�k�@�q�N���&����e����Э��(�����71C<�� ������o����Asu����s�ߐ�-C�[�c�LG3R޶(��y�����H�~C=E|�}.q�w'v���6�n�-5a�QS�m�����������ƀ�K�GLB�<�˔��"�zף���w�����E��w��c�D/�Aa
����~9��6��?9K�G&�$�H��2I,��4��ծ%�c��{�R"�g�� �5�lfy�V)��59�Y9�w��A��1��1s���Y4Bu����F�\�-��FBt@��bz�֦�p����aZqy� �?�\�R�ꯌvwٶr*Lv�s��Ǌ(�ħ�4=W�8�j���K�$B�flٖ)t����0�*���L!5��W�w.� �i���V�X΀�{�\&%!�},�K�}���MX�B�駅R������>��.��K�Uw/�x���f������7�d���ͤ���l���ø�p��:ŔX��@���/�d��������;<�i�}���:m,��~a�.�H�����ox�������woA�����<�1ғ��Vγ=���>�L\�x!^�Ͷ�<�4�e-�2(│�����?v�a;+����Xt����Jç	]�H�l�&��q�͛����@Z����[;X��KS���������Y��@�D�'���!v�M������#7H�������<��\�����{�J|�������6L͡�������-���E�KjC�g�A��V0E�oc�ݍS��>�Dx��{� =*l���kd1���A����D�>�u�+>�͗�ud?��=�[$��d`�4�U��Cy|�%���$?��Rr�8uXDޣ����k�"O�a�"��`d{|UX��4�����T)��vCO��{�Qf�Z\t�WJ���q�*I|�򟍸h	���_�~�����%\����})�Ϟ(�bqsB^���	����J��s�R����M3����ޕ�׋r�����V�L��zʄ��Ϧ�ĸ_��"a��<��o@�v��ߵgu;�L2k�c��n^>�(����S���N�"�}6�?�������f�ݚ�?��H�PSf՗�k���Z�W_(���W���>�i$�M/dA=�����	;���O784�H0��t���8�"q���#�Z�ʐ�1�F�E�^�R��)�����:�Nh1����ۚ��}&�֚
��0��ڋ��R\E��ܞ�h��y;/yZ��X�N��L蜤=����.�8�FJe��d~�}��&H����7ZGϏ��/��uX������v�&f���Qwn)�^0��w������	5�5�4ٱ������vV����^M��1rظ!gQ2ć�A��h�d��'��d��r@��W�����V7�i��c�(�,������橷��j�x�<�a��_t�E	���>�&�82���ܚ��R.+̳��8Vɾ��?IH�^_X���Ą��]��;��V�%4�4'��٥�S����d���
��I	Y���(2t�� �Y���A:sp8[��?N�zs2��/�E?l�Q��srS���?@JϢH���S���pC�U�36�e�����I��%��+j�XJ>�)C�5!Y����}SQ��nA��s��T��L=��`�3����1^��A��)���-}��"Y
����b����Z�nz�+k�DB:#v	ݓ����r)��P�����0��.Hc�Yu���S>4�W��5�$$�;i�J�Y���ß�&1'��B�Z6M��T��?Q�Z	��yE��0Mk��4l��=�V�ߎZ�з�cu�-�3�HbC3����ihB���d&���	�(��w�g����,�?�O> �v�E1(�#q������R��J�?!-X�Ǻ�o �l7߶U��=�H��]�ϛީ���2yP3@p����:z���Yч"�@̬Pz����|I9P��bvFԢL���c�H]�)M�Uq���_��y`��.�i�#]^X�[�*��V��eh�BEn��[!���SY5~�j\	�v���.l�,Mk��>_F�ګ��8�<���8� R<e���bC5@�t��ň����|xa�CdS'��-��5���q�Z�x�=��u�w�#F#�w�fp��ߢ0��i�z���f��]Z~�s{p�e��pou����F"8��CT[�5�����'=��WJ�9�*��h�l�~��BD��G/����-ŝ��D��=jX_iD)��;SW�bt%��2�l�.�_�"S���c4�uJ������إ��v�Ć2�lW���1.L>L�:�l̪P�%����@�/�US/A�1�%0D���	Ks�^����AI/#��U.r��v�=�N�����>�Q	��k��4L��-�w9q���9QfŇcg[no�Έ������U&�rm�lə���9y ؇j4��(�oY���Q�y��kŌp�+���B{�����C��q �� .�K�"����6*I�Z����[�ka�W�^��W��7E_��r����?�m���|y���8�>����no��O�%?#�l�u����6!?�k���!��[�e���438��Y(+]Q�9ñ~C=�௜�#.��p�o�/Y`�3��4z����,�o��nBT���4֙���?��B�Oa	�2T�pL���Q�F��~x���凜�+���&�'@��-�I�D®I�B�I�D���Iq���X��@zy6�G�W2L�~x�V$8'�v�?�쐪XB�#|��︧��KB�OI5�0(96P�ϼ0�c�3{��rj��<Ve���!S�RW���;|�&{�, ������@Sr�)��[(2o��&��w��_BdzH���k�j*2^	
n����?�A���	�������7{_�O(����k��J�@]g�����I|�� 4�u6����'�D��G~u�.�L`���3=�>>����r[pH���5�&�X3�ծ�=��A=p?yza����g��ח\��b�kw�}"ל�<ɞ��aMK���o0N��ϣ�.M��������#�.D�i��r��	���{�\�������゘ݯlx&��	���D����Ͳ�s3��T���EF��	W<�e���#5����c��[|��+߹[���#%Rm'y� ��I�ci�s����b|ܽո�5N1�*v��i��p4�������ƌp`�wyʹ+��ʒ���'4��۩���m*�+S�C�$��b�B�k�}��3Ơ���S��ϙ����N\)Jq���.�^�`$��Lwx^�_tŪ,����TJ�&˖�G��G��C������v����#����դ�-��kQ�ךy�A�$��N���N>�\���gwQ�&��k�8@W+�ػl�'�X��	��Kb;^oL��͹8eo�ocg:��c�ϑI��
d>�8hRDH;���$��{�o��9�<��Ta��p�)����������1�k�k��U�	!0�H�3 �3L�&��#�F�3o|���'���W����,.0bK���ҡ�OO\}#��F޷���,҇���F�Q���j����9�����eM���=�{;w�+b�;F�ht��&��
D�<�'N�e��j^Vk��ؿ�lw���q[*���.L8�[��]/t�-}��Sl`C�U�Sz̡7���<�;��O>nJmc��	���
ϳ	�&�T��2f�JH^=��w��:bj��V�����[ɌC�����Lk ��~�.1.�r�h�G#�Cg�	12|/�@�� )ة�]U��'s���>���y%V0mrm`އ��	�	��M7�6��u ��R�r������}�⯍�1�<�	 b�f��Ŕ�����P�Q�-vr��iذ
�d5�nɏvb��^2���Q���''Zہ;-���OO7t����@=�q��t(W�;�j�����	�� a�phDHEjl��"��_�G���;�!�ҊnzAh���@
�<iH"����Mn���s綌�B�?�R�э�$��=)�r�/�㙮��;¸x�e�[]c�D"��4����Pթ�}J�'�qYN,���$fߣJмD$�r�%JӶi���zH%�ē�$�e�к(JW�ݩ��(?�Z[�P��R���y�$�f��3��a[�?��_ŵ�)[����ET�����_���\�C���
H_Ie��ֿa�Ji�����D6��I�mQ�m���rgM�=�)���	/6?ӄS8$ES��U�V�D�Ub���V&n�p1.�wxaP�+��,s�$��o^k��hBf/��"����M���!�5��O�l��	�j-���C�bҾȪ�s#���S�~��j��I��_8��uXPζpDYG��!�RFvKO���B�S��P�)�=Ձ��(Jиm'���iC9z��W�!V�vR^h91�zC�A��Vvj�V��/�7�!5������?��Y`Ʊ�3�\@�u霠(n��	�%�05?mǒm�w���|HF凭��i�m��Hu����2���{m�i!m�R����Ũ/ %a/@�G����A�T@��c����/��:��5ޗ��v�5���䝯�\^k��CWG\-�u6����7Q:B$E�x��,s�6��Gו�J�9zwX$$�A�ɥ��>��W]p��)��Q�)i%Qض��GG@paA��u�q�P�'��%`�9ٯTń���%�P��!�ݠ�(�~h7�
��SY8�,��}.��Y�e\-��{���M!8yb.��uƈ�p�z=@�Y��f,�R�&d@�A�E������v ~������)�u��+t���R��.9���+�$�M|j���-���`��a������k%t��;��Z*�8��5B)|Uh��ӕ�xM��?�(��aM$u6�����*�C��6�'�V�E�a�<�`�R�E�X�D���?!����R�[��b㎤ܔ�I��]3<�y������8�(�����大��c߂��il'M>��S�����5H�t�%��Cg���P��#����e.�\mJƏe��]&�gF�$4��Q���O�(�`����*h5ص �gt�Yr��X��XvnEk�rz�yW�\�P�/�G^��#���1�Y����N��;�OG2hUǬ��i�Ձ+��E�۟��]�`�R}��9�sgL�//�>.'��*ċG�1S�T�<5���F-�C^'��oF֧u�1ǥ��"L,���u�|H5sNI��� ]���P�<8=��<��ŗV�,3>���~�_
���{�!�g�)�ݬ�БIRLI��U�pĆ���@�鵯���Za��X'NǥUJ����O�]�r��Ai�2>��s�WJ*O��=v��0�oF����\�F!~�E�-�5I��*��ֿ�nK;vn�{�G�����[����*c�̢��|�ΰ�)R�[9 ��)z��|�k�a�Uy��.g{�;l�`>�T��vM����4z߿�g�/���7&%���r�_��U����M��c_p�E�Ǵ�I&���G�Im�WmϹ�b*&�	�P��Wʤ�'8u��
2@K?���]׃Uޢ�2+��q���2�k�!=a,��F���ut��OIvH>(����}�Nd���~&���I�Ęs�e��4�u��m�Y
mZ�}(n���)ީ�	�A���0ԯ�H0ZNUj��P[�V��ǣmd�:&ݡgC@�l��(�?�UT��[/���2GH��3/6���&�����;O�p��
�y���/2�싚CZ3s�u�M�?�d%�t�8��O��Mw�m�%��t|�,R?��FIA�8��_9�����dJ���a�v[#x��Ώ�u�*���U�9���I	x!	�f�ʩ�z�h�'��.���Hwr��� iD�<=����?��J9�i�����t]U��S�� UK�K��T件R8TE2O~�'�3
r��I���>$�V'��^;1!C�EY�Ƶj��c�ڽo��%��S�RhF�*e��t�Ŋ�����A�W��`�A���!���5���:+��h�~�!����ۛ~�Q���� �c)�`���3Č�S���_Ҍ�
���µҖE��e3(����^�6A��s��7�-�~z�B�W8^MLѻ�R*5y�07'#���s�*�9d��Aa���E�����U�xs��&�3�`�WE�����B<����]� �=��SE*.��K%��?��0GV���XmS�♪��%���
w瞉�AT������� �<�V�}VN��bDm��l�F۬8�����S5֛��7��T*qC����+��n�5
_X�^��f�&"=ҩ!P���gG����jl����M��c��a^�j���}s�sf-���l��̽��w� I�7rM���^m�/���x��#!�t���:�ˌ�Zǚw�xy�7��K�UnI����~��� 0�0�|/N��\e�vE�θ�-�:�)L�K���z4�=�5J�d��n�FxN��T�x!E��H��7ܟk��	���K�߰G�d�D
�;҇���⟥�aV�!��>�PJ@�����]=_Fy�vC�eD�.�5�,��DKq��GG�m��aQ�MR;#bfY��s"̳��=�b||�<�{'A�g�;*Kr+;ZR&>9lZ�
�Z�b�%:d�-=������c`"�,�{@9�:���1{��_�{P\{D2��2����ۂh+6PvI
�$YB�8��:��T�/�p�/�l2��A#��������.���-��c��^�E�}{���m]'k45�!fS2�О(���9���t��M�	&�ӊ� X:��%��<w�Z��*�JYJIL��rg ���Coŋ鲔��o
f����Dkld���Ҫyo�~JW��1[Y�[x?MêOl�oG���T�%��f�JUTP;��L >`�~����&R:�X ��~p����ǕeT&B��g�ѯ�ҫ	Ĳ�B��bB�b�xlNE9��pEͽ���eW��B�$�a\&X��휂��t~�^��uGBأ���'�M����_·�;���D�G�g�\i�\,��,h���*�1۵\LqW�ٷbn�z��3ԋ1�t�o��Jg�Pn���pŀ�A_J��1�.�q�}�$z�]k����ɧ�Z��!�`�$�1&͚�O�Q@���ƫ��I�+7��cvߤ�g��S�
�/�ye=�$��7wa�$!�UU)�?��[��j�_z��b=��\2�<�����MϺ�ӥM,�dO�x���x~�ʞa�N���=���L�ƝY��TU�#>Z��ä�\���;l����3������_�U������uZ���Zy@��w˅ǿ=�M+!\��O}FV?���[��k<����Ja:�p�����0�� ~Wt�{v#������l��&X���,�x�<�7��B89�Dm_�Y�$���k��'Ĳ��<�'6H������Ǡ���{��z;s�´�ρ~*΄]���O�isc��?�׺��A��A���	�e���ۓ-Ҷ�}}�Ž_��=��j(�AK-ܹO��?�=Yٿj!'��n7�>'E��6�e�!B%�V�B>[�:���������J���20cX+�>���hpXE��k('��!f���a6�m?��U�U�M�ww��W����C�G@�k�Rhɘ��T��-�ac-`e�-f$���-�4��)���FM�/V�!�g��"M���1��K���6f��L��ƾ���BWڛuA0��5��mqjy�;у�>��7�������TWryգؗ�|oA'�d�9�["ԟڱ�sс���)���1�B:�%D0	�㠈���� �tL�̒n�P>7'@O�<s|����чo��~t0P���-`
#�'ۭ乲)8?��^�<����������_�y��o.3u7=%��7��أ:`��X������L�d��lS�;j,K�ʴ+bZI$��>�3�p������]�����9;۫�ù$�`z�k���O?<[c͐S�1���<MQ�}gH�Np��m�/��CV-�ח��?U6��,����Zx�縿��F�uk1� �\>�u$l*e���pC�=�=�2|tv�e��7zn�;�L:�g�2��S޻�``��V�WNY��$ޘ���V����j��(���6d%�ك��:I`kx�EL�ڸ/ȈF�������X�gF�KU�1��SE�t��z��b�bg39T^9����&&����G"� =�xc-d�2qrz�ӳ�[GG�}~��ȭPU��7�T�䅒q����bJ��8�?�in�C�W�p����u�,�/"���g0D�
�2�9�D�b�~R6�#L- |7�����c�Ym�l8h���x�tm�*QL_�M�u�M�)["����VIwğ����N슓�b����&��'�)p�ld���Nd�J�^������#�Y��<��7���
6�+G_0g��t�I4	g�홁F�'#�2�2T:Л�k���G��v#!Zd�+Χ�_Ґ �oc[�GМ'��g��_���z$��E��L�F��`��i�.�!�c��%����g�O0���k��f<�b�\��X�ڗϸ�)�I��BE���Ō�(%��й���7-�Qv�]��M7;��Bަ���{�"�$-��&�}���˫+y����$<�:%_��
�zξt�:��<��,5~Y�����+3>��1�J$T�6 ���m¨�>�J&x��y@Ȥq�haQڎR}��я�;��{�g�������"�i7B����`O���z��mp��TKl#��vO9)�ʿQ�w2�#ya"wC����D�
TI
pQ>x���-XV�=��!��x��R��j/�H,�U=�2B�e��v]n���K9�yrLƠ0�9�E`q�Pǿ����AZn&KX;��?��˦3�?��\�5R[�OeMe���øH4��/�=@1ܚ X�,�y�]�~�5�T����2!qG�xx	v$���ڒ_z2���^ϰ�=���v�Xۓ�����R�Z�e#�*͊���*�����w�>��(DpBB@y���g�3�Y��^�t�X0���)7W��v;�%���e��h�BIr=�����KH�$��_�݉.��ˈ�������O-{R~��y��5Et�푗lG�K���o?��-ɀDd�Łl�]� ��	�l���X7��5����jZ*�N�GϤ�9�/O7ς��P\ݿ: .[�����Bq	D�d�`x����u�������p	v��"�?g[�͇�3YHh&���ښ��P�:,8����*��$���OD�g�Y�|������r�NBU���޿����(�rC��{���S)�ܝ��l�����C��Ś��i��zk*�<C/�&��$�z�r�Th��E��W>��V^�r�;z+�޷h��`� �%L�ZL���|�ߡI�B++�Y���Վ�,BwJ���x`���XI��c��0a6};#�Ժ�)��Xt��'��9��c =S�{1׷8��m�@)����X�i��c� /���)*�n��ZM{�Wd�iI{\6¡�n�����@�=3G2S�A��_O?�ș�O�s�f��".�K�]�Kٴ�R����)<�~�VK��.�U�h?ݾ��j"��%���â��YV.��j �%��d�����Z2��'f-�7�� ;�/��RRd۽�+`_�d�"��O_��A۵�]��|��e:̂�f�sᴚ�
���&8LϠu��+��ו�����[��`"�����U�p��-v����Т]����۫�0��ţ�K��\$��L8x�o?xeY靟I���H�-y��1�7���ˏy0����X�,�[cC#��O������*Y�^�V�L��I[�J�d���i�vEl	�)k>3���f]K_7���Ȳ&d�1��� ����=��\؋\���|���$�y���K����4Ǣ�x�B�:�G�z�A��A���H�������>�Wf���*d&����}�z�杯���q|2���d�-IWQ�vU������W�b��J�,`S�*Yf�d��M7�h#�y�6�/��J[e։i�9</�1*9��*)ED��H(���P�UBa��VTUT��{��n8���ԘIQk��&���VC�O��;���߲� ���RNFI��FLm���0����jw�{����*���5X������(��^�i6�d-v)	���Ӧ���e���2�r��$)|�����5�_�q �4�hZJ��u��.f�&}��"O��m�
�� k�`u���T����F�"YcJ;�&_v�I/u?CTs�Y2Ӹ�㾬�q/˅p�`��Z@eD���Z��.���/a
w�*�n"�d�}���"Ms�9�kk��L��2'r�M殕���#�ᇶ�t�?F�g���)eU���*!��3,��cL����X	KY��!Іs�*������C����֔��Ѽ¶��5�s�%��T�"ՙdZ�oq(C�c�y��X,�壙7h��<x�WJx��R��MyY�+^��Y,��H!�����S1u\(�4*o�t�f�Z�	K�[ˌn����L�Y���Ng?����"����5"M�x��%9�8�N�����I���gZj�f6R�tE��f΅~e�y���	L!qЕA�r,��㫘�2�Ҷ(H!G�y�����E�VzlQL�i��?=�g�66���HJ9X-��d�+���Q&,����|��&H�����(&3�5��df�ݷI�%Ϭ��bA{�ï�^�)\�S�=��3����ѪI�hH�e����凿�*`Y#��'�:�\�R�u��N%=Ѿ.��W�0�L	T���D��P%m(��N�C�(0����s)=b�7$*)��g�c+�^�v
��Bh6�����$�?����X�s�p��ꪓ�r�cś�k�tշ�������gi�A��/ro&6Ȣ�����j��;�[�����`mx��1[�b��D�B�����-��&V�S�G�{��
9$�#J���?.5��w\8֮H�^.��m�%�)�,+c>���W�kf�f�m�3��4�R9y=(�y1%����m�y��k:-R���2�]Q���l[�*�*�r�T�Ϻ(�����ܠ>GP�K`���O�|
w9��E�ў��*�E�M�����US��fT���o�0�rm	l��jzR^F3���c�����_I��B�]���5G�4�Rpq��|�.y-�#�h!��ṳ7���Lf�k�p�ρ;�+b�������������8D���ڕ2{��e��ۓ�x���:�mֿ�"!�� ��1����mc�,��;|�Rd}N�)+��C	>$	3�t�|��MD�̶�]��Ă��"�`;Sf;R�u��%��<��cm|a����x�	aݮ'a���9&�SJyf�ڪ��ʯ��q ��4�k��}ה��x5;���r�U�}��1�h�Lx|���H+Jt���h��w6��AH������s�|4}w`�h����|v�q,��hY�q�P{2�HYe&w��~9U�0�L64 �Y��/@�؄���S�"���H��j����"ԉ?��vIw�Oj�!��9��,�M֣�\�\ץ3�m�kb���)R4��Nd�z�Y�Wju����5)��C��m�8{Cw�5�xSl�r
_3�KP��D���qH���XƆًu�q�¥fQǕ$�����������t���g,���^���/O��}�`u=$nb?&�V��<���WnG*�vW�mMCav^6H�*�ƒ��%��C��k���=�\�@��Bs�eQ����V��9x�#Yٟ��m��9�DHPv_m��߱N��51�'�,��CP���$�>��C����Ur���ݎ]���Ӷ��K��[�:q�:}UA!�Θ��h,����'7��4se�I/d��x.!��[��#�SR���l�rGR6�:���_��⼒nt�3-�-��z�'(2���5�O�獏��h_]�^!��*�1�������:�����;�sn#��/$v7���2�Q��h͛��}�du�����WY��w�p���	j�nB����-�ȵ���?謨��G��bn��i�-U��o���إ�iK�Gj�{	�4TD�1X�w6`2T��1'tO��Vx�ȘZ����1ĺ�L?�1,���
��鳷WN?��t������R�+,IYZ6�� %ˡ�ǾPj�v�:�Ǚ.sd���~W��pޤ��g��I��g���J�u,�!a�qB��I����l%�8G��{�����.��k*��$n4�7'�V\�M��B�P���2P�
�=�S��֧@*띘�޻���-��$��.O��ץ<�;��VUS�	����3��"�Pg������5�^r`���F��y�����>牣��4:��]�Y�Y���S�\롪��I��"U��F!攴6�9,��T�����0�����{J}NO!�'c7O��f�Ի\Q^��Ԉ%K���{��6�?�~f�wR8U��xv��1�s1��H*�[6T�H��B�Ew�A��㐳�������i`�>��3f��%�ȁ�;L�wM>����������l�k�����2��"�Z�𿑑TW��PK   �cW��*��~ ̋ /   images/243361b7-2241-4a0b-aa59-149fc34d5bc9.png�UWL�۸;�!k�n��ܛ��N��]���\w��v��q��ߘ�nV]ՒZ�SV�BC&B  h2��  ���_dla3 @��S�#Wv�3���	 �g&� (�i�/��Р�~K#u��A�����F ���)��k,f� ���5�)��Od!��I��|�.��ĸ7x������q���6�0����t���D���D!R
0	u*؆_jq��`���i��br�B�� �E��{>���;��+͏����p��	 ��J�D䑇M��z��܎վ��d���R>��b�}r$A�c2'G(n���`kD ����S���4"MR�����_:��)�G
�K���C@����g�/"�$td���ݑ'���O�����f|S�v,�.��!Oޏ8��1T��C�X�w�L
��tc_.�o8������-��L�냯w�)�5S��Yf���eTѽ�=f�\~Z� {�ǖ��`����ef�a	���,��K�s Cn���;�L���4X���lʵn���X��L]+(����V����#W*�2j�(�0���k�k$��!hj�F_�i�áL�M��p~��uvSv#�~%�i}�D]�˲,���˺�I3�������@�#�qAd�R\ec�\L�5'}����0�ȵ�nJ+�r�
�T}b�8/��Kf#&B��C�"��?� L����c�~�
�A��\ F��0��D�[Bl
�UF���b�AN拾'Ӆ^�Q���u���0�$����+�m��-9h�.D3��$��L��3��gY)T&��t��k��0�q�<���[��P��$����m<`ٞ���������k��=�7�m �oq����)&��8�VE�/<Yb ?^YuN�;Rɏ@K��<>�f�9�c����i���|��A���S��'SI�0�4���\m������X�	�Q�q"dq�FYSqR#R�S}ǽ��zҍ�j��x����������W������y2�'a��w��%Z�Z�Z�[tZ|פ��C��^vv�����H�0���P������a��ъ�h�.�,I�S����H�}W�C`�O��U� ��d����/MOo�$#>
�˔�)�3\f��"��@Y� �Pn��iip�d�C�U�ZE<�=���թ�����N����n]ճP^�Kݔ������P���G�ln�2�w2��p�x���oj�jH?F������G�~d���唉4*�T����J�L=6p6�4D4��%��̨���*>פ���k7�`7~m��t�7���6CHL E�	9�;�v��Y���x�A��������(�ȍSȊ��c��ۂ�Jhᛕ��ļvE��I���3��+!5{��{.���y���F������PD*�^� `2�IlQ���[�9Ẩ`zvq��]ĆV'�<'MF�d�a{�]����g�[�;)4y�<TdT"42bl4�`�`�UԐ��HSbF�2nOCyS�b;�s�wCcKlP�B��nki0�"�a�6�p`|�a�b�4�w!�g�i��k���I���O�>�&�&\������#>5�z�}A��O�_�6�ӍH��׭�F�i6LB&�u��Ϋ>Mg��N�O��6�t�n��O/x�I^I�yx:\�q��O�x'\�O��o���׶�w�����"&�A� =ׁ��*G��瑉eơ��U�s�s�s��[uf��zN�?��p��պ�v^x1pSv�yls�xYuGf�Q���T�m�S ��_��9�V�����-�U�M�UzE{Mx;y�ɄN��D釅G�E��߾nuY�&O��$zֻ��5�U���L����i�r��p:H@J�����w�:;������ZY+��ٟ�7�)
<	�H��G8�_�����y=}��nC6S�<*N×���Z��u���m^��=t� n��^�G�(Usک]��{C�,H�H8]��<8;��m�F�	�tG}�n1.Q�z"����!��)I��b�&�����N�����aX��x����_"��r8x��Ǐ3�HS@�V�9ВLŖQ�t�A�z�4/�'i:I/�ArߓCSt,k܏D��6 cSc�c+�'��np^�IS��I6����!��5�-|6wvpMp?�.�+,��ƙO_�l�<SRXLw6�[����>��/�v��j��W]���a>y<�z7yPP�$,���o�XQ�滃h�F��^�>sA6��ZM��+#�����7$�hVi�K͗m|v��ʽˈ��/h7���*�6ډ�\��ʅ/��Ηqj�K���]��7�^�\^ǟ[��˛�O|�|��/a�\�\\1lKBN~���n�Xz���ї-)	:²w�`F�v��&���R��ruE
4ʦ�*�M�M\'�$W%�W��u�^-�N�՞��˳6�݋.Ǘ�;�)��'�9V:s���N��ϜV���:�G>f��]����R������X�pX),fU�<N5�dMf)p��6�9w.�p���3V�ؽlt9�x��󺵷�y�Ot/�n�s|?���1n>�%		1����l�M^�vvu.�H
�,]x=I�6xF�Q�N�8D�l���܏�`~6�ՏF��Vz}�aZ����x�����8��[��n���io���^�o���>�<]� ��!�9��~�>����w:��R B;;�{97
Hui*H��sC�Of�a�_R�/s���1� ��0�l���v�2,.QM��d��t�p���ۣ� �wMט����&�ϯb4^�����;*���w� �5�I��� 
 ���ډ��k���m{��}$��)��UM Å��#B^��-~h�cC�۟@�od2��T��|���Q^I�:��^i�o�{Vv:x*�=��AT'N���4�o���Eth������������A���@^����7`��qwk��004�!�)�---�=::j�-]�>x{+��;�}an�ya���Y�%Vf��}ւU f軯��*KU�TPXUXP _TD�s��ؠiiy���i�G6���ֶ\y|��I��ކ3��8���b����l}��*�06��2qf�Ȭ�����=3][Kv��/'&�*IKMeHώދV��9@J��d����+=*�[NK��M3*��������=�qM�HE�O��{͊O��?�ȫ�Π���x�"Ǩ�ZX�Fގˀ_�%%�==��MMM��M�������+*�O+N'3�2�OOO���~?�ע���C�M��m1�'{"<��i}6]�h�����������㸸8
��v���{���Ɯ	���1'� ���i��'Mj�<{={���w 9f;;;��Yi�z
L�pY@N�M��aU(5�qy8�w47��;A��R�]�ޗK]Ym��H��-'������!v6v��8g����{�������	�؜��̜�Ռ��O���30�ͼ?�����a�ߓX����鉢�$(��M�=��;K���Ά����ܧ���'��[��C2�۹�W�et?�F����;�=&���I�����"�����n��}w�x�M���$FR-r��*���,ŧO
�����l����{��ۊA��QB�܆�@�����1��4]�F�%�$2�Q"�w�o+�������Rr,�[>�6�7���+}|���:��jr����>D>�{{{= N�M�󧄝������T ��Q/��,��(	8��iA��� � 0K���艖֫�IT<�J���u$�����p�����KdY<�5�P4��N)�ɠ��*�e�(N��(�u�w�9
�ӕ������6�v��٥!�C3S�n��������Ws&��k:����2W3��ԍw������.���gg���]+�[����)}��ֹ��쬽��ڍ7`rL�C��gbc��^*J{�EX;��Y�]�r*N�N(����g�0�FcƗ���`�_��zJ�<��˳�ɿ�|U���B��V=��� �����`	f���Mb\vk��P:�-1�������\_�0�>�S�/�� ����X��22䤥�^_�z Æ�9P���Q䄁�NH[E�J\Bb`g``@J.b��D��}��l�� B�-ޢ;�:����ҽڮC��\�]6f���6�7
K�5Ф�nP�H<�=:3�މ~�ϦsQ�� d�@5�J.m,�Hag=&%��*h�K���*~���%2�m�b��� �΃ke�g@m�_]���q���@���5)H�Èյ�0{%= �ZP���V���u	�"�sY�}�C򰐞7�>����8� g�w�i))�lhy5��2���Ĭ���Y_��Ϟ)����C�{�O����oa=1��8i-%������~>�M\Bs2���Q��WWa`��Ä�~j"0{�BOS[�?���D�K]���_9G�-�#��v�N���`*����Lwkع`��q��Z}��0fs�	-h��w~58��vu����YO5���w��b�"�_�r3����0�=D���F*����R�fl���'%��er�m����c��$��v�����c6�_!#I��;�+d,\��s2�x>Z�^�bCS�&��f7���oi+k����k�Z�R7��a�*,�#�~�m�<���YF$k�?���s�)�K��%��C�F�����Pڥq'6��[��)	
��|�L������u>��>��I�jO\~�z<�!J��A� u�>��:��b���@x-�J�MA�W��䇉A���h������2�	������٬o��H����=�����֔�1��[v�SK�zk+ӵu��w瓓U�m|����O�|���G�\���$OIj.*�$΁Mu�$�����pi��B�Piƭ�l��pn_�øθEPFC�%x��R�u/�iz�ƃ��S^���&��r�q<=O},&�.X)I���ESe1�Q}{�Y�بCC�q�C&e&Ui�<� ��� |��4z��s��-���p}{����*^��"|��T<Z�*Q63��C���s?�c�T~<�Tܻ��*s����Νɦ��111(�3��GZ�L£�6BQ�M7k��+:�ߊ�\��4�u�LI�X9�q��2�B~]y��m鵙��!��@m�<ɽ����W�ːr_����e��R 	�|Ln>��f8��}��W
������U�+r'S��%
��W�۹�D���}�����Hdx���4&��VTRY[{E]O�����飱��vic�F�d����0��ַ�����0O/�̛��^D�bwke�[�)�������tV��}"�9�*1�]S<ԸB̗ !J �p�����>̩�hz�e��)�(���;_Eu$���ـ����g��̓���xe���b��48+$����N�-k�,�w�lѳ���F`�1G��\;/\/G����):/a�q������BخI��y%���җpȸ"\)���mlF
1���m�O�~�!�M������DK �e�?�3���e�ɁS]-�_�� ��vr3;��>T�:�¤��6$p�r(��1�Z�`��iTI�b]�ߺ�l��iU�����k��m'(��U�0=��,�h-O����8Q�g��<�[}F��8=�3�Ɔ�� ����/��bm
q��;0�_l�z4�+�%@?��>b���\��,�x�������X���ed��4�R�������T��éd��`��P�q~>C���
����6��*�E�>�����!me�P/be`'�3��C�����蟟��D�Q���ᷲ	@T��OT"��M�n8�t�4T\�
�a�u�l�dA�r�i�G;P1G���F=��������Vyn�6��wF#r�\� 'L��_��l�>��O�.���͕xH��?`�.O,*�&C�Z��D�������zz˩�8�0Bz��8��}%Y���`���9炝�`�x� ��m3�R�����������f��6��;��@n�Z�������!���ű6�OM��E��OC���/(����ұ`~�Y=2猰@&ݚ�`�85�[K��H-�8�_����fJ����/���]/d�ݍ���UA��W�Z+3���d�~!�^rnc�M�DrǾ���rz0��٩�c���P}6m�RB��y)�ǚ��.9�@���o�u�c�5dݨI����W�%QH�#[^��x��$O C�i�anU�)�a��C��H���i?��J������B�LP�� ��B?\!0�inij �vN�?���k���*xS!�NI���C?�P:�5��
�{��Q���t(�V�_O=����K�����q���!kg��9QVi�Ɣ���9!��sZȬް`��x,�}&�X8�Q��zvw�K0��;�k�B*9'��g)Y�6p��dV|#}��WE�����>Xd33�*.d�A���ޙ��,�ɖM(��� �C;�M7:~�T( " ��M��Lh��Ա�c-lP����O��c�z}�A�!�jt�"�g� �=�Hy��D�A9�4��l���Z�XyL��x�Z����Ady�"�Q7(�^��y���X3���T�B��O��4���J��42���0�yX��"*�lh"�p�l�`o��x)(_c�cH�O4��߿��=gf���Y�/NN�ߢaZ�&Y�BW�k9K�a�2kO#���?��JѴ�d�g�}o���"�w�����>J���ˤ����ˆ|�'�}s��������:^;A��".-+�v�8����={6�`��*��{+���:����pU�?�Lgfi�I,���M�dF��)�[h��qE;Bl�i�LR�1sE��I&@�9o�
*W"W�\2U ,�	b8�UC��{�Ơv-[�@��1�YB|�B�QX{���
sU07��c��g���9��u�-=,[�}���c`cl��K�K�g}��#�z@��e	yu4��뻵�N�G���lV|(�[�/�q�7��kRs��2_�+E��
�тg�}�	!���´�̄�5��}���I�ɶ�B�W����y�r[R��:�U��N�,������|��M��%=�7���^{gLy�=sNJ��<-ȇ��lN�Yk[��cJ��<�R�))º�욏�,L�a,�<oO)��^a�Ol
_�d�}�Q�6A�8���{w�M�j�w��>��-�Y}a���q�09d,����_K�e��ɀ�F��� !�wKv������&�F��y�}r �EgEX�
�:�	u���3`K�H��wI�#�-3��Ê���yI-�{[�i�)9�C�߀����w�����d���B��f�|?�|Q����t� ڐv�_wc����FW]﻿a�4O��ty�tPȁPx���w�u�4քBk0;ҡs�rwD��KR�/@8VK��}��j�l��R[���������������{�&p&ˎKJI��}ޑٰ[�J}�׏���Q��0�Q�^�V�=���7��%��e���;�ž�q2��SZ��w�3��%�	~�f}�7�Q���q���s_`����n�/њ�qў{n��;z�,$4����(��c�������'mhn�n��7`_ַ��vw�qV�	������拘�h�T�����ۆ����wF��<3� ��Q�W
f��B���u�-��N�8���C����TW��lF��@Y�pt2����sU��V9 $�U��l�2˶5�g�=�M��Y�{<�i�Й����=idp�۾Yj���Q���BL�ұ^C��.�Й�i�9[܁8����/�(�8甆Ò	��'�,��yu����<���$2��Q��v�`�F��x���K�!��J�h���⧼���������u̫����%�������-	�i�z/y��@ɴCq���A���w��ܹh��ޜ_]�c��jz����0�ݙS;0a�����+XV��-9�l���� |�eF�b����>|���׊[jdS�Wߍ	�����a�ʵe����~z�M���mĐ��	�L�(d����]���q���F�����W�����?K��b�_�Fq�.�pHN��ͯ�-ݕ�ҭ�A�K���������ǫ��؂��������$'��E�-g��'%.��K�q7�R��������t�؎O�<b���c>�i�!���T�9y�A��������@�M�B�@���I�ī[%p�*ӛyj�h��YB	@��F�Ŭ��/}��!\Bf�:Cu��m�X�:��/�5Ģ-�� S���A��;2�L�Q/�+|Ϧ�)�����R �U ������Q�H���C��B�{#��bApڛo�5�gRzj�$.#|�:)h���?'c�&���]UC�\9��S49�c5Ԧw�y��.Q>��;��`\�aNҒa5�������J�Rf3_�[�2/C9�$b)�y.BӅ.����+C�P��	+S�=��ޏ�˫<�:��F����=:C����7�A���nyu�F�ۅ�����	�&�~�X���VY.ש	�,��b	"��@R�]mI}�k�y&�I��F	��ޤ�b��<i�ñ��T^E
0�Ywf�tHDO=;��}y��;\�._��C��`�2C9�ܧ�Z�rx�
��,��X=����Lu�R>>�qo9��
WƄk���g_{�\��zP�,�̳���勴v�O��}��ŋ�˿T��C"׏W\�^��4z3�S���Cv`�s���iTO�U���xo_l�7:��Z��.����vK�9xO��uyZ��������\ƒ��9��������]�jAh�n�[�}!���z�DQ�G.�2P:>а��	$���f��{\���MYIPؼ��j�hM{g�s�������J��K�L�uG7�3��#\"c7%-��c��ә�M��r�
B��K�'�W�����ř*�ac�	f��$��$�Ba'�#�!H����?�D-���;s�hB4n� �~[�wQ�ӥ�b17&2_z��R�Ub}�|X�*����Ŝs�Qj�86����z3��^�&�S�y�k���;/<;x�:����8nDt�(�3TK�f(U�~q�^���u��p[k~,��L�ȝ��*���i<y�sa<g4����N�2=�����eG�絙|���/W8�����:K���aQ[�e�W;�o�Μ�s�J�!eH\��!$0SD�x),���W�<�]
�9�^���Pvo$0^}
�v��Q[�*w٥�Ddl�M���T&������}oC��f�J�f%���I�}���7���U2n�92�m�6�LRcya���p~�� �ha�c=y���E��BcK��?�c�C�/K���<�3����b�r������254�@�������E�`:%'���t6�~���h�$\4�2%��!b�;2�>��SF����n����Y���ޝܢ��[�Z����ɻa�~\tS�Ʃ���������ΐ�� ���'�o�p[��q`m,�0KE6qx�����2� Ꝋķ�2@r��kq���D��G��s)4gn`��J�8�!�Q�t�剥�(���n�*y�IQ��E�)eJ�g�b�`�1I�e��|ᛷ�0Ӳ5b��
S�.�������
[�E]A��-�Eɕ�E���̺v.�('���:,����6��.�z�8-��Ǭ�7�F�'=*N��s�S\��7�A��P�7Wݜ��-�ςk�$V6��!?M9-5�d���r��G�=b����2\�q���>*6ѓZ4�ݻ�&�˵�r)�EĶ���k�/ۭ~���<E���x��6��������1N�=.�����g<m�44X��@(�%��D�'|w��Z��ҕ�sV6�4��H=��a	��Bp�WQm}�6�֒��N�˖	EڅL�����:|����p�6�nq�'U�7Q��x� �� ��Y�&���d�u��E�J��0�_Yh�lx�Җ	_t
�rJN��"1�?(L�XςV#��/��8
]��I��r����¸J���1��ɒr|���3�<�Ƣ�M�F%G�M�߃�X2�X!^��	lrӣg����(b����2��R>���JQo����\;S��o&����a>�do5��J+����Wy�y�x�LhU���r����-�L�X05�s��Vz����C�:/���R	�x��w�/p��U���aC�-�����6���(��;$��1�{PBO;'��@ޱȚe-|������W��F���+�*9$b���.N��$v��߇������y�}�v��7��H�ϲ��b����NU8k����"]�f������n8� >ݴB���wK.\��`����ó��x�|��2fU����Ύc���D-a��4�_��P����W��Ͳ��z2�"�L�B��Ǝ*�����ڰ�R��L�!���SnOJ�f9�_�,�@cVk-ܪ����9|0��K�}�$�P{����qw�eE,��g*L9

�e[�Gt���x)���Aܦ�5G�3Ye_U=�d�U=������C�:aZ(����fl���?�5f�"�W.y�Hg�v��=w�����˙K�]ĺ[�>������f.R!�[����f�f��[4�>�Z�/�|�ڼ�NL�u�	��zNls�p��C����������]�p(����7���e�T�[��|θB@� �\�i�%������#Y--�������ȏq=�kNK殃²I$2��yzJb��8��o�MM��2O3[[[Rѹ2��8�2����G	=o���������&%�! %� �������^]i�V�)�����Og_�r~����,FHy3ĄK�H�p�Pakk��R�y{m.����8��yŞC�;�^0��W!��ܮ� P!Q~G�� ������;7l*1u�?|5�a�yZ`4TK�;<�6�j��4=�kTvSx��.��P���@���l8��ه�M��l��������pq]����*O��̛�bZľa4疉���4<�9b(��F�A�KN��_�F9�v����u Y =��R[�X��V-��6n����
+[zb��p���#<�����+UO'ʴ3�y���c�h�c��.��n��1u�a�x�ր?\z���E(&�Ԣ!I7Os�K]c�lm-jm\��܆j�{HA�G����uY�Z��&����O7�gĈ�:���گ�~���I��d����n��A��|Eŝ'͵��PԽ�dg㓌j�:��q����4ߏ}Yو@	|�A���;?����Y�nL_j�����K���Z�[�������3�8BA����j��$�������x�OajU4��9�I��r+�?;!DZ���:�`�;k��2lN����-�9�0�٭�I�90���N���)�)kjz��_L�i���PrJF;;���I�ad��u�\���҅xj��}��3�3,Q<?p��ӫzhgf�j�O���v&Ξ�
 �Ց�\xO�ֻr�z>d�j����dx/��&�~kF�H=�5�w�I�j���*��|mM0����b�-�8j��ʝVE��4䰲uU�ѹ[�l^�zXw��j}���9���w2����x���걧�cz~��5�]�ydD�3t*%� AR�Sdc�Jc�ʪ�M�|�L���F�R�N���]��(�K]�}�O����C�a����(j���s�O/�l�M���jvea��0$�<������S}�>>��8�WZ��1P?�^�]A*$%<�����z�p���rw[qzv��k��fb�n��_rǓqL �8�SQW���S:)j��|�{kɤ� S���/���r�B2Z��9_��%v@,}?��l��i|���*m�iWEHE�l�b�_��@SrLE���%��/��>��v>�7NO!W`�?R?��7�|�^o44����Վ Քe@H�!ը!ר��vnCH�..ՠ�$�>�kJ�۩.�f0`����i��2!�׾�2҆�Z�>ׂ�2̀�7�[�'���)���	!�v��&��rڄ������>#�G^EG�I=7zV~�V�G*~ө���Y���i\L3:z���T"�S�"�'�ޫ��h�QR�4���#���U|�ٯ�=X����΂Y�C�ǯ��_�J|x�A��3.�4�����Ĉ��&�?\o�]r2�:�G s(�ׁmm+}{R�oB�}�� ����Ha�=f�?x`����0<��7����yv�!	�73��QT��h��=Y�i����w6L �L�#;f�gh���+y��B9v��Hp�P��l�)�!["�B�X�$�	�KW{JD��`��F�(�s(�#�������ت��rC}A�ai������/ˋ�������Y���a[cg��[g
�����(t)H<�v��4:V�}nY�l��[�%	z��Ӎ��[C�sz>��s,�E� ,������}E?��>�aYZ=��-����{:`�׾
V+6���ɮ��������&��R�v�5�l�`\i�_gkM��ෘ\������ྛ8��W{��
:���q�͚d�8�Z-�H��Y>��"E���7��G)xw��w"��<w�¯����^�.]
?�2�h�$�R�|�^��ڟ�N� ��?�l���T8��$�F��7uu�����+�,��N��ܙ��0y�u�,l3� x�PY)��׾�����x|Y�SQmh"�?#p- j�� ^��Ȫ�;@��@��C�?F(Y��
���
u<_O)����V�pJ
��������?�J(�ð6_���A�]C�E�k~��y�{�)��.b�j��D����������\�惱���%a���G�۴!�W��`� W�"XǺ���iq�'���_M�����~Ms]����e����9��5\&I�cs�g��s�X�ю�A���G���#�[�UNb���4��Q)!!Q���WQ�v�;NO�Dك���~-��w����8�|�N��{�{u�%�n��G0X]��Uf�=�Mhȕ��k�I*���n�v}J�'C\ƕ��l*) v�����ߙ������r��u�k53 �1v� 5?�p@��h�����'~�f$�0�G��bfu�P5������W��'&�/N�b��8zJ�a�k������>��F��Mۃ���l@`����L���LƟ���c��P�Q�ՅP�2�r?W5�(��e�O������M�aC����z�}K��^}YfZ�3V!�W��\82��²���f���Nf6{�Dx��U�+��I���'��$8�Rd��%$o^�s}����� �@E����k�Dg�M�Ⱦ,�F�F:]^�Ȋ�l� ��C+�W����&��]���qwCM��"���6�Kػ�k��r��PqǦ���I|�m�'_;�1q��&@�<�\�:\�{���gǏd�كqFYmU>N�a�ٻ`F5(�O�Ten�n�V�o%�(�=��L�4{82������j�(lY�k�ҙg�i��cc��9�**W �Ʒ���2���='��Y�OU�ve09O��+��E��:���S�no���2D$��W��4y�as�Q�"��{Pv���YB[��]�+�_��&nY������V����X���]�W�l}������S���b���`6�~Y�[Jw�0�����^H����?���]�ϋ-�D��v2TT��o�L�\���>�2�h��R�ɤ�(p��b%9��0U��%b~`r2[Cץ���kU�l����Ѐ�e.'G�����J��ApOp^���d���...'{���>�fW����7�k0R�k+++��"v�h��P����i�3L���C
6��y���$W6u�{j@u!�-�����*Ԉ�B�DZ����v�B��ާ�"9ϯ+U���{~���7�-S!�"������b.�.�b�z���iWEu3���ǟ�	�)*��ȕ=>n ֩��>�<�dU�$�<匱VS;G�&��C�l��vƓ����/�������2N�z�>�tNHN�ӘM�F���F�&�������:Z��cȖ:p\�tձ�,Ղ4����,��.*�U�͕�I�k�&�r� q����!G�u=`����J��CH��U�gq����E��̰���R3e�2�ց�޼���M���]g>�+���k��P����Vnmy��j4iw���;F���ꌎ�����R��:G+�^liUڎ�����֖��B91��(�� y�yd �C����*l�TT�c��u4e��Ul�g@	V;�֡��E�]�m	����TWyNJ?>����h����:w���Tu�x=��<O�>v\�K��������R�n �FN��E/S�C8�^i�hL�B��u��
�@�Ƙ� �Z�qyl��>Ϻ�b}]�q��I~��;��#Ҙ�Ua�䇜F�d��������'�!���������hb�����D%�"�X�g��?h�3��Z��J�Z _cuvq\aa	����IH�Aq\`7QŪ��yy�=�qqOR�r(*��O�>���+��o:1JA�^mr��:��)��l��}�����������M���Qy�q�k�q r�NR��b��O[Z|3�*#������ߟ�JczV���w&�~`��U��ã���;Aֻ���7j��Sg`��j�>��V�3\��e��4WW��0��<���p�#�lyP���xcu쉷0��h5?[��}�*���Q��x�d�����\��O l>�e��
�i	��i���u߷�l)�&�B|W��(K16�l`n���y�R�޵f���iZ�� �b�Bk7-�e7���{�j����C�}�l?za>���o�ďo$���}h�0�x�|�)�묉�J;�� �̂S�Q�/6 k��G���ne�V�[�^Y��}�REZ����W���y��;/��I��E�@n���F�w���u^~�3]��ڣ@=�,+ɡ!zL^ܼ� g#�a��� ��ا�ϧg��79Z���)���;��H�K(�+O�������7�/�{���K�bX{��p���b���i֒U�GrD#0������2�1��Js&��_z�Y¨��H�Qq7e18���c�*J�U ��;SJ~�%-�^7'���'��?����ޏ߄��K�(����$�IxÜv1�	Kq�
���bw{\���qmG��4_���+���(����#3��d�WDa��5�4X7Z�|R�����'�ά���!�k�hV#<���!|wۆ�e���������灙��$E�T�S���"dӱ���ʖ@�'����J�|ٜ�X� �X�>.ϱ��hi�nfn�.f&��!��U�rj[�����[`)d�����B�Dg��9Lp&��%��ۙ���J�MF"oF-��^ք�*��O;y��%\n��y���(�*�j0|E�k��Byy@�[`�|M^�mw=��S�^�f�©]
�]�>;�A9L:uз�F"A��-�Wl�TKf��6����\r#L5U�zd��$݌W��\���`9-D^�߃}�*τO��z�(�����Š��6��O�M�2i��S)�����ôƙ�z)�)O���^�F*}���'n���;�9咥�.����R����wUn��,b%��]%�f��"��T���P����k&�������[FD���W|?3o���U�o�j�j`eֵ�M��>|�Ȃ���s^�U�e2&�%m�w�l�p�N�/0����v�6�=���`���#�64�b�	F0j�ܶ˻�AӦ]b7fpA��QմC�Jf�l�q,�2QS�HVڭ�5��ȴ'0Hm�p B��tMؽoUw��|�}�s����Z�_�x�d&��o��%(	��w�g�!��$,Q�5�2��vܞ~�K�lx�|hgqJj�#���:��X��֬�C	�H6��/}\����%�,J2HwW K�f����~��a+���9r�ţ���$P���*�ob�}��,h���Yf��ʷ��� \�vpAA����ݬ~՝�E'>�o�L�*K��>�Iu�^����w]�"~�2N&Ԭ���j;6��d����>)�c������-��8����9`nͺ���5��	����+晩�(ָ���8�Y���:��M&�ߝ�p�d��0�_��[�vf!/�w8����P�?�'��T�XS� 4@˿9yJ�R8�J���P�
D�jm1a�+up�L�JJ
�1,�Z �d7����#΂��qf�$GP��pqXQ�D�u���Y��r��E� ����g��y�ٹH�;��,D��z��� �����E�����3z�[.��ٳb��|�7<x裑���#C��O8ANxvÆأN=�e�3ke5��֢�N�:Tw�KA/��U&��*?��69;-(�*����/��K���Қ�cg勇v�_϶���/)<�Ҧ[{��linY��\��Q�|Q8�i�L�a1��ZG55����Zh��2�͹hde�H?�8"U�P�OWg���ԫ����7�"s2�w��i�K�6
�5��t���.��"�Q�7N�b��͏f-1'/��@vs9�f�ǔ��.�_��w�|�9�Z.�����������3G8�����RP��)�,rɍ��$��YJ���9�;��.�D���:e��p��3#ə�5{�ך�u'_/����ݑ`ώ=�~���	<������l[�������~����+[�����ҕ�B��$Uc�f��L��"�>��|��2�� R�����F�q �t<�32a���H���T&�љ��V(��6MVM�{�ÑFxh��p2�BR��R�7%I.>�)F�3
OC-uq�Pg�����D~nަښ�Z�r�O֯X��߼μ�~iGD������7"��F�2Ǿums�
��Id�8��)xF�6m��PIY��svտ�<sk�������d�J���AmC����w�]�z����}�~6���}�X��_��[���|CO2�D�I *Y���3���9���S�N�JX�X �x&���0����5ג�O��6��˄4*���`��b5�v���򠴼"����",ߚ��+��LxZ��h��E���m�<P�M����NIV���G�r�yy��災��ǭ�55_^�`��n���.���<}ћ�Z}a��?GgFoS��{�r�2"��[0�C�D0�:�4 �e�4Y���mc�}Y`���&�$:F��8�3t�A�����cfBW{W�K/�����_���e�GΖi<��-���^2x��WW~�3�����±a�{c����p�s�(�6��j��S� 	�|YC�@����&ud8b���s�͸����$�8t���%e��Kc��?Q8vzX,#\L��j��mhI�$��F����� �H��4�7�pd�C(3Ȼ�*��ohh���7\�tɜ���w\�a�՟��o<�����Q�җ�y~R-QG�j>]i\\;@HDM(Zt.׌8��i�=~}
9ԍ6r)��y� �FG��Ɩ�^ٲ��x�WΖ�<��-���^2x��'������v�$��!�)<��BP����8���'���A��F���:E��4����8�i�a+ ����xOwW0]<��l�O"�����y�`�~e� g�8���9�t*X#�;%Z	�C���<��)[�t��/�'�o�����޷�����ν��|��F��e�;JR��@��v�*�)I@{f�,��.8P*��h�sQ<m��[2������mٲ�O~��W�x�m�φ5Bc�����>�.n��w�@�;�Qr:1L�w��c@Y''��dF�rG$��gSpHz#�ݢjc�sW����d��{��g*�ul�ly��ٗ�;�j��d,�:'2݅���0��;��Iրiv]���q��	����ŅAaa~PXT�RW[�wW\���o{�Oy0�����۽��۞^�t����+(�9�/�p.�B�<��� �w��i��m���Ll��8��+�f��ѭ��8��<���O�ǂ����/���oٿ=�l��G�gê~�����?��S(.)^]�_�w
��cA�y"C���-D�3IL�ihQQ!�^s5Il�҆�9�̥O�Kը �6x��4L�˴4G���5{,($�1�fj����q9\��Ӣ��>��9� �
�-;'G�	��I�-���߬�g���������\�|�����%q*�/9�-𮷾�o����;x�oQ�� �\�ԙҚ"�E`�]!��1�70w�N�f
�a����*H���Y�Ɂ�ߔ���3�Hd48r��[���z;����6�g��i���]�غ{w�����?p��;:;߈:#�<���Z^�T�"9��;<��XS�iD�d�J
��� �A��\L�h�5s��K��ԶH�
8c� 3�����qQ�xG]x��HV�Ǒ�t��������18��To��K0Ǡ��Tu7��#���WW�YDA_[�tI�?��`-���O�߳w��::;���Q"yP&�A#�1�\�u�]"m��DUf���M��Ԕ4gmY��=� ��4�ˑ{±��������KV/���w����\�y&��#�3iM����/n�R�e۶�~�{�34�7 �˓q%�d�֗!�u���'h�J�k2D]4��F���i.���:C�V��q�h��&�[r���~��1PE�ଽKS����\��Ԯ���F��BVDj8+��&5{��kt��d����)h��ɤ���X�2�fWpG�=?`���E���[oz�������(,�7޼�'O<�۶�~N��LIq�J�D����w��r�Vb��9K�h-<y��d
����=	.1�#n��:e�p�QJ9	=�I ۡh~�L0�Z�ۮ����{��gϤa=��Ik�}]4�C�:m-9�%�ut\�s�������A��	f�'��lFތ���?��1Й��M���qۑ`VT\,�^���f�ˈ�}�6D��#�� {
�o
�	S�{b-��.'@۸T�RG��YF�-�%�s{7֔��4=���t:��8>��І��,*�o�H��?{�ez.�����w�z������?���E��#���iw�ƅ_B�Ř�"�e��]v���kR�Tګ�7:ͩ |�,
t ���Yrg������v�����^~��7_y�SJ�)�����_�d,��Օ���9������H�m`��G��SM
P+.�B�J��Ç��o;*D6�=��m(�a�+b1���.irz�ne���%E��d�� '��H����)B�ӶM�?�9�ON@�׶�}���I������,v��]Zf�Sy#�K?9�px,).zdQ�¿�h�W�*�/4����6�s�����w�ȱ������	�v��1�2s�H���6π�nי��9 ��J�Kќצ�6�D�i �%�#C�lWM]up�m7�ɇ����L��������i��{��wvu��������U�##�ãC5��,/P�j Y3..*B�u�l�x�X��އIgd�*MA�����nCWb�5��d��Hq[t� �57�N��锨��΢?�2�F��[4ϋ��U���u���LK<�`�����7N@˂����ق��<=�9H���TUWu��e�ܸf���/�3�t�_�w��O��t����炱��a=]Ư"�Ǝ��#��ݤc�zi_��u�W�h?�S��N��4�`��2VAq~�b�ҽ����wݰ�ڦ3����������g��{�,����>��3wAo}Q$	#Q�Ç��>)d���Q���0���z�$���]TX�Ҡ��"(�o۱+رc� � &�tz���Ҭ��g;e��OsL�E�=%�q�9ר@G��V�6��MF���!nL���YnO�DHo |�ر�-#+���[@<�NNbP+GK��(��kV����������;����֭]���>��e�ԗ���g���@��z��_{�7a��m����M��(������[�n�U��/��/��LX��ケ���Gj�����g�{��]]�Q yt��vEj{wJ����3z�d�tY�N"a J�wiqOP�4tyEe�v�ZQf۲eK��6F�3k����9��1&��o��E�<��3��u�n�t䪒w���R�6�QS��;ǂ��5�k�:�G����>���3�V'�,v�����̠��eK���[��j��C��8	�Y:o�ٗw|bh02ob|��bPu�ML)�e��ǉ�H�+�]%^���"�6�)��������OHwt��z$�6P�T�Ç�{��Ǿv�u�=�C���x@���`,���헿��϶��_E��m+����>���`L�������,%�E<t��"���y㑁�` 2(�� ���o^x��`��}�m�V3D�J��L�ŀ�<���g���k�%M-� �ю+��f�ysLU������X���fB1H���<��`�3�^P���S�YYY�o˗.�{S�`~h���`��\������	��u������6,�ך\3�Ŧ%0�[�^�P%V#�.e0G��vT���b��S�N�$���Pu�]�o��w៟:��~�M=��^���ytG#�۷�x��/��ɮή����zz%2�Lr�ʐv���N����� >�e3��7�l.����~�@�)--*����+ķo��!���f�K-�m`�G���ǅPG"�͕`G����b�m�]#т��\M��۴(�X���f����b��|�!�����:��l]�h��׮^�ú�rO|��g�?��c�7�v�����ѿ���y\��]���L��>8݈�90�L��0�!�X�ZDW�	I�[�V��x�#$������|ݺk_7���9�{�����<��S�6��mo�(��� <6&�� :ъ�q��y����^q�,�d^Sf:�Ę���S!��Ι*/--�-_��s^�}�Va�k�Z�ׅ��{#�Y�z|A��kL�sL���y����^�h�q��5��YP�J�����J
_#~��щ�l-Em��r�JJ�~�b������+w���������5k ���p�?b*�҆��;�LA���Q�O�v��P;�x���FҜN�f����g�Y?:أ���ӻz��}7�～����XϿw�[��W^�w��=oii�����-��:�� ��^e-LeR9X��V��I�������e���F����3��������j�ye�f��e���k[d���_�5ͮ�;�s�N ����'cRA�����;��	򮟜uuQ�r���Y< ~~?f&����%K%�%/�WV����K��b��Ȝ�q�z�A,]P9��+�����o#ƞ��lX,UG\#̞ܓSpa=0�W�EK.��z%+�KIL"w�.`�Ĉ�ht0���c��ulσ���L���<������. <��3�=��c;��`~�5����f�+YE�����٪���LrԺR�Y�#A��eS8�>������VG�@�Ih$�]���ࡃA,z���b�-��P��Y:��0��mC�������
^�|��6�$�y'����p�
��Ӡ&�[}�Jq��� �F��-]���pǶ����-pV,p��;��ɳ��-�������e"k�(e��T^��#��%�@�z�Z�����D�	-j2�Ѝ\eۚ(9r�PG��U�@��4�����0�u	^�y�_���ZοoN[`˞ݵ�����ۗ_~e�(��ݠd�B�Yt�֦Ϭ �)q
��*)FS��f�8�gKg3�U��>�g�E��X�$����� FCV�O��e2�'�w8*�66F�
ԩR��G�|>��+3:H1�
�舘o��ls~_���G����_����9}2���8�X��ឮ��b����$Y3�le���&c(�����Ď��N	X�[�u����uw����"k[d'�)�:x����������z�������w���y�#�=��i����sGA���NA!����������L=�v0�(U�f misʾ��e�2.57�� ��;�;���.Q�C���}�.�Zc�-�gd6�i����1��9� w��#(.�n�7ky��������EgWg���p֜�Q��y�,�/�X�P�����mY9 �Bl	���\x�赩z�Ǭ�CF�vc�N�w��o/5�f�N�:A���X�]O��D��~M�k9��9k����w�z���I��$dY)�Ⱥ���}�BNq�1^��7�Im uM��fD�㘭�4�\����'a�Lx�:G1��NEOW�l3�|�t;a��i��k�!�!<#��LP�Bc�v]4t�:K
�L�sAѴ�,H�o����ކ�{n��Q��y�C�v�e�1
����E���d���he�N�y�d&��]M��a�p`��v�+�i��e:R�����Xr��ح��U=��������=���o����ԓ�=1>�������>��� ��`u���Q3�]z�^B5;����xKBR5���&c�ɱZt��85��� �����>�"�!ͩ�4~\��쳹����s:�r$��L(��yg�A�}ZG�ϕ6?!������^�t�ɜ<�Ay�,_��;UO���C�G�kD�%;���(��K\�h��(	mQ�����ѩ�͂�:>���XRSs�;vݓy:���t���3g-��Ï�ܽs��1Ԥ�$���$;3'(��*k�>���&��Ήb�"���)U�(�B/�ik��ձ�]-U/�0Ȇ{í�m@���	K}���~����R�Z�f
ǌ;�j�S�ֳ��-�6�=���V5�h����ch:_3��p�a+����:;;o|��9s����-p-p٪�,�\A~A?�d
!��5b{��S����˭%Ur�N�iw��vH&N�d�N�76��_���ֺ����O�j�=s�O>��L��W�a���⢒`�Aaq!#hd�\�&������Lb2����tl϶>o����L7��f�c�x�~:���H�c�:����붍����΃��u�#B�D����G��)YN#~�߹����g�ohph��=�K����[�[�~^�SE�a�"��%����tr!g Ho��v�o�~͈Y�ܮ�p�rh�%�֬a��"��ǎ��t��%���?]�ɿ���7��dz��,�ĦMeG��8��/�9۷
�^�_�0� pA��@�WЏt:�DG��� ��KVk��3�����˄U�X�֌���]����#�s���&:�i~���\؀��9||��E��y�Y*`�A^s=��5ж;��~{��T��j_��)?v����;1��8M�^R3�`ނ�dg��ea�	��P�A��T�][�뀂|� ��S���G�,���Ǧ�43�x:�|I��}�K_|�~�Ï"b�������}���7�Z�rE��ͿgnZ "2��z��b/8�丘*�+�rZt�g���,j��L�e,��x�*�����>g��a-nj����t�R�F�Z9_����@"u�)�c��m��7c�Ξ�����:����~W�h���5<�OO�Z���%#�`��g"k�77]T���K=��޲y<6��	t�0�F�y��8�t��Y��.i��8��  ���k��d��tD�ad�"����B���OM
������������'#��kh�HtuSc�?��{�����^}��[�����9U���I`|�mS��D�\LA�_3/X�dY���r��������X���&� km^��:���I�v��* >#c��	[�LT���U{>�f'��w'S������x�;�g����p{�8�?���y�O�����������	��㽜 ǁt&�~F8���&�/o��+�U��������<�5���YX;F��Xz0ɩ��|'�3e.k�h^v,�Y�+-&���B<��������k��X�WOI����/~��������5�l1�u&A�����Hm[k�u�_ݲ����G��x���/���"�w�������~������\~��`ݺ�`�f�hc�<�e�7�����jR�"���2�}ۘΔ4S񣨛S�U.6�d�:��^��Gw5y�(���<�֠����lm�7O�Ɲ�N��/�>T�ҎO�����=�8��J�$D0�ʂ��[rr����=�< ��q��M�I�_:箓܃�ΆTPR00޼�K�,���[�-P[]�pKsˮ����S3PGg��FS�	k�\�ɐvf	����	k:ZU��[�A�MI�#��T�:�����4�2�{:��u��T~�Уcc)��Mg��YX\�b��%���L�y��������[���뿾���ޞ��e������2Ƹ�&匌�\��u���w�]�=�Į�|�_�x��Wm�zݺ�S1����Z�С�e�e���r����R����K���!�����S�8�s
98������\j.�LZ#�N������R�|4r���F�z�#�IF��0��;��Ϣ���B��S�]��vVz�nX�-�����uo\ĭ� �$���:�4�vT�2Q��vW�~ Ei��t��31����eɒ����K�O��{�r����<���zz�.'u<s�Q�(w��59� ����4}�뒡�t��g���:��~0*�"C�#�Wl9���n��U��mN ��C��"ѡ��� E���.F>�����҉��>�/�|��������*�LD&��KJ����׊Elwt0�ڻ�G����Q��5"tD(f�$�cC#�8�"���z�kԷ47_��/n����]wݶk֭o;	;�Mγ �뮺�lW�ڒ��8匠Lҙ�S8A�)v��y�|��6%68�tTw�I��� W�e�Z�Evl��)��e�Ԁr�^�ᴛ9Lᗕ�ɘFk��������~�y��.<u�ֱd�ai���:/d�K��;ܗ ?�C�22���8���z�ƫ��s����?~nZ`�����6�����Ŝ���:��O�ǥ��`���bz���+(`�5�'�ʶ�r/H	�u2�u,:8� "W�:�<Y��	@߶s�[��;ߞ��V>>9�=4<L�.��D jJIAyb���q,d�l�0�y:#3#)�^��̬�C9Y{����ܜ�Ʀ ��)��`lYTA�~]F@����
bT�QCF���hm��g_8�����[��{�]s;��ʓ5���\X�`ss���>�'����C�A*R_�ێ�3o���
Q�us�zs@}֓��IRԈ��S���u��V�S�Y�м���X���o�C��u�o��óύ�F�h:�"b�J-�*t8�z�B$'a��U�u����ci�� �r���(N�����ɴG_���ի^���s�[���8_��,ُaK�p}.N�B��*䬌�9Na/ �3kƋ�d��;n]	w��K`@���6�G��dI�A�AԠ������035� �����hV��h�<��0�v�_tdge����t�'23��� ��y�	����E���;a�\Q�)Nl*.c":='
鳓͑��:04��֑hQt rUkk�U[�m{ߣO>���_�¿�]�z���Χ���Uu��6uu�=�����ȱ�;��!ʀ�\㨇�=-�U ��R�D�
�1�&'i/7������L�Z������5�'��<����*pjt�ly��1��v9f�zF@gt��7��q8JERG��N`��dm�f��H�E�P�#�#b��"{�Ԟ�\��y�e�)��$1o׊+Α�������@}M��?�0������J���
FR1l��Pn�����VV���c(�o��5!�IN	u�sM�(���9�:���Яذ~/���9�� T��!��ΉRSR@J����7�Z"�4�JiX����6zYI���u����ّ����#;;��<�ޏ��_|��nx�M�����g�G;�}ll,�Ʒ��g�v��PwGw��$jޢ��0A��8/�i��g3ґ��ҍ3�������x�kdNOZJ8����ML08g��̴�M]���t�|�M-�HLz��l֗��=�q<*�K��d��0�׮��"}:�s@�/N���4��{�z)����f�3Z>�~�����%e����Whvgf����R��)�R��C�NR���G��q����ȭ�N�9r^�\�I��	ꃃ���'/�_v|O�ϰ�� t���֪�⢾���V�8���Xs���e%IR#G���`1�,q���al���[���2���IM�Id¨�sƦF���hoߍ��1
����ڵk{����#�S�}^��[��(����O>z�W��C��)�.֞4�<�a`�#�LR�D� y���HWھ��si��#�Q �Pj��"nK�kj����W���p���}���m��#ޜ��鸳7��N�X��gjdn�̣��<6I��E�����/�V�;Rd��.@��y�y�L�w�ϟ����M���.v��������3]wh%��k���'>��5��sVr׭���:�h�X'�M,�P�6�I�U���<r�����W�x���_]X_������T�VO�ᦦ��~�[��e��2�.�IB*_��1Lߚd�ե;c�x��X���:F���L�T̖�T+����������խ��W���Ճ��;����u뾼n�7_u��9�W���w�~�_��-[��i�t֞F1���΁,��JTM�5Ȼ"���nh�0';��7~ca��;}�s"�Y[��7���]���,���*�cA�X�6��.\��[z�Tܸ��C?Z���&��9�GC�����~��v||�N��ht��>WUY%��l����%������w�-p�[`Q]��7�����ԛ8�!5Y^��2�+ʋt�鸻��㶾��+�����X�����(C��d 2�AzNN^�fǎ]��膝�w���e˷>��s�J
��)*,<��a?���2!��n��ϟ=����۷����M����z�0�X�-h�\�u���ۈ�0�Ч�f�:��M�r c��b��4e�f'�����񡑥CѥM��~����}�/��W\����z�[|���~��|�����r������ӓ 4�����h兣���?��Np^@��Xr!�ۄ`�n�l�#�Y�.#v$��t����R���qQ�#�Z��%�ҥML��At}�v|&���L���ʖ�i�s/!C'F���f�?s��ݸ(@=ϱn�H�:}Qq�8�ii)P�+�aü��r�O�'�o��`-����)�]�3t��;��YI ����ϒ%.W�F��2ㅵt>c�[̘`��U⅖�1؜��*+G�����F��������컵 /�V,J�pi��ܜ���n�TTP�f�����#y� +Su3C���r��߳u[����������E`��S�Y"��b���mS�A��j�p�,�S�=~4��>u�g�7�� �;��F#��{���߷w�o�����V���뮽v���+FO�����b����Ư�[����V^n�7a��2��������o�D��<)L�����{�V�#
{�$���.c(��iq�i8�`���WR�'��m�w��$)�d�s��������It�"i}W��9)5��I_�>�׀��DH�
ql�+D�=��Q�.Y��/����[�[�(+-ٗ��ӆ�B�C�e\k����qq�=�"y����[S��F2pXG
�Wa�WN��s�y���~��^ڶc+j�o����t=��:-9�h&6[��3P�l�̵����{�3{f#�>�BGVz����'
��dd��%'MƆZ���*��Hyv4������`$?'Ƃ���A��c�v*�O�z��6�I]��6 �$'� �dɃ`'5MFIXX��g5C����ؒ���%-M�wmݶㅿ���µW^��+��=��o��h�����?���kV�'��YN��1==J=hpz�k��)j x�K��E�r��;C�)�^Y�gmf��ŻÈ��SU�\�b�dr��dH[��]i�3@'��	 �㿛2��y�n�
AX�y������Cxn�9�Rj�3�n0�E��竔�4�z_Џ}|�CdR��b��W@7_4��ss������N�y�����[���{zJݕ�(�(Y3�~���, �'��,a������@Jj\t��%�'�2<<��$��s�v���Gq8��}cKid 2o0��������|��b��+�X�t�����g]d�ڣ=鷧�b��)��
��'u����s{�|,#sp$�@-<��0��,,*Jʊ��rD��Q���4.�|s�6x��~)��&M�T{2��<����^R؃����%1j��BeoW�/=|���/���?��߼��k����xl���8�M�������o�s|O���������X	^�?��
q��-�|����Ս��sv����%Ql�U�*g����E�Jfq��DY��562��E���@:�P��La@\�2��TgdB�!.E���� glyi���!Ǣ?���Ld�Ld�<�z{{��@5���
(HK[VN�@mM�7ͫe6�߼�N��e������am���S���G!�2�� ����ҥ��]�	@w�2n�p-m��#G&1ru�V�82�~R�9��#^V_�h���m]=����W92<R
�Т޾����=+{��+��,��W��,T�&b9��`=dh��ӯ)���'����#�8�~�a��� �r��]h9(*F��((-,ʪ˃^DB�aH�B�s4� fT�-��O�f�/=R�m��<��MMJ��?��wi�"Ik�@F� zrC{S�۷����?����o����ի�\�~�'���Su��}��<�������{YsS�/PF8k�̐@[	iA��4�</#����
D�h7���+Eo:�_� ���*��wM&J"sQ����ֺ�͍�'�͎��m���h�wu
X_�m��aix������\��gSA��L"tu^\d�j�$���}*�mѹi�3u��?%a����~�	kH�o^�tɮ�Z)�F��q 7v��E'���q��0�f���_�t��)v�sE��+K�Һ&m����/�_�;��,��PSQF_���w���|�б&��D.t���E������L����Fzj�W�%�O��Ը�{R�槳i@=�ĺ����� �\"�����;u���F���1h�"�cXY��E�ę���!SI=������V9P��������<�����_|a�j>���l�j��S����C�<]�Tlނ���5��<�Ep��Cϻ�������JcϷ�������!����R_�K'��� �d��(��d�5�ݼ�3 �99�"�ʺ{xܡE�iS�M��r�Oz�.>k{�1�1�8k�����ś���?��ꌲaC9J��_�n�<�(X��5�Hql�#��!�.����p^��9���>���?�/_�^/�k��sk������4�k+W:fxMI���	wm>���k5D�ӄ��M�B�xXc��妳���V�,�q���i����?�Z�`>{�xg�Yۮ�'��u���C���w"���͚F
D; �'�8�tA�C]o��Ƒ��pOw�9%%A>�S���p^A0�h=�{/�#��a�a��2ES<gf��N���DRT)�Am�?(?Kt;�BA�=*�vt����v�K/���~�����g������ʩ��3�,~���~���݅ŭ���w�_W������a������߼iϾ���将0�0�fD��eL��RؙѬ	�XK��P�ӼX �����B��9~�(��Jh#O���ik�p�7��1�R�wѹ���~�o�g�0��?�=�4��-3`�7�K�;S�$�i��:l�����t|:�s8@���D��	f)����<(ȉ&���LV{�T�5������Z ��6D胸s�-b�87G�^���qD8�t�uݟ:����,[�[�T��P.Z�	��vAD��[��AyY�����ʋ��Ⱦ7��/H��Õ���it���C�SV����u�Ԯ`2?;��"Z�ȽQM�t��"*e�Ζ�3&iQ{��>�A߂�y�����f0:b��`�c�C�\ꉩ`x�C��
sSSK�M�n�z���c7l���5k^�~�/��}���9t��;�s�R��=ڏ�{WA~{ai�o<p����ֽ�:鱅��Ӿ��'�������?�ߤ�v�������(c���8�S��z�����G��΃���K*@���L��R*���!��i�-suv��-�.���k*�i8"�]�|�r��U.m�,�P &w)�=�q�}���i�g {�����<8p`�h����-�==3]J%E�ߺn�O�;���o�- `BNr�{��p���M�*[�@���s���~؀�ǛO��)�}�5����L�O
�Oj��,��iϬ*=��.F����,�lw��H��iXX�@v�[d"�1��b 籡� 6	����dD5�л�B�>T\��W�k����x��!L)Q�s�<�I���!^��!i��i��+-M�������\<�7����|��G����ߏ�����]v`բ��M?���_�W�Ww�����`�5��9Y�9�Սm�o y�}�{���o�t���/�t^Y������z�� �������6ms�U;3�5�'�-�Vc&�iԭ����H'.	���C�t��-���J��ą��5�p[.R0��]���h�� �3´���f�W���V�U`�<mP���:8�x���1g#++����s�>0�Ɍg�>�1U���͋-��z]���8�@GLz�\���ά5"fp�O[=��F���r"� �ZyO����������|�??#=�^\�tZU�����I$���z8"�g�"�
�؅�0��x.�9y���� �o:�l�PT�:laeyP���E�>��NKC�Ϟvܱ���Vb;�v����N���`
&�Y�e469`L{0<;T�Y�eЎ�~߁������?}���_sͣW_�����ǟ����o���hp��D�|6����yUy9yU9�-�5m��Ғ�����^�`�#��?T^Tx����'W"�|�Oy��{z{o#3�<��wUcSp6�dkѲv-�����~l{�y�j?�b��C�&(�l�3Qb�D�L�;1���LLK=Z���'�=ƄC���;V�Oc�ԛ��)���9$��|_1Ji�C����k.Vq��ec��J�}"K�(����#�Ͽ�~��>:?�ſ�R�@]I��W��`���qP��(�άѸ���xV0�K�X#r��AȢ���ר;1��)��'c���f^�ɏ�e4��1c|�������ɒ��D���T���D���	ԴǨ��4��Ӑx�HL�pnz���Ӆ(�[��s�C����"���`4�G=vNH\B����T66X� 8�"���$�/���S�3dǳ�@��щʡ����cGo|�嗷~��>�����n���}�k_�5��tOk-�@��x��c�o8m(�ĸ�h$R���W���u��c��E��G�y�k���m]^��g�̉u2۴��%���|�O>��ݷ�z��4\+*�����(��9���E0���t�5��Ү��lK��S�'*�)h�T���3�
HmFo{M�p�K�1�ψ��h�6�8nq�|gk%`�9�X���6K��|���޼�i:j��o(�:�<��xi�zWWW��5�ǆыb3�F*p�B�i
BM_��꫾s2����[�[�g[ <�qՅ xgG�W�
W@7�=lhO����=כ.:\��>>3sRX}R]�?�ƻ��:�ׇ�952�964�/�7��\;�߷~vt���O��i.�X�� ��d>`�f��'��2]�4�T�py!��8(B�>��:�+�"ؾs ����mo��Q��j!�s('�V<{�i��J�Α%X�e�}
Y�(��C�$Hx�mhjn��܋/��g���!����#~Q膙��$�m�8�t~2V|�C��3���}	�#�����?x�m���Ƿ������VWU�^�h�Yw�L�ˏ�/E~�-w�]�� Da}R��`�N�DF��H��X�b�Ė0�<mʛE���B�64{�Ѳ��Y{f������U�F��2UMDh�@gN��Z�w����e���=�,ZK7�{8�nN�9L��!��N2����Ōh;Gr���ͅ�"���}kkk���<榦&96�9��y�t��7|�e˽�논��c� d@����?��)�$Ҳ�*�T���@���)D�ͨi�
�[d�!�c�k����['HR��	.z@���W_�՞�c�	�p���܉�����+�{z�0Z>���T� ��I �4�ol?0��6D�HuO��ў i�2�����^�R;{�+;~�7�Q��&��̸x����_:��Ң�!	�$����X�'Sƃ鑉<�����gS�B�-�����!�����58A�� ڇ�;�ѐ�MGԶ��XӪ�����:�/}���ϛ��yu5;�-j8)�S��ZZ�r>��?�x{G������W"�A cJ��f�x�J�+6!�qrS�**�12�����5Q���>�'`m�������q�d�J8u.����)`���e�}�o�|�BF�!��>?����`�qU9��;���մUN���y��`)��T*��=�`�?� %��/�,0�K
K���9����=�Aa	t*ˠW��;���W/[�uN�d��z���u��"��$����8��0ʬ�6r�&oǥ��z�.:��Cʴ�n����`�I�\��_���e��e����Gc��ߝ,�Ԍ��^��n���d�@���@���p�,�=��5��	���dF"�d�u�=AAy�}���¼��� �B:�{8��䕂�5�Y�0R��Y�(H��PN�Ɠj1�ce?�PF��H�3%?�7(8�p���5��	L���Ϣ�m��	�^g��� A6!�__^�)sEGWǊ�G�����������ϟ�ե��ϯ�f���Ea߿�˿���p���z�;�k�/��Q�"1����y�S���&	���@tk}��L�m��S]/&f(��O ��� 0����Z�X���"�q�6ev�d����I4�U��͉Kn|i�Yoi~������Y�@�� �)\a�=��T:%oyLt��"���Q7OE&����O�IY���~p�W����u��7{o�S]]����h���f�>1`�R�ʫaz��Q,��+�j�8���)�~i�����sz`���Åc��Ý�"m��������k�ʛ!�0���_]$_��4�c�AVaA��>�C�e�h{���PЏ�Y�l���t��N�&ӞiztL�HX�8�D	77[I]J��`���z�x��K��D��.e���SZc�z���i ��&U�E���������]����z�k#�RSU�T[Vv�d�H$���bx�����c��5�y�[�\̚pRJ��4�*�Oޏ�[	�3Re�Z��rs��E7����#G�ֻ�0�]T�Y��=I|�>8nt����X��n��:�c�i��n���y��6i;!�]~?����"U��a��]��Q�s�=K�ٿ�����;l��{yإۥ����	r0�uf6::;H��.^���o���?���k:N���o��������`w�K��Z[d�p덄��K��$(D]�����a�Zv�G�?��J)�����<ﻧ���ND�F�z�w�i�`�l42P552� �D���5z��H��f��ЅH��2�ɺҠ�l<h�}#v��q�dj_F�*),��+O���F;Sьd��ּxw�xt���D�r��q`�:@M�a˖�;>��$�Ǟӟ@3������x�!9�����f��]o:t���9ه0�cǿ|��%�iŲ�N0962��isE�]]��(-�z߂��h=���_��!CP�B^G`fo4����I�2+�Pbj� ��wF�	y��� _WW+#q{��f]��q��;L���� ?F�2┥GX	���=j��fm��Hy�&g�#uq��9+p?6Z� ��~��8�1�B�
��p��8��8mȌK��2����cΡT��=�o���o�������Wu�u�[�[�[@DA��ǈ�>��S���c�[Υݏ[[$����k�v���{��+DgD"�9>��3���S��S
)�vޟ��+km����r�`{�-c}�K���ڔ�HNR��HkSYn_�۠\�lD��
S]�E5�,̽�4�F%����E`�D��%1��g$���~yi��I$������]r�PLGiUS�Q���Z�4<��c`	�e�y֪����� �۱�J�I+�K�V`4��Ntv������Ntutd�{�����ȟ�a������!n� ?�`͈�#Iԣ�K$.�J�p~>���j}ٴ� �Py�(]0�+�R���::�Q(����t��y��y�ŵ����1Q���f������2 ovq���jc��5��.�=aJ��T̙�ϐz�. �x+�{/���ؙ^<38�p4J��N{��6>�ܻ�}���s߽֕�{�)\�~So��� d��6��8��c����OL��v.Z�윬I��Z��YL)6��������^c�̪�y�����h_�HG�����[��;�O4�Ej��0�Ǩ �#�r ��S�T`!���z ���g����8� �:��Ј���@��)��>'��L����W�]MO�`���¬��2͇�{=s�XFօ;)�Q�F7���=Ñ��[!j��;�+��2���L��j益$+ӿ�}����)��Oٿ���[���H
��k����$@12/E���F��@�(�� /1��ǂ4�^8�)?��/-@&8F�}(0�o�ir�NS�)�/�ӑX�@��@�GI՟��T��@Zu|��P݌�fM��ʮ�`��y���㎧��?.U/ut��a��9�7�(���%ǽrժ������M��>�:�n�Voo��g*�i�r����z���ys��9�։�$ә#��u^J���kShk�Z�/�y@�E:����J�	s��<��^�|�@[ۺ����F�;�a&����I����6��L�#����
���tc��F�?cH�"�S� �!D�<�R8s�;b�J���D�ᚸ��5��}F�����],�� ��e��W�Z�|�-2죯��{$ �M��x'@	���|8)�)�HQI�{-x$r1J�g�r=�W٣�~y8m���޽{Y�V�39	�B<mS���\�?[�X��4:z��fMa QDK�m�_:��f�7����t��K�+�I����O�l�'��y<�n�<I-]���QƠ�M�����4��;�+�楳�b�w�~L�q���th�>��̛7OT������k�Wan�g���u�7�8�EǓ~���Z�^�t����A5pO]
G�a��6�^7�QT"Tp�`gk�/��}y@?�_�$ޓY_ݏ�x�9��hOO�P{�ځ��7���^��E������!m��l,�y� ���`0=Y��=�!�_�����f2�UH�L�p.6�A2��\v��L�M"x�f(��R��3��QH���wp"ٙenIIq�Zl�r�
q(���7.�g�yP��3n?����D� {�В�E fmhb�zD�r�⸘ X�s���ǍҦ�����&�[Slmd�(#pJ��9��#w��虓ӌ�B�Ho�8�@&�����k?�l�ۉ�t�z�T�Wn�s���Z(6e6Cd0���u�Ŭ�@�5���H�#s��$
T���
�}ߓ���HY";{`ɒş�`~���[�uZ ��µ_@ �z���,��P��"�p
�>Z���j׿<�t���b��#�������'
���S���tuUF��.��u�������%�ѱ�q�� �e@�??/7(�)*�󃎼�`'Gg��e�{ WR_�  �T<k/I��'c�d���� �7͑���r�#J��1��	�tْ����+�B��*yԟ��{8g�-Is"�B�D�<�Q�%�d9���O��*�������cuZ=Z^� ^��0�ð�!2��6�u�>S��@G���8�h�����#�e�N?�h�����$���� 3|!Y-�@�NUӀO����!�>٫��d�my,�kM]�'�@m�����2f<�ΰ0[���W85*�����O������[�[�gZ Nu�<���l��d�H<v���h=ޯ�T&E�
R��i�h�=��"���6����#��h�ر�hkۊ�֎k"�Wew���F�F�&��<�/ө /�ـ2�!/쩶�-�Ғ�q3H_K� �lnvm3����6���͆�LM���t鲥��?�~(�e�͍*� 
f/4ҾLc��d�# sF˒��kt�z��`�jB�� Xz����:�\7��B��"�̈�3�)FCW��I�|cc�K�Ca7�)'��ِ�%�:&f1H�"4�hQ�8	 ���k��nN�����|&�)�n�Ջ���^�o��/��]]\�]0��l����}t[*OA��[���;m�V��v啕AuM5	�?�lÆ��T��TZ�����.:�OL��8�Y:jQ���A�kk���^9K��`(������e�C	�Y<�ii\R�Nz@�΢����c]=��m��6����qKW{Ǣ������)H/��5Z��h������9��:��/"�)s�{��Y"�C*�h��D����� PK ����=�`@���e}zl��q�٣D@=qf�T��`�L/3ʧ��LFì3��*�\œu�nF��`�ә�����c*1J�b,=��.?^5���D����E��Ǡ5z���ǬJ �%Q������Þ�?�������<�.�-��V;��D-1IM�:I86����)o�m�xM4 T�G�n��6���L���
�6�A���(���QB(*+
*+�ظa݇o��
�Q�����������X5�� ��i�c(%2�(r \%BDV���t�9�	��UT �YTk.(�2)�x
�r$3-ݧ���{&?#��l����DO���;�ꛏ�l�?��l�jJ���������Nlm�����F�t�w��#팒ڥl*�n�R�V7ƶ��냷���¤f�5����4e7k����<�Ǔ
 b�ɚ�	��dd���{S$��y겳g���ŜB���1Yȥ�,�5���>d*@�m�Q�z'ӛ�od�kkZbn:/ �p#�ِ^~���Vt�$�O���;�nf�6[ٿM�=�ꁻ���Q&2,vq�h�;6�[�+�~ն9��t�0����K��A,�^�n��~�g\��L��~_�� ��D�O�yTt��\��l���.�&iL�� o@	��xH�T�V��L.N� ַ�ʾ��>���c\�'��,Z�zՎ+����Y�쿒�2�	:nB��\�~c���$�蓧�xڊ&B% D��F�N'@������}�{�
�к����H���$�1��2���M��o>Ǜ��Md� O�廉�r��q<��/���Hl�c-ip���9���Lbv!�?�;"v�ú��1�y1�u :	(���dO?>��n�mf��~�p��@���bMגƿ�q/�d�9OG�Ѵ(��4�@O��a�}��*y$�1���l@�cqc�/�Z�s�_���q��M����[�b�@ot,	��f6c����l	L�V��H�S=^�˞���o�Y:�\�+p0jπ>�HX_:�U�3���5���_ g�tjz_*�ӠΎiF�RTM@��F~*.�h�:F�)�~�MY�e
Z���a*5m�;OB2�)p!�u"�H<�6NIZe�� 3҄���0�y�J����Y7r���-`�Ys̒���sD�~kE�|�����}`���G6�i�X�Q����2�N�V#���>w΅|'��a���[����!�N'۳�/:�^y���`]Rj��y���O�nVb�w`&����,Ɉv��Gݺ�ULN���w��O���r����.*�F���Xs�;|�H����+ZV3��8�\\]�k����I2tX�D)�jvf�����I���n���5/ �9��&���$Ǔ ��Zvuc=	NdYꙥ'u�I�w�<��Q�X�q�������8�s"���-����v=ݽ �a�,<G��8X�}�<����	NB����k"�ʺ>f�'�V��w`�<[7����� `��k��ۻ����>��ؐN��E=�f�m�|�������-������(q������,K��5F��+�䭾�9+�H�8��gԍ�^��Pbp)x�\٘���+��d����� �&���'������[��k{��Y�?�[�Ҵ�@d���b.�.���ȩ����ʝ�u���2��%�4=k�N��� �/�5��BYs����������y��p[k����ӵ�S��uD~Oa��Ө�Α����r�B���8�V9{�U����i���0�T�d�Q�b-� h�"5�I�3zg?;�aH�cʛ�����r�Bd�{	zL�kߵ:=��jJI��Օ<&�eG.1�'i�r�<��e���N�0���E��j����ϤC���B.��:�p��O ��\��P��w�m����g`�Y\h�9|/�li��Ѹ��tVG�����񲦖�����~Q3����x˟��Ϋ�Z��yx�s������XC�s�?-*�k��"p�Id��Ѻ���k�^���Ć5 w ���<vE����I���m�W>�!���z
��� i�t a�G
$sj�.ݮQ(�yx�L��q-�vײF �W??���7K�vo_�Lwc�7EM���d_��qH�c<��+�N8F�z2O�,s���8�uj�iN뱟��vr��J� ѐw�{k�2a��R�4��%z����dE�^�?9��] 5�`ύ�F�:A�هD˝���p+��LE�y)qÜI���<��% :>��� ��v��T~o�=��ao�Ѹd�;�L��<h�����֭����w-�O��::�������8�$�I ��������2����zD��Ҡ�9�ѵ�e�Lde��2�Pb�
�I�<������F}�I G����h�Ȇ�N�T�VkK����-�.���:�d5:'0���t�/_�<x�/��H�r���#K�i�xO��:8�iu��Ep��k����J�ֵn�� !�׼U�֍�1��XP;]����N;���4��`��-f��'DX�c�Fg���Hx�N�՛��Q�t���L{؊� z�*��<k:��M1��K��)���u��,��g��ϋ��������"z��0z�D9qZ�u��v��G���|?��e�%[���>g��doo�}������5$�)��%GY=\P�u�)p�k�V�L ;X�ˤ�%y��-�6ș��i@��Lg{Aa�IX�>�������=���k'��RG'�PN��3��LG����*�o���fYg��y��d�ҥ�=��#�7��@<�x�D��+5q *�s�&��e���L%)�{@R�p�V/�z�,��<q�H�����֤�C�����1��X��L�#�q���B���,�*$�q�Yֶ����udA�Cz��X~��9|���y�I @,�l�^g$.�n�����Z��x�[�A�n'�?�I��9]��K������&��<2�?_X�`�?U��y\�h��\4�g��9T�K��5��AJ���L�S�Ra2�,����
qk�(v���R��ŵK|�~��Y�����[��t�%ܙ�,��q�(e�/�D��͌`��m�:O��	ȿ��:O������|�ȹLY3'P�`�\go�c ��)h�笭;"&�q��N���J�R�Α�\
Y��nw�g�'<kG<�eޙF��O
�&8cl���U;]��0�\ߗ�X���?��D]��N>2�	�B#`��3Z�I�����t]��p7�7��F�_/v|Wf ���8�X�m$;���dM�3�S��f-.܇��m��p���HAa�LMMu�b9�����P-���z���H!����0p�u�k�d�z����v�+yں� {]�4e��T&���̌����O�V>B?k��m�}���W��^SSӕ��}����u������	��H��c =;�|	Dr"IszP�;�i��B1P]c�t����E�a�(<P��q�Z}����g���r�*Q="Z��	x�NP�c��u|*�i�&��}�J@�:�NT�����	c�=;P��(8	2������t I��9�]<^n�'ֶF�x��3���dm�vq�s�y�S�I���:�,��<��D:���F@π.���T�Cd����Y`���8��i�K�h���V~W+A���.���|�<�������������������#�����oD@�J���s��,�1u� �@< 0���M6$J��32{���:�:�@$�f�b��Ik/.-~�T���S��y�������?���lOO６���[[�ޅT�*��+Y'���1�7��	`P�yeEUp���u�u��g�=��e��݋�l:�	��Z"~�40��T5���{�-'4�k��)j����'�u�b�u����m��֋)J��9'��BNH*>�Ji��٧m��F��e/�F�v�����Y��`M�DDgp|�	�xM'��e$b��@�N����*���u:+��u��)p6x��}�9�4?�f���a���B@���9��3Av{uuu�`�B��<�������@kG�5��+'���Ӈ��RJ�<e<ch%�8�;��Z�ʱEg���ɕ�t���3��ܜce��=�by�b�9�müZ���y?�������%��}��������yYOwO9�ռ�����dɒ%��ܘ�f=9�y昻N�!h\i��	�'s�9�)_a]��7۵�6��n���9%i�vN�e�C\uڂ�iu�3�"���	tTE�6Y�.� ��>��D�UE�x(�+�D�t:�N���)8��A=��XM�ƲZ�:���E(F���:KL��i��ʓz�?,;��HJJK��JM>��g>�������� �gb�j:�}�[�8�&;+s�������[���@��HΏ|��QJ�I�pP�g���&`9&d-�;6�E@���5�31�7c�8U�W/Y9�{@?kͱm���c?�V��i����W<t�}=9�.�% �	|��p;�K����b���ƭ,�Q�h�z5S���EC�G��8O�qe6����h~�՘�.g�m\v0�ܔ$�T���i�IuͱWM����պ�E��a.T�S!�~�t�ɵƲ�<��ݛcb%�q8�'��q�w���ùA��r Sc�!HM������L�ώ�����,c]q,�R�5��z���L��b��S��OB�!�/�(��5��P]up��~�p�.=�rES󱫣�T��3�Z�����s4`�����mm���kt<?G�:a�+	�Y9�������ɩ���Zl�n����ྙ�o�-�����Z�����N��mL3
�a�&�A!��'�K��s�U�4�Ir���"�'Q-.����|��n���Nl��x��3#]?�K��]{��&���mg��#W9���p���%�g8�L���(t,u�U��Zi�ϳ�`^�e�N���:[�rs�U��΅�,����Qc�Ǒ�N���d�!����8��c���������AB�e�=p� �������YPSW���noЩ|��-�-p�-��?����O�2n%CÃ��4�5tZ&G�̶�p]X��Fz30��TG��s��%bM�S68MP�l����w�_���Zl�o��O-{���lkmMko�D2��' �ҧ���x	�K@�7��4����*⢠|b�G��:<�8f U\R\�D�L�m����f^�����
����~��#��E����$4��؅���5��h^�X���2C 7@f�k�[�a�	Sd���,g�<����T�ua\�K���΍dtJ�(�Q�S1��9�y�r6�,Hk�n�+�s�$�!m.8N�X�H����ߧ��6���6����U'5>q�����.84��_���z�0Jh�f�5ةEZw3�&n��m�
� ;�.L�ө�Gf�r2(�n�z�{���~��������ߛ�����qOO���B�9�<UUUV2c��4��֙��!��H��m�'}� �
��#��%@�DSp"�U���N�;���;�V\7��%����mY���~�pL#�eU\�����Ѝ3e��"�/i{f���.ǧ��ۅ���c�X����H.J����tXӶt�I�2z����q6������6sڔ�`փ���CW!Y͈XD�F@(��^Y]l۾���[n9���>M��y\0���>�ӧ~����b�&�\3e�d0�o"��$ݮk�1��J��X�D8Eh͑5�ʖ`r���Ɋ��㺊��䦓����4�\��S�������&�6�G����J�zK�(�B��j�m��Pb=��Q���D"��f��{��8~ԥ�	F<qxr�U�GIs���Q��	b�3%?���'=w�jMaf:��yRK*�e����7uF�=L�K+��KEh\�� �����0�u;[�^�+����|
���Z�������}�x�=��5��5�@i�����Fg��X&�1E���m|������h
u��WUU��DwO��>�>�/?|���?x��#�n�D�$�h��8�H�9������n{���Y7�Vqn:��t�@�57/�k��ں�M�cR�c�9���~�sw>��S=�4��<���~�|��M`& 22$x�D�� ���S�XU���D*#+Ҳ*��<Q|��ۆ��܎'�E�Q0A�.b0�K�Qx�4C���c��	�$ʩL�"��ˬR�ե��"�SIU� (�Ko;��2^��H<f�����}�$�����a;�Q�hWf )Ťy�ql)A�2����C��l�KW����\;Sl�pe������&���P��Y��G�U;7�X�7�N98���;#�?z��?��*����8BT�ԅ�+��m�-|�8N��5Z�ꄵ*�KL¬!��xNWc�j� 0��%8��ř�~������O��'��8 tq@�u�b�:�tFy���2ܜs;�KR@�Gw�i�$ ���E�T��I.�-�����sB�*�ik���p�4�����+�M��R��?�ؓH��F����Z����7S�TO�)h��Y`���=]�.7����x�	�<�W���g�w!���.��,��Z��,�caFB$f]T�����덟�@l�~ǃ���d%ˍc_��2!�_J	�̅�'4���@D�D�3���cm��ޯ\২?|o���������H��Q	Zf%��VT7��K��&Ʌ�)	�Z��,-�u��{��5��K6���r�Ơ�P}�<U�9ś�S4�\��3�w>���]R^�hACCPQY)l��~���
	�@M]v�x�{Nw9Ay����j2��N�������r�%+FI��0�Ļ����@$���8�$��M�T$j�j&��sy�OM+������d*���Z���lq�����U�Ď�d5� �C[� ��@(�I�^��9I����t��R�o���\1
�uoc���gD�3�mR�,{˜t~�aLgRb��������7�<?3�� h�h��sp�e���9��[�R���C-�������ʦfGESHf
��,2hR��(j��P�IW�9W�Lm�e�<I�|ƦDr�x��,�Xc�6���WS�������Z�<���6�����l��5��J֏���G�/zd.:{%�Ǵ�K�w����Q�nLyӼB7JP�Y4�Hg����ƈ�5�y3�wPJ�
)�5$����g�J��(7is*j�?�Q�E�V��6��'i�v�ݖ���򌉯�mJ���B9ZҌ즑��Z�`�j��{��Zfi~��mq'(�إ�Oz���hB���vdLm���L��w�D�xm���q�
^9�	u����\�q��y>���{\Rh�d>������zEoOO0��G���j��A�����m�r���d9�,��9?jR
kq�@d��ee�O]�����5��ӵ�y|߁�~���?���[ZZL��b�x����N*���n/��z�"G��l�"�-�"������E�L�k=��pm�Ѻ��I��wf�?!��Y��4���Udc��V�O�s����B�f/��8�@�[��dڊ�7>��	�b���zP$�ʹ�4��\+7����҄8:�w6j�a�4>.�#�=��7�ڇ.i��s�cd)�j�d��/)8���;�-����(�SU^TUW�CX�����f�U��E�o�����w����C�����/�sZ�n�������[�2�i`�ȕ�[�ފn%S�C���5o�3)&���������z����c�s�޶�����Ƿ}����-��W�I>��*�n֖F �T.��M4&8�-I�n�0UPִ6�U��E�FP����x����IZ����c|s[k˰1���E��1�ZKo+��C@�CkG7�}�Z�V�9.�_)�h^H%x^�i��ZX3����(4#�.��_~� ŕB�dɵ�DZ��� �Y�Ii�7`�>Ǧb;6#hNW������oQ����n�kgg���<t:3#H��#g+���]E���A�����}�����zp��_��ŋ�ז��r�9>E��y\�xuǁ��>�؟vut��tuKGK���Qn�ɥ>g�j`ckO�O$k�*�u5M�}��?�s�9�y9�>�X[SCY�Ӿy@?mӝ�7"*�������?��}��uс����-Q"�f�H0��8�k�*Vr����y��0O�sl=slrI93����I$j�P2�ǜ��I���*�1$z	4���p6���$��dP	� x.��|�Ȅ	o���J謰R/b����>7�b4t�lk2^����x�H�yz��G=KSel/Sr�3����?Ϝ�ö�L�㦦��d8I��NO�uژ�a���6s��L }�H�K�;"����sU��=�Fx&��o ��b���Rs��;p�@���?|�'�W[�c��e�4��ܞ��Ӽ.Lj�*z��G>��ܼ��v8�X7y����o�f�3K���#~b<y<F�c��# �lJҪ��YP_�ŵK�j4u�7�i�s��}��}���_�n��[�_/`����KK˴O��Ih�̍�M0K�s�4q�f��u]2�S�u�bXhcϷw*'���$�	R
�<�$S�Bl#�<��6g�������l}�҃��`c��S��3����y�v�HS�i-d"��He[��m�
?�Ύ���&�r�ֳ�HP���5sxMEE���9�e��Oq<<F��I�Jo?3.�g�\2�z�LA
>���0�ho�ϙ�T���x13����t[���QG�a��s���utt����*�pYeů������U�W~Cw.[�0r.�E�Y��^���:�����+�D6s�u�p���^��y�Cd<+Cj���K�N�-�u����9�K%Ņ�/^����k[�ׂg��O<�T�?�_>~�����MLd�%����9sA�b&S�3�ձ���F��~�7H�'܅U�����XÙ¤0��D��bg>i5r�K�3]= $(�L�U��8�H] ]  ����Y3�a�@��e)n�'�8�I���|m� Mg��#�1��<�qq(�^z�܆����'��T�d
P��5Ev2��$�1J�xڠ`��s:Hyl���/�_�q��P��f!����0�o���{�l��;���nO��� ����� �9(ā--m��r��߳c�k������D}}�-j8�b�B�������)Z��6���SOm�}��rݳ#�� �:B�x��ʌ�����������jr}�iĺÌj:����|Έ�����U+0����<��>���w����/��W>���~_AQQ�2�ƦX��cc��"F�F����~r"��N��ѷSRc4I���(���Ho3�60�@q�(k�(euc;�$�t�����1�5F�2j�%��f�G=rz�:�T�6���G:��g�vK��q�Z�6�h���W��e%�q���#S���|:6��H;��U��.B%bb�����$��{2J�C���ߏ����c�s*��
0!��U�XoG{[__���X��9&�6��ߝN���?�C_]I�Mw�SS��	���ή�c�//,*�����ѻz���_�_�p�7/Y�i�|��7oo�_`�ǟ}yË/������]ȌEpCޕ��j���=w�.����:bdҤ�8��k3��=��yA~^P\\�y�Ϟ������Y�����f��[Z^�Z[[��H�5S�P�0
$ �!O��D'$J%�K���l�N9[�\������]ݜ *� $X�۫x:N��M�'(�^vmg̦�fD8���'�8$�aҦ&#\g��b�l;�L ]�tj��O��oZ�T����I�P���9���c-�����X758�(ZCN�C����k+����!�aJq�Ɯ��C0�t9�	9=��߬�@>��x�3F��:G:��=ɍJ�S8��T�|'��~�a� 8 �aiIdKM_wOaka�eE�%�8t�U;wn�����E�\�fm�Y8=�.�.
<�i��ǟ|��M�;�Q�@Ã��)���+�c������5��(�h]`�0��;�!Z��Y�����d�Ϋ��ʆe�ψ��9zZ����71��+��2}���Xĩ�F�VF�)�R�eTHb��� �	�v��Ⱥ�4���m�́;�Ϡx
�c�cN�z�A(ZO�pB|mXɤ�>��n1�Dp$zA�7�:u5nֿ�A��CS�`��5=������G@��]��Qܜ���}�MMt��5����%!5t����n����hZ��5�L�k+Z��΁��$��u�Gܸ1��o�㓡-�o�G~�.����9{L	�Io>#~���9�?�=���4��$)��33��q�F �Y��H��O�)b6��Dn{^ޱ�Goܱs�e�e�>���۲t��//Z�`��U�������[��[`��c5>��g��Z������:�Z���YN�(m�L���\�����u���$�j���d��d%�K�iPJ;gb=ຜ�`��9�g//[��3��=��)K���|�?wOoo��^�aCQSK�0+%Җe\�Z@�S�U<G�!��Ӓ�*g��1"n`CL`3��g��z2@��kS�M真#@��I����0�)p�4Դ��ԅpG%:�X�vivRpi+9���8��-'|�La��ah�d$��Ia���&�53r�̕F�$�2"�C��쬀2�v���3�g���R�<n�$��x�ԑW��<[�hK����Sσ0�j�S^��Ƕ� �G���R�8N��w��w��3ڦ�$�sj�9����v���6�1�YkӓJzڅ_(y�
��\(�!�> <&�ERz��kolYp,�Ђ��w�SPRt�c��̖�����K�]�jU�<e���.(���\����|�W����A�ublX/� �Ņ4`Y�WW�u�'ץw�>r�����o*q����`ұ��`*c> =;/;Z[[��|�)�I�Y�N���q��O==oϞ}_C��F�΃��D�$hh��'��*����BT�2�qT�[SȌ���F�nuj>���L�1�Q��]��hU����-�n�yɈUW��64ʟ�m���լ	xB�c!�u�ڗ���9兢�<�D�l��O��)z<�3U���)�i,����G��ʼ�ia4,Y'k�N��R��w::�=YSJ<.����q䪍F�u@�x���475a_�K���Ngj�����{���[2����>��U�^� il;+]��@�7��p��j�t�$�7Y�2���PH~(mL�������^[W��˖m�lŊ�q�^���]�xe۾���~�o�
�������m�p���,����� �]m�	w☽�d[�Ld���d�nN�@�+���4���
�-�����\��V���){��LY��k�����ވ�iZW�UFs&#:/o�ih.]̔QZ*�`��*
G�3}D@Q ��S��8P��*�~��N]3���~�&ѕ��T��53=͡% ��E��ɺ�[@[j��$��.�M f
��֙�f���hS��hJ-�Mc�3@���c��-/u,|�LBr���9Ԅ��Ni_�qˌcMH��B3Q�Ōy��t(� !@޿�g�|sGdF��k��BIٌ��e*��6k��A3T���9��s�A�O� ��;�~g59W��*1��?��[�Ӊ����C��hd0����v�v,m:ָ�����w���/_��O���?�`~�ޥx�����n�^زg�#�?�O���N:ȫc�jY��*\W5�� ���<�k����L����Du�	�h��v3h(�E�
!�E%�G�/]�Wg������9w�Бkv���~(�I:|xtD"?.��I���dR����-��f��]"n��@6q�'�k����,MwآB�q<y]-��_�uh�k�.ނ���<G@u�q�w���P�2Έ��1���O�u�-����!�J&��G�읏���sL��)��Ro�ߒ
gi�� ��&�
��'��d��Ɲ�i/F��3��8fKp,lY�w�wM��H�!Z'�P�b�!4EoS�����\h�ڀ87i��Y��؎�	�޺%�ѻ���4���D�y�Ǳ�����PDLyN����?2)8�U�w�ZUT\��P������G/^�@}ݼ�K��.��9ti�C�^�qx�SO?��������3� ̱�r�
�0Y�C�f)N�9�2��9�-�ś������#��\�~def#͞�"@�-�C`P��;��u��Y|��L[�4��A �^z���'�nb�7	��t�y����QO���&_#��'��Xj\ �m�Lq�=-�j!���-`��p��\m��D��IB�M�q���R�Ƃ'O��J�p�6'����{��.	z\V��(�<~�|�.��s���k����C�l^~9ܩg��τo�(�8X6,�����2�mE祤�D��nݺU����l�@~�~��\D��N�~�+�@�n\z\9��1{�S�.J�,
��)��n�Cx�aP�D�ʕ-ȷ�st����@����������?��~����?�r������v�-�Ԧ�^|��ط�����"`�#�85��!t8xq=�����q
�iǵ���-vm⑙�d�DFd��������AQy��/�t�5�����8����?��v�]���/�]$:xo4:��iQ99"\�5����x�Kp4�M�"�v�lΚ��ٽ"��DU$j�����e;��NJ��e�I��r�������4���� &inG�S�5r��Q�yUK'�hY@�� ��Ԛ��!��{����H���	��K��������:������̱���r��%EA-j����FG@濙Ex�W��A�W������y��$��V /��@ssK��ܪ)tqDTW���c��au��L~Q����5:�]��g o��<�uy�%��H��k6,�u�������#55U��.Y�u��\�l���́���En�o=��v���ɦc�6tw���|@�Y�!:��SMr����Z�Q��s�6�����vw]1! 7'Z��p�S�����*�ʂ�҂��K����g��>�~6�z
�lni����O��w�;��yz.�1c�O`�)e@�A� �3*�p0S��pwl~|"�'�*��|��T.�r�5�6�+R���)�b�!�.r�'5��'#PfH�6-�&p[��5g��rظ%�u FDO�dM�CV�&M�q�;[_��sR�J�F��8=��YŁ p�R ?�΅��˥�"w���-3b�ls��H'j˖-q8f��l�
�p�:g�F��vL���-YqN���0�o���xe}aքQ6�)*:�����������2
le�[�QH�)�t\W�dl��m �Oa��c�v¾޾"8����6>z��%%����+_������޸���O�;���oz�,��ћ��SϿ���7�i{k��h_/��Q�ba@A ��`�� ����u�AV�Ws��S�n�p;�ۓÓ��	5�,���<��s�����7�]��ٲ���ϖeOb�;w�۲e맻{zߍ�sY�9=�7@a��$IpSH�y�p�5�T�LL��z�ʰZ:��Y��k�[��L�A�"M�����}�
�2
TR��N�a/q	T��ۅail>)�	
�e*�+<O��VW���vk�ˑ^'1%L����1�<�Wz���4G�3`����:�l~aa��t�Tq%	� �6�)�"���DA;]�؞|���رc�	/=����Kɸ	����W��O����b��q�ݻ�ĝ)��(��ߢ$��|"D�z{�9Ε���Y��c��+_"�n�a�F��(��ʄ`�����S�#�-r�C/)z|?
��<�L0[n
Xl/-+�U?�7,zb^uu��ŋL��$�~����ٳ�����^���v���m�����H�c���S���:�u���;�]7zmʿܨf��5��w�\�9�7�k|OF���@�;?(.+�\wIPV^����6��M��������ϖe�~w��1��W����o%ә��ĸ�1�JE� M���/�Mx�F��%�#	�Ew��a�ah��񤺽��5t!��L��U���5i�%�٧�֭�k�o{�6�uN��J:��eL��,v�d�F�-`'����J�ʂ2��0�ܢ~�1��R��|��Uԛ腳�Ͽ�zT ���s��HS]z��>s�������{����Le�+p������:�O�}f*JKQb�К(Yk���X��:�f<������H$�#�]����Sp���左���I����8Q(w�\{�~w[�X��GR�$�(���� �kaAagii��ob��E?\���i�r��?OK�%��?���7���o���o��l�T2�o��]v�o���W���B������6-t��V�N�y�����Х��b����AiEI����~�=������y@?����޶}�B(y���@��Q��ɰ�@-���Q���<��-f�"4f6�%�[X��� �����l'O8�!e�����L9��!��Z=�љՓ�����/�s�a{��]�.���;A���yGj��&7-u.��߁�8 {��=YR�W����[�j�H��m�%�Ď��@PekX-\��Y|?#�'�1
f�O�$�MX���$+!����Xm���s����Q������`�2�oll"\��1s�����i𻺲A����7�bw���n�9V��q�KdsYNш��C��.�l(��GqX$"a�;	����ag���H�`��������#����т{�\�Ώ{=�̥���4>���۾cׇ�;�p���N���2~SX�(l%�i�#�5�kI�������jZb�$	�2��gs�9����ڧ�C.�gЋ1L���h�a邿��[�tq����U��������W�,ߺu�?��&o�Ƙ>���h�֖�6N�v��S���Ty��Έ]fnSY7��p
^��B��)܆�r�U�z{<B��,Ol�ǥ_�ʹ˴����5)k��PE�z�S����
c-[���q�X���S)	((���\ۙհ��2�m�!Qa�)!�A�v�-�Y���7�����g�`��$=���E��:>Qu�	r�J]�t��$���x��<޳�3���v����,�z��-Ph+��1Z4���F�v�����7��E<s�tq��Yj>q��4��"vI⋞�>�YW��	�p�g#rσ�f��U�F���,���E��/[��gF��!<����(_~�����֚N�q���\�uO3�X���M�U�ru���	���i�����.�%�N6#t^�v%�3��Y+^a��On��\�f�Ywl=����dv�}��e[�m�\_��#��Q�$��id��> @�Ȝ�iN#%8l�HT�'�KF��V4���c�Z�h�H��O���P�+��Y��窥�e���I���M]���^!m9���8	p'�h���6%;����Z�W��<W;0��w%Ü?��A�#'���Ό�]|�`�R���c�[��t�Zx�<F�<~�Ow��x�N~/�p:]Y$�,$��؇�6��3���z����+|	Ȓ��h^�\����e�o+mH������uw�{۞�����0�h��ۚ-�W|�s�x��U���"a�3���K�@������a�4r ��hii顺����ͫ������x�U^��d��ϴ��#��^��F8��_Gg�>I�QLK�ZC�'��″�\$�5;>��Ĥ���rJkpc�F� E=]u�ymq����
4Վ�yaA����m���oz��s�3z@?V�g �W����Toj�>;q�i�htP � �jS�<]��I��d�6X���`'�*����P2�������m?�^�H*p���`ɨ���������q�S�UK��!�}���\�n�.�hN\��,�����8��ɸZ���`�	T#�^�Fnn�8+n�	���(���x�2�9#���nѻ}���8o}cK�$B��<���|H#�;u��F���u*�)��^ 2Y{[{p���!S�欻��e��	�1�}�ND(�'�_!�I��I����Y"�2&�w��g�9
a@�!�W�WǍu'^�>GG�c�@2p�$�C�I��Dv��ɲ�Ҧ���=�UU��iX��e��e~��9Z�.�9�ڑ�kϞ�[�n��#G����ٓ��Gj��5�k'��x��-#v"���dy�2D�$�fՑ��R����k%gN���T!��wPZR��а���{���seo���һv�^�c���ȯ�I�Z�I!#�l��I���* �O$)I�kJ��G����t���ү��Ie'��0�y�s�梏���V�%�9�#R����x���WB@#��!@�y\R6p9tb�_�v3� �i��	�V����N��bF���D�٥����mៜ�����>�Ke[�펀ލ)j`�Jf�� KFl�NiGt	�����g�}��l��{�}������*�7�v5q�� ����fT�.�lId��G��]���B� >~S��;��gk,oN�}x���%�2⸹(��+����qJ8ɏ~ U	�f����x����Y\Rr��/̫�{�����W_�y.M��������Ʒ����DQ� 7W���RUE���̓���51��HRhn]����Nd���3�I���\3a���ѕ˗��5W\����������e?��37A��F����X�d��O�����p�1}m�n���0Ep�گE�V'�EԄQ,"�e��Q]\wF�N�Ep��DmMS��p��B ���=��%k��P�<QZWM�Z��7�XsP�}�*�\Q^��q��_`��3` _QY�>ӈ&�e;_7����	 <��ѺJ�B��9|�1��K�<�c�&u~q�ql^l�Ҕ��긞�a�Np�1��[XHD���oʌ��q����,ț��ه�Y���#�l\h�D/�<ns�̎v^XVE�8��<��!�B��q�!�Im�+E�x����7�0���#Uv�wV�6�ܰ7χ!���g����u�5^�+w�xS�Y�L��/ l;p���m���Ç~����5 �FHS�=Yc�c1�ғwf.m�T��f�]�a07���.�6�Z�uH��8�e�f�fKKgaa�TMM��.۰�K��u�f�g�}�֝;v|ndllA|i[���)���,��	��� �΍�.�@Z�Ֆ
W[T�N�`5�I�'(#4��i[S������{�5L��
�E���g��g.*;$�y��7���<g4lu}~�Ԕ��`�7�������~t�ݙ��3*6�t��d�Ir�;�������x�s�3���#��=;wɢa�d4x��
2^��|oqq1�
\]-K<v�tɌ�g_xN~/S�S������1������Te�q������'*|J�%������68[�4z���-d'�N�C�9�W����P�u��wH�)�?@��۵cL��iyq�������B9��JcIi�����{�������y����jͽoڵ�z��w:t��M�#}�CCY7��3k6���a<3'k3_	�V~3�8ҩ�϶Ƅ�O=���hm���:�"�ulʅ���$�ܫ�ʾy������W]w��=�����ɧ�yCWW�g;::��d8N&�� ZԔq���SҽAi�b���If e�	�V�BcF�ª�r��%��{�����DgM��+-�Bߧ�h�˙�Ք�&�L,eQ���g,.#X�������MÜ���a�9V��{y\�yA�]�=ѓx��\M������E�?|70ퟓ��>��Z;��)�,I�߷/8���x�4��^2$���! �x@��P!�N0gt��K/��޷G�cݟi;����)�@�
ԗ��n\�x�Kg����x����0Sʦ�3+H�3'24
���"s_Gzs@l˲�N�(��V!�-��$/�0��<&s��촗}�<���$��v9I�^<JK�6������V�W쭭��IeE�Ko�u��u���:v>w��+[�ڳ�� ����"�}I� O�P:G�ζ���<�Dv��,�7!׫:�v-��bk��pfo:�/�� �݇�AL��x���3�q^� �K ]�����_�q�o�u��d����CC��=�����zttlq+��9�V96%����M�@��?'�qAF*���(�#:eS�HNT,���z�_e�kz���E�ZK�:����ə���y��	O-o�����_���I��0ծ�m��q��YF���߼`+ X
+���q�%m�������KK[��X�<.Ɨ�K��9>�-R�ÊM�6�kd�Z�k��y��ኽ�"g�\��TN�6&��T��`ѢE�K/n
���ER�֟j���V�C%��L�����h��ɕ`���_�����,5rl�M��ƹ�EEI<�7���(��7�7n^3=
��� am��s��1�o!����(�<����9�xq��EL%��	�-��ID�}�Ȇ����"N�,���Q�� ��A�6a<--���M`Ԏ����R�8�����q!�97/��R��w�-�Ȃ�d�}Ś�*Z�o��|i���v��0wwuv��>G�?��:�G\#\�A��.ܓx��h��/o|�x�(�z�z2����	��f�,�%� �G�0p����4�9k����K�Z�h�o���{��/�{@?��G��^z�7�56އ��J��b�Y�hS�X#2驖�q^$-��X-%��:84(�c�7JzݝČ�,� �0�c�����,��{xBb�ƶ�\/2xB��f3/�H�*��x2L�I��uh��
���bq����d�:ntSY#���ӯ7�@��p|f[~�lȑ2�2�c��ҝ�����9|W�?��f�Yu�(�c�G��"��?�I��x"���Ɩ���NS�d�#u��$���J2 �Gs$��ϥ�H�/]�Ldd�٪{�t; �� G��3��KDx\T�L�X3���2�]P9W�jn���4L튠i���.��h��ԼE�vN��yb��;FBb�@"y:rj�#�qD�����Ӊp|9.a��]:$K�;�L{�y����IHy6�W��\UQ�x����Դ�lX�� �m�Z`ב��CG/9v��:�ΞeCP�e���0 �I�_�L��ua�H�X�S�[�~"���#ALrR��4��Da(��q�\��r�+���Lz�)�Z�[eE��V,��;�r���id�g���<�Ӛ;v������a��A0.���Z���	B���J��x�K���H����O&#���S��L1�QmY�4�0[�H��i#���m�n)l*��5�⍩QM+��4g��)fK�&HzP�㵃�O�6n,�Y(�$���ˋ� �;/8u�YQͶ��k�����#�d�x��&;�ԭ�.�:�q�(�/~iC��6a;����t#Gq�C��������Q����)�q8�+$j�j'���z�����L{:tdxs�򪫠�4��nM��v�u�=Ih���<�������Š�:�76b�^T��
'��E/z����vP�cG����J�ӈZ;l_��(Z��z��;9��8p�mj<�`ҫ�Bx$/��r�|��HAj20�L���a��O.��wg�5M�~8��F؊��p]M�U������4�TU�nX�J��Z�hKG�Ѧ�z �����Ύ�#���(����X9�$�8鹎왬-8?9 R�-�X��sP֢.)��:��t��TKY<W��	�R�+Ѭ�s�z� ���8ۼ��X@�i��Z����{��w�W�ʕ�o�m��{�e<�ē7���g�]]W`�J��&gk��"� ��8eO</��;{��[I�2��R���H�8 �2����)M�n\����XU,!^SrNE�ea�r�՘���%ݮ�� ���-^�*�a,���E�<�_���J���2M�U��3�6Pg]Jj�n+�=�Z�-)a<�(}h�r�S��T�T6�`Ir��9�k�oRZ� ujsv��P�^�C�ع�l������4��yu�X���w(�]�c ӕ�%W�3�ed+��	t ��o��������NOK@YfCgW��"��� �3#��:UE9R�u~�q7e���1�F-|���_X6Ǣ+;�w�]<5#*�Q�3�_�E��=�,o��>g:���M>m��s��h��#~��O��C�<�x����n�l�����G�.�'��9����~dfƲr�� �ъ����˞����Z[]ՅL���n9?�����$-���-� ��mjlz_Wg�F6-J���R�������*�h�)�zy0�������:vN���fqf����i&�����)��$�C��HI�N<�:��dbm6;&�Q8���˗-��w��'����f�OӼ?��C~������;{z{kG�:��8S�<�H<!��K����K��bL��:h��,���5�c򃌜(�A/QOp�q�� wF��}2��Җ�jL�[
S ��R����2|ܩ�9�S�XV�c�H�Ǧ��f>[[�-��Z�%P	���8x{��Ô{��>u|n#���+��T� �!�,��bA~�D�ܿ9.V;��1c�[� �s���;�"�F2�S~N�p ����I�=-5�r&Ś���P:.|j7�,3>1@P�+r���e�	��а��_�������f��g7��4tt�����y3����Z���踎[���HI��r������\9��5�� �4�4�9ik��4�T/�{� �3ҍȥ��ۯ����5�'w"�TO�X[WsX��	�k�G�-H+�E����k������Ж���3�D���n��Y�B�Y��~3�y�<��98n}iG���}e��O"E�������.8ͥ�����Lio�9|��ʶ���C��J�^7F"��(ERHk%'f���ڸR��f7u)r�;O����>�9��u���s	�t��^������:���ѩ'G�|z	&������|��_��`.��?�N��g}��������7�E�@~�N0��IB8�M�xTLD{����mg�J�/��$�ț^"����0O�t�}�����Y|?�����Z �{�g�gk I���er2�@�¥��ES.N'J�C���Ead]�u�7��P­O$v�jvC�iE6ԥ�ܱ/���ܞ6���V@%�%�����uu��N9�L;gze�:�ФH�"����'є��1͘\��1�����Ĩ7j,)�ذ*���((��:��3gΜ^����Z����7F���q{���������{V}����.]n�2n56���n��}&rܝ��p��(]�\y1��{��;tgu�-�T�mn)��n o4-)��K�0��v8���++^y�Yg���_���}��v�=��-��b�6�������ޓ���~�p���ڣ�
�w4�M�ݻ(BU?��px�ǋ/�J�<	U�y�re���8�O�^w&�tB��=t_��#j&�wO� �2�ɛQ�����z�g#���[���k�q����:u�S���iVg�V9mܺfvk�ޮ!:[ղ�����/^|㜮�K.�v�1G���w��+��}��7n\�I�jO^ѳe�;w�.����@%�Ft��QdF_�!t�yr۫�����ع��<�5�)��idM�P�щ�k��I� y�ɥ��à��u:af��8T9�]s��z�!o��׼����NB�O|�=������������-�W�)tuw�-�H��j�!\l�@��=s���2����R��L� ʊ�J�[�%�iޓW	��dyvy�"Q�|1ǎV����+�͗/�s��P� 1H,!^�����e�|!���Jo��W����i*��<U�	�9,o#�+V7��y]��0�]wBf�XEA]���yd?�b#s���q���1Ε�4��Ӌr�(�q|�g^]y����杯{�Ѫ����>ͼ �7���XQ�p<��0jW����K�Y-X�ؑG���}�EW����=��ky��G��_��bE�Α��F�����`�atx�c�n��;�:^a�j�$�El�<Nh^�������,��ƘE
���<����f��<�ۣ��a�pc��7�
ɕ�uUr��t@٬�Z�G���aٟ�Z�O��B�״n���E�ظ�u�HF� VDY��b,[�\[۸�~�~���G�̞s˼�ݷ,�7o�ڔze�q��������}=�'64��l�ڲy���Q���z�n_%�ŚY�X������Z�.{�.y�%�����:q��D��+��bX�� ��߸E�=����i�����OD,��A�і�C�F4TC��"���j���Ⱥ*g~�a�W��^������1	���F6l�4�c��[�}�wީ�څxn�/��"�b%z��!p�`�n�L��U���bÉ��z_�������G�����O���d�[��g�*E;Y�.>nQ<�9J�a�7ij]��P�?F�4���)��Fȴ�P!�g���r�7��W[�e���r���T��/�Q�ї�.ki��b-{�x.�m^�+�ޢ|���y�ku[q��X�·��ܪE����5�ə񣔉�J]���C����Zu�y�V��6.oO�z�֏��b�ރ������v�j���^�S^r?���p{��nظ�;z_.r?yb|�P낐�8�&	�[XO����8�}��M �->�5�M4�d�p������D{��@�q=YD���k����Q�r-i�F2�k1�F#1��{�M�sD,�oƆæ-��2W{/�$4'z2Q3R
��{��L���#�\�BM}�-m-c�)ϭW���Y��K����s�~ޜ���̚�/nPQ�ᕋ��������֭�R���m{�\y�mܲ����k4ri�ι��C��*h���3���v�]{}�=����wU���}������P
3�<���������81�C��?qf\ڔ�R0F���Z�+g=�z�an�Pe��P]L��9��E?'2�+_����W���S|+?�H�?�����o.^�d�CW��#Q�5�N�o"t��f;7�2Yzgx@CkYM%��ݵJ����uO��� �d� )r��~VYQ7��& ��87S�Q�86R���<�{Vv�����L�E\�Pc�5.�x�c��]��k�����6W�l���a��9<o<�c#Q��ݧ	u̓'/�9C=�*L�ހ�WX��5�!;�3Z���xBrD9"R���*���l�\}򓟴�����Y�m��{�g��Ezmʵѣ��l��+W���x�ǖ/��O�!���[�nذq�=���"uW��hЊ�Q�&�n�����F�봖����쭪^w]{4^2<���,B����}�7�,1��Ȟ�WF����:����:^���KC�Ǌ��v��#�b�(Q���4�P�s�s��T(�Gf� J~�6����h�Aj���^�y���Z���Ͻ�5���������_�>]��*��HW��U,��Z,�gΜ1���9������ɸ[<�k�\?�v�>�M[��Gg����948�����<�cv����ܹ�8�S������f�5��V��PR:N��٫�� q'���as�"��Y��V�,m�yt�d�-���Z����x�Z}������N����ʤ8���x���N��M�(�y�����Z�bſ}�a��3���A|�����S �g��o������C�w�a���'�p��ƛ�R�M��D&��{KO��i�J�CuO�_מkt26M����R��!Cۘ�"�^��̰4Ͱ��B�E}�z�mȊ튶@����J�F6�B,s�}z��]#6� �0� |�3��<�j�� 	��1�&\>�!�.Du����Q��.e5ȳ�=-��c�"�m�VþK��{�c]��7o�l-&]�G���g��9Ї���ڿq͵խ��j�j��m��ަ��c+b'����kad��˞
�CV�|�	ǯ����M������裏.QU�K���R�q��U��:%Wi��q��o��yq��ֹv�X���c�9�H��1��&,x^¢��D͆]�F�A�~%@�$���ͻ1���)�HCH>�� � ���M�|�vNv}y���AL[��	������0��^�vn|�VN���gW�u�=�k4pr� @Tu��ݏ�uT�����QՆ������P{[�v��+]�M�����@[K󠮽1]��Lj��k=�R�@63ys4��Y�i!.3��f�hmOU��t��&�&�\�����'&[�GF:����u��׿���]�w���u�ttj_��^թVɶI��g�\��â;����Wu�\K밢K=�]8��u�[�/�d͆����!������u's'u�� ��I��:�4��tyϣ1L$=�Sc���2���.[��׮��g�rJ�w�����|+�|��}�s��G5o�%6ͼ��f�ۻӪ��Y�M�R�Җ���sb$g��ҽ�щe�~�@M�:�r����
Û�����,7�#�#�n+�Ԃ������K��OŔ�t�6oN��@�s�|Sm�,_�fQ�X|�A��Dh�6�B�<���mh��]�Σ�v	Y�X�Î�gȡB���+o��2X�9���1�(d��Ǡ!O��ܢW�CҜz�<�������Z�W#ON8�&��T样��]�B����GV�X��9�S"�z�a�����>��t����q׿�s_����_.�ꨝ}���Um/9wt�<�i�Cǣ��	�M��}�$H�+��2�ͱ�mG���͍8!M��;��=�����R�xaq}�ǵ�5����8u�-��xuś�S(/��"FR�K��uiZO�s�:W�"�I|KK��?n��S56\B�"r3��eʔV�c��9s�����@�$�d�)��P�^M��ń�G&t�O�u�Z;�"��j��#��Ă!%�/n��S&wOL�"��麦�뻛�k`�dS�K��I�]���&�o�'�hꄊ�L%<^�.��2�0
��4���j{�}~�4���j藏Go��!j7��O%Bk�>�~�qx={�u勍�ߏLl��>a�����/��(�li�@��"u����7�Y�fnY�|��^t���;��c������KB�@�n�cG~��W����-�^�y��QX���E5$b���D܊7a�f����ԭڂҹ�@H���yxUh}�T�H��Ǻ�:l�O3f5!<�q7 �2^w�,�7Dbbq�S��T�<	6�ܮ�:7�F/��-'Ţ��#��;�ڄY�gl����HS�����I�M��R�N���,��S���T�ǡj���E��U�Un�BEy���`�͹��m��Vm޲ٌ*w�L����1��������u,�M9�W�^���������U��8�Ik�������p�޺u��۶]���y�܏S]�"��f�����ϩ�C��y��a�qM��nr������v7�~ J�F,.�Fc�V�b/E�q���Jj�ä�&TK���O���h��k!��#-�now����`0�0�Ԭk��\;?_J����df�ہ��mϑA`�=U�^w1���R�>�<��U��|JZ�֫�S,E�206ƈ�˧���Z�;U�*�rc�0��p�H�X�v��kS*�a-TmQ���/�����9v&�Bd�t�љ�W�ň��牴o�r�O�N�������6���=�AW�?�+��o�g�Ju��hL�<s^�c��E��� sB��@�;�R#�Y��5�9G�1s��<�e����k�:��Þ��Z�o��HB�	Pj�n��7�r��>��w=�n��D���E!oj���Ϛ�$<[�+��X�Qi����\Z��Be�RԆ�չw����q"���.-Eł5��b#f1��l{�W��;�(�q�Rm�'E+������ym�1{��16�S�C(B���)�ⅇ�~��O��E��ո�l�5ǋ�6��>88�_�����ݫ�9���>�0����TK�,u*�}�����y]mK	C��%�P�~������6Cm-ʗ�U�٣�8��v��M�l��:���UDQ�����}��d�.ٱc�k�?_�~To�B�{�E������Vx^ד����Z:���G���j�H�yl������?օyӐ�:ߕ�]��ۮQ72��'&�=����7WD�k�C�.��9<�q���u����W1��.�Z����:30J���.e7��Yu�)H�j-��-�p��r�����'�yËw2��|\>�
�(P�d�z��`�Z_Ð�E������
k�z��3��S�������Qܛ���/5(��~��i���N�X�a�������vMؗhD{��/��J*�ÚaҠ�PO�`H�#?I��ʙC�;�Ɲ뤑n)2u��T��SE���̒A>��#�8�O~�): ~$�?�k��;�]�|𝏮{��[�lY��:��W���H�QZ�s�� yI��N=�� ��,]��*y�Q��Fd��Ԫ]��x�-mZ�x�l��yRd���F[�eA`�{��U�.��Ó5O��Pu���KPO����"/��U)�,�m��a�����i���B5;6�(K��7�Ѝw��Hܼ�_�ya�Ĺs����p��S�<jP|�>`�`��5_��5��o�GqK�]�5�oL "�Ѻ̯ɢB�K/�n�d��*j���b^��I��,�K���\��(Bl�h�T�����g���p쑇�W��g�r�G��77����k?x㦍�lڼ����c�OoU7��`�>2:�Eq����u�w�������*���S�y|g����CԐN�N��=�?#�"���li�@f�i-�77Չ4��JJq!�p/��G����9��0M�b�)q^J=O5OS4�-a'3�Kt�C�jp�2/s��\���q�C���d��X�Ɓ7�Z�A�f��۫f��x��͌x֊��#)�^�++�;����͸����N�%"R�z�Z_M�s�<�F�C��#�[�(�s����g� �lŅ.��>�w5��u��&��=Y������s��]R>گ�t����i��h�(� ֱ������PI��x��U��N��tĵ)_>[�K󺻷-^��ߎ<��9���v��=@�����E]��o���K�����X�}#�hQ�\si�E'�W1�֞�-e4�+�^~� Bʐ�"����DH�b�.�(<���E�[�h}�ņ`��}S�˿�)�f�E��($X�GH�����v/�,t�mɘ�V������Q� pΡ���S�Ef��V�7g^6�z>�-i<��5P&��Qc�
��Jp6g�,r᝵�;a	�xM�έ�H��
udK�#F���׭[W]u�U^�Ā��{�#C Bo2�p��w�'�;T���˗-��)k�ݹ����N\C.�黾��>�.����w���S�F����j״2C�4ћ tk��(���O5�"�RA߂�j���5�+�]��pu9~7Y���9!8AX�xgA.�96�У�1�;�X��x�䲉 ����gax�������L�>K�5��E�֨B��W��
A���Q�v�5F�BO�&����y�)*~��5�ms��pc��̃7�<b�x.{$�-��H'�����'#�f O@��X�1܋ǘ�s�5�_�y�A���cx�+��؊��\�wk��T��h�Y����S\�5�I��0��|�'(ּ�|��p��67��aBʀ��f�"EՉ��D{�x����a���իV]�a���I�e!~��;�������9���ƾL�/ch���䭱�Axxz��bF��
��HL{�66�YX�C鱹�z�75mGV�b� Z��BTq��.~,K[bF�w4�!�R@d�E)�1��o���Btz�.�}�7�_=joVx� �(��ͅ����q��C��Y��ƪ�Fo>�����Ƭs�����Qp�"#�0�Jhx�ni�<�dm"�����f2��}����ߵ���橪\פ6��d�����_�b�#��
�d����;�#��%(�q��%�X�b���/Xp׉G�W� �ǅ睍�y�_���]�{v��7�j����?jtd�KU϶�N���zT�]D�����Z`sF@����Q���oFmF��*�q�m�w�f�ҜT�b�62�0��7B�E�D�,�WIzG��4�V�Hޣ$wh�G؛(@���2.vcC�X�嚏U�8A�\�֜y�~J��ηx��������R9~��t��5�^��8�A��G�	���1Ἂ>@�+�=��I�HZ������y��c���u��?/�w1������i��y"�=�f5��
�p�o'W����'�	K���4�(���GNjL:�6C#��Rd��ϿL���z�9�<�i��?��$t!��d�g����D�/>t�a���Ǭ/�� �%c.�*F���B�{��}�'YҺ��)�"w�<$c��6j������L�x�4�
�^�c�f��r����8���O�*��yꮪ�Ƈ����n�rZ!�&�f���Գ����և�p���H��3�$��R�g!� g��,1Z���PySB�f��f�c�KxU�I�E8JN��.��B�K�"D���p��V�R�̙Oޫ�uth�w�ҕ�7�]峟�L��㏙:�ӎ��M�C����E��+-�/r�!�:����x��@��  ��IDATQ,��l�^��w�k��ݙR�:\X�fgo��J}�V�}u6@CFP�M�r�Y0��g�0
�c����>e��.������G-�����뿐��po�Q-�]��?�{�.�Pt�� ���V��2�"W�Ƥ>LM5Ε�b��WY[��W����E<$Fh�'�Ҏ�������W�1`�mX_��k0H3�;�<Tn�^30���)rn<'��0Fϩs �O�d ��uj$A#�
����('�愫�c��U�������I#t��u�vΥ���0\�g�:۟t�.��E�&L�����R�5�i��U������p��|��Ï��٧��s�����5d���Gߣ��}�q6Qg��Ǹ�7u7݄��͋Ԧ�c���:�<fm��^�\l��wi�/~���sr�4�Uq��p=s�P�c�0˕����2������=��0��9z�Q���m�C7յR���ڰ���8c!��ݸ��o>g��y�(�s����}���/-I�3�E�,�5�Y�U폍�f���m��)����n�Y�:6�F�K�^��~�F�ͻ�Q���4h�����+r�8҄���*���u?��לt�_�����K��}���:ޭܯ��9�����yI�@��;{�عc6��|���i�.!y�XB���״W�"���kC�sF��zT���bB��	����ǵ���c�p�Bw-�=��n��<���ȓ�{z�p��X�I�em�X:_"C\�A�A.���H�aX��pqԝ<9�]�F4~�8N��}�k�f�j���iO���8��s�����5�87��7��ec�Jr7���c�� �^S"do�� �Z�.��D�*�K�ecj�>k9��e��8�n�Kr��Q�[
�[��2������I�ӥM�[�}������%/}	�%ϋ���z衹����_,?�sV�>�Bn�54���D�� ��El�~]d�JU���-e�����جؔ�3l�rQ[4,�h�;��$�.J�"bKŻw���E#�=C�%jgܬ��w*��{	~�ڱ��YʀH�<_ϫ���Mɭj��q��=xD�h���yos�D��D�\�:��<��+�ˀ��Dq��*�ⵍ�lH(��Y�5���i����D���r���7%(�G��f��"�W����sW\a��-mͻ_r���v��_�1�/U�)C��8��ө���}�v�C���n�Awώ�nX��U[6o;Smp�ʐ뤳���hS�R#ϑ�e#+�_( ����hb�g|�FD�hq�H�Md<0��٥���w7�M|A\CaT��AY�y�h�{O�H��R�J�7����F������E�`cKh��X+��9�F�9���������7F	�w��pƋv,�}�}�a��֢ak.����
��L���xx��rq�X��A)$���g�:�(�+�eހ텼��7�����3�/"��o�fSMЉA;ڃ��A��Y�|9wRe
�W,���e��sء�^��#���yr{A�e�����/\��URJRU�Ͱ���PGB�C�m$x�%T��q�`��F�>9G��bsj�H��f���i&�I�^���F��Y�X�,��iV�M.�B_H��Q�av��<:��v�1��%��t^�g��&��#φ��\x!���z�blw��!?[X^�[l�!�S3Lʦ��&.����be{�{��W�������{ɵMU���Wc{��'�����^lԒ��x���o�>���U���oK[�/y�%}��^���d�ﳏq֋N$�~=�+������Va�����_$}��D��L�N�T�n�%�%^X��,}�ڛ��c�WlZ�6��d�ӌ�kU�"\+�"N믋p@P��=��X�a3��B�:�y����w�ޯ?�/9����Yګ�-=UjUx|�������Q0ZK=������GT*�L\���|�!o�����Ǘj��D �3YY[-r`Y��S�,D���j| ����F!�2{���za��^yoCy>^���aT�����m�������^�/��Ɵ�4$[)|��C��ra'ռyӿ�Պ����[]y�A]}�!>������Y�/XB���O���~u��֭[��3�6��[mJ}��m*^�� :�c5�1r��	��h�BU�<y��V�Z<̺�[6	*}لJТZ��@��K'[\&2���N�e��K�Sa�Xx����E�����X�战'��UWV�5�ì���!yE'�	�I���[p|�^���F�Kc8�����@�yٴY�����eCg�ɰ<p�G^�r��O����-�5�+���@�"�9��Dջ�A�Oj\zU�O�{����K�L���腫W��Z���}����mӳ��~�ߙ��gǲ���W�3��yT��`@�Ǭ���8�Uϗ���+�R�5�\M{@��H�	Ia����{���䱟4�R*�c���׼E��K���E�H�	k�B���wJ�0}�&�-w�o�@D��Wؗ3l�
i<;�͸�#���T��3.�m�u7��|rXC�<|O!�B˭)���� z�=�_�j[��o//��Y�{��X���}!��x��/�S|g1�4" �9��q�n��~��Mʍ�m����kO�f�;���Ύ���ꑇ�7oxի��{~�^����ӻ��o|�OU���'�����q�,
��P�N��[/��d�)dW!o<B�^N��[����h��"�Ell\��m�/U�^��Um�!��w�:��)O������c��n��w�X�o.�.��=���ҦTwc� gJ�峴X�<mJ�����a�/(k��'6+�zR8�.�Z[�e�P�jQ��W��^�"$Q��̵>��%�@���f�/�����I�f�+�kEoVT(�h*s���`�����#��a�[l��b��e/��������>��g�ޯCs��������[6-�:;�`�%=�{NPO�*]����yVX�THh�S,g�΄�b�Z��"P�1�~���f��&�~$�3�ƍDJ�%a��뫑0r#!j5�q;>���i˛�����pK�9:M�DĿ'%�H���Gx>RY�_��4�c��	��}�D��u`Q8�`�A=�o%&kǿ�3�a�c_;6�u��7b6�Ý�I�X*�{��x���{�%�e���(��̭�Ͱ�s�GK� �v^D%Kϼ��2������3����7��N�3w^��T���+����i'��2������
l�ַo|�7��0a�1�����0�F��X0�����G�]���ZЬڼ���B��̃ԉF��M^���k	�a=�A[�	t�6�aGo�`+B)*��4�on1��"%���y��>���J)���(���i�>�P�Cg��,�Xg�-�Ro�v'��FV���^F�Mò潸��f<V�t��#���8b9<n������&�ߦ���:�6����:�ŋ���|�2o���uW���Z����i�Zu�����F]-o?#k�>Q�'t��;\w��M�=�躗���<K�t��j:H5)]� �)*fc6m�'�%�y}�\�Ng���Wz���0 ��)��8e��]���%c�A7<�:>����k�^Wň��q[��wk��H�y�5��U)N���,��!@͟�7y�
�R �Ǜ�sN�	R��k�B�A�&BU��<�Q���27����)ѸڹԿd?>�K����l^D�LP��N�x�}�v� p����j�DY�ރnpf���N�"���ޛ.�aۿ t
[-��oQ�n�S�5�~
�S�.͐9�\�3g@��7h:�V���5���'��_P��<�ԛo��ͷ�u��4�/n������_Y�mY�ޖ�%�ӅY K���E�����7��(dsJ�Ō��־,����"Y�}bQ�
T���� �HU�Q�V�����w6��*�}}��<g�j�Nϭ�Θ���7�U�(^b^��$﹩uj5�t%�[V&9?��د����Kn��i˂̰��j�i��cǺ��IqLV"�P��Z�v���B��l<�U�����2LF���,v�(��wL>�;����0n����sʙ3���FN0����G�~�?v�u7�w����B����P�
�W�W]�͹CC+����8uG����O���ǲh����v ��q������?��]�ծ3
�D�f���-Q"+�k�)�,B��4ҴȖ{��Vu]�W��N5iVNb����+浖�w�UQn2U�wa�7z�A�ea͸��Rl���z�_�\͌^Σ�U��҇��/���m{r�:F���9��	��~�c������q�@�(΀9D,<��d�!��m��zR4�o����,��}��~քt���;f�0���9�-�7�cR{������+b}��Ν����zۯ�������;sGo�UAB�Q@(l�A��lba3]\V�VH2�Y��Y�"�r!G.,�լ=L�V�����E&��6_��)�P���E�a*��=��(�ALٲ}����#D"��12�Y��A9�5�CL�(ry[��7od����6!+��&\�!j�-�>_�]��X��$�y�jZk)>���{^-b�U*v��f�3�E5��,�n��P�c)y7�-���^}���{�#d�'���ҥK/�������������_v����v�wO߾�g��[�z���%d��g���;w�N3'�d#;]�a���6���5���S5��J���@��&����!w֌y�~�����ʢS�i��~�s��׌��������cNtы5��|{]Y��kI6���Q�z�jv??'W�ZY�_Q�k� �y��u8<T�6���y;`����iP3
H�&���<߿�P����S����3E+�"\�M%���Ǡ�H�S̾EO����LGۮ0�7�,Y��K�,��'�����k_G���з��v�p÷߹a�7���xҭ5D�����i3>��������7�S*�ḻ�� �z��^�Z�ϱ[xN��ro��փs���?��F�����x�ͭqo� E��.ϵC��Ѷe��b�H��m>�s�ː�B��{L��<Q���y�dZA�Jl��PX�Wl�6
�8f)X�=ۢ1�D����{{[x-���ꆐ?ƽS=�z0������65��݁2�T�Gn�1��5I��o�>���یp��U����6�ۯ~����֛�U�۳�����[�E��p���ϐ�d�ޓ6o�r��!�Ѱ��V���D�5K�7�~tmB斛�b;76=�٣HF?���1(T+�x�X��X��2k�D�I:�}�m��Fr~R>>,n;�#�q��y����������ɹ���B@RcN��+�|�}�uKh�7��U^+��5���TB�ƽ/�a�[�9�|Es�D�hg-��תs�37i�z��4�[f�dn�o-iM6<��-��ͳf��ڒ%�>�x���v���c�>�	��ǟXt�u׿��ǟ��m۶7�ر�ꕬ綞[��y�:�:�Ch���Db�xУZ�K)Px�3�
/!���J~�Ȋ�J����`|1c@����y�^zs6�*��R�-J�b��Vs��ؘ�0�n�DāsW%��g
�ltIK�R�����FW+�)��ri����G�r��B/6ǰ���90Nx<�QX�����ٔ��1A�{U A��pl��A%�n����)�׾���_���ުJ�4<<�Ϧ�i?<��S��O����0�糏�'�Ի���G�=|���sw���ixg���׷J�w���h�fvG��kt�n�X�y�I!��xN3au:9n#v�&��!3ͥX�	����m�1D���[K�ԏ��p�ҟ����OF�+��|<�m^�������9��\�f��5zɱ>��X��@-~7#$N��݋��hY�u��u˭^�[�`���~>��Z�����6oA��"�Ì�wx��Կ�D"	�C�!���{�'@�"�ŗ�r�N<���jҳ�r����&���g���u�_J4�<���S)����i���[Ř&p3��6��;�V�A�w�Dj��Bj>#�^/
c�X.��(�ɪ�Y ����U��5h�2O�c�6!*;GԪJ��t-���!1Hohh�,�Z�v _hl6�a�S��E'|�V�V�F�]-����n�.�j���"w�>
�,B@�Y���]�cG.�&�������u�y��~���.��(X�5�=�B���t��|���W|���r�UJ�d/��}=��-�>��;�˅���d�;�P�������u�s�޲�댁���u�;>>y����*��:4�u�@�Vo�v!K�<���� �#�����㒳��|���Ɣ�2ό�bD�܊�XZ���'��9�ܽ��nx�Pv��w�U�d����qh=��Z'�x���3���B9�n��o������ojuLڵ�h��= ����1]Њ�yJ��~7ϻ(��_�k���H�	=&�ko�A0����,�̲�K�t��/ݜk��x��m���n����}�ݯ�뮻����_���[�l��� ,Q�&�Z��f���.zi��k=���mC�	a\�\ж��R�#�o��b�KX/S�Ͽ�\#T<Ko�o���-ҵ0�>��J����I6�B��O��Y>�pL�bA�q`yq_�R��8� ����M�c����{*�X��D#�u:B���1����O��l:$�h�sB�EC���*�g�\M��8��9���Dc����{
"�}W���k��M�z��S�}?7�����v
�_���7�ڮ�}��m���Ti�dt.]@��(�6�k�n]D\k�C�&v��9�^�_S�e͔�9��D;B��5��DZ�:�(���j7��׺�A�%�;���B��5/�r�%����c!��7W�]#���m���hܜd�1�Е��0�m�i�.)��p���t7�	5J'ksأ��Y7�;0�O��Q��ufUP��M�U��ܞ����tͺa��y_X�t���:�$���A�yI�*~[��/]��{��e�7o��:l$H���3� �<��v��0�մ��y[{���A�@�y��&��n\���M%b����E:���)?�&��t&->���^����l�T=����41�٬sDdd��ʳMl��k�m4�[5�+�M���Q_���l����h�Ÿ`�*��X�x2��"
z�x�ܬ�L�o��bvGC^�y"{��O���Xx����s3qm�T��s��/�WNܵ�|������u�a��w�駟��U�W����[;sw8�8����
�7|���4�a������D��422�xl��J#*�T{���i9�P͈M0���S�3r*�[�P�֩�:�к2BGyQ��v������篹�c1��qƑ��-{Ώ��='����zȝ��>�hOo?�<��0��=���X������kܿ�V���,�n�xu={�s�,/n[��ΤXK���#g]ư�`��:��%7�uMCS�4��mF��m--���?/����}ک�Y��@�yG������>����:�[��H��T�f<���Tex�]�^�D��C��m�;��0�������Z�]�^@�luQ�h#�ԖAe:��|�D�d�s�����l]� "f!r.,HP���O@sa�)S4:�V1~���gct���
]��x���]�0�9�.��Z�HAI%����\�=$�9H�?�c!�0�c*Q�/�b  �ߣ��͘�@��a:%A
@��n�B�绁��B�e�~���_��aY߬6Y����[��o��_��X����O9�_���A���{?��,�]س��t��ר��y�+���V�V���1��$gk��R2o]3�Z7tM���[/@�=k��</�{�م�kEf����j,����J�G̏��ţ6�-�������5�j�ȩ��R���ztϽ�8�������,�-ܔ$14�d3E���FQx�Ma��0��D1µ�Ǥ�Q���9g�MʍE��GN]{�?���^>�+B���n]��}���{�|�l��p�e�UL�����1��.ċGiB"Ǭ]�̈�'��ІBd�PC��rCǃ�}�x f;�=��=���E��onx�z�	DDˏcY6S�cc�1��u���p���C�%��X�&�Q�L�/as�����ǋ�G���p;�:�3!Bc�>1,��q`��z7�?62��gb�z��[�wxD:�7�X6��ex) $��)���������/�w���ѸQ�{đG��$�g{�y������6ěpG�D�fKr���O��x����*uN,��emo��m\�u���75;��Mʫ���2΂��!|����6�7������+�i�����H�v�&OŹ���c΀ր{��u8u�Bx�I�$�U�",�oa���"��б�و�＞�G͘��ʙ�@Ժx���c��	v���1�}�U�32�z$[}���wU�vü�so_8oA�I�e���Y-�B��λf_v�'��c�=~����p��\���r��P��.>N!8+�y��/9e ����PQ� ~Y��`���l�S���|��q��䖾�nU8b�-��y(����S�0`���o�1�~��;��R�V/����1Bi-F�Z;I����e�8V��F~ŭ]���&ϛ<=�O�h��ú�{�G��xo9ϭ��l���V!:U2��g�`݈6X�z�$9�E{[��I?܊���c����CU3u�>���zS�����7����z��Y3����N\9��:��o���&y�34v��eOZ���Ô���n���q	J��ބ�S�"w3�aG�<���E$��&�ٸ.��m��b��1d% ��7^��e�ly.�L�{�~������C�-�X���xn��xo_�%g�Mр��(^�u����}�+����۬����z�<.�|��wk�u���_�;��3_t*�y�G<o��K/��{���ZlS�<	�Q�z�B�-�Z�٥!.Shr�1Ԥ|j�)d_[��`+�&Dn��h*C�Qoax��Ex��R�\6V�F�83���q������Zr���}0�-T����tf�GH�H�Uq���we9o��3��	!���7�_b�(�[搭�e�t�w+Qn����1O����'��Ot�8�us\?���Q g������ j����l�MQ�n��
�:;fY��Y�|�E ftδ>T��[�S]�~�WW)QA�p�O��&z���t�G���o��^{��^嘷4/Z{,�Ao��*W����[4v��HI�؁�����#�Jzx�ĝ�IԦ[��v�+�f9w�C��QU�W55�C%�Ժ�U�;q�\�M"On��vK����_5�k�� U��YSh@��+�>i�����!�FJ�^XH�'�y��{�2����%��j�e�9F45�Lvl���<��(��4�k�آ�����w̝�u��!ݵx���'�9�ͼ=</����Q_���O�mV��'բbC�-��@������iV�~�B�б�� Ţyd�ݖS	�G,Ū�)����=׬yY�{|�$	ze�[��h�֥��F�ZO�Ř=�n�F�=y��H}q�bfp�6�҆�{JZ�~���<e���Ԍ�KGQOD�i�@&ܢ�~�p�\�����",�	��Q6H��/ <��G^��!�ذ(^�3G9r��G�Bz֫�TuuwW[�n��qx�|p�l�b�B����qmn[42�{+W���\����i��W�_��D�'#p�qG�όw�r}��i���M����~�FE��\5:$aܥ�K��L��b���l��07����!�B���cD����tI�!�,җ��ƀVU�����\���9�n��Q��̹բ�%^˿s�%��]>:F�k��R�F}z��@�98jK�!ң�ڡ�����c��3�=k��f̜�X����S�_���9�?�������������3f1[[��M�X
�G)�2�fz���J���6)W�㧷nQ<����{�x��"|��vBo�R��Y.���޳��u��$E����4R-[rd�� @rא5�m��b4K�Ds�<�<�Rh��a��x�>�]�lx�q�ԣp�I��R�|��S�Ќ��E3A�aE�z��Y�r_d�f����s��f��N[���`�p���y_���3=ܮ���߰a}�̓a�QG�n��M���?���,_���SO=uݯ��/M~�����5��#p��C y���>�����Ｇ�p����_�s�+������Z161�\�v�v������6����S�����}=z_<-���X�{���y	��1�.���xw��n��V��}�:1C�1�=��b�ͧzm��w�M��rQ�X��^�Wn�:Iv� ����Y����?lmi�����^�/�����Wk{./��п��S.��N]mH�I8Ha��3�Ң	ϓ�b���a�:R(HA@\�\�\�ѧm+�~T��^�V�^{�<H[P���vR���aBZ.lS'p/��r��~�c��}�\u�c��<!3�����x�cDl���#��{�ǿ����q�V^o�:(�-;�Xó6�ǰ(�>�8᳙Ҟw�m���s�K�йy�����u�!k������{�ܷh�ªwǎJ�ߐ��Շ�3�8�/��>��?z{_`�����rm�{?�8�أ .�;t_�{M3���noi��ܬ5<S�K�ѯ�?D$�H{��щ��Z�jm�Ԧu�"��f	���L�ͧ"z�����a����O����E{�yc��B4ˣ!��Kѯe�v�kO�=k���׈���O��+c|��^��t��a��y�p�I����}@�]w�3��������Y␙�G�b�7����UkmeX���2�%^�D��]2�ɪoTw�&9E�
��H�zͽ%�rc�$�ƿ�`Xh��r:G*^M��v�F�;�8�zA����#J��16�
���/�K��#��z�=)�H7�f��(����u�]Q��g��!l�+��ء(�T�ʂ����q�4���rgS�&��L;6�q���x�(��x)EU����y�=�ܣtʴ�+�/��Ͻ�5o_s�1;�-x�x�	k��9������8��^7mlr�E�+=��f8�+��ڤ�ѥ��nmZ6M��=���U��l��69�ڃ����^mgS�)b��&͚5o�R*��3U{WGg�E���kV]�iD��m��w��lО�#����5����'�iin��&�;�Ȭ7yί���	Є~�׮ִ�ө�O�ֳ@@�6Ȭ�J�^��J�u�j���+ك�!�]S�,U����}��'�N=�"7�ɦ���.d��+&�X�𦴦�O�.�dʗ�b�zrT��e6� >.��:�6�P�����n�~����q��̴7��ԭe��+�5�x��k<_77|�r>��c񷔼_������3�����\J��B�v|�~���vnLM#�αs:�щz��;w�'�1��k�w��c��8���.x��qƋ7��.�|v"��!p̡6Rv��X���C���=�f����̦�=z�!��s���%hB�uo��|R"Nd^`fU���3�-P�mݳ�*�x�#�r�摖�v����y=��m|���#��=� ����U��P0����{�=��|����}��r\6r�:DZ!R������Fu����u|�j-:�a��meL�"9�
��PO�yխ܋R@ÑxcYy.���Q'N� xp,^��(���#L�t5��V`��EDO&�}�K�;������'�?K�E��������b�%i�_�srF�$�s��?��^s͵�������^�Y@�ATSC�����4!�Rq��y�� i��g.��z.a�!�y������^�^�	�X�[}>x�E�)�c�.���@�H���\��#��Q�
�˽�ƫ�ȥh�B�<��2�����(��<c�g���N����o�$�g�V�>���]�9۶�k���vLʡ=�׶�3�i�͚5[B2/ӸMH͋��sfW��ϯ�.]ҳm������^�������ٯ�|e"�$�/X���/�>���L\x���J����������ڽ��W$ވ��wH�1��}��X`�7��kM��C�x�5�o�R#�m�f7���Z	��HltlԼ�f&���B�Qu���_�Sl8�vֵƃQ�E"lg�q`�\�k?��)ԕc��`9s
�(j�8OF��\xO�tz��6KTǅj���K.�#
|b{(C��f�2��!��/�'��
��bf�1P��
z�d}
��w�s�
��v���N}��k׮ɑ�ϯ�(?M"�<MXB߸q�Z�B��(�
e##�R�>A^^�%#r�%dο!D���PS���)����[J�*��PIn��+ć�	�@�f#�x}���=�eD���N��T��Q��*�n�6�lH��!{��*PE��7�<���L�|O���fy���}�Q�S�������_��mx�$�MT�O�t[Q��9��xJ7M���pžif��~��4�E䎗N��Y�v>�����[�YcWל�C=�]��k��4��|y"�$�KXB���~�Z̦��e����Ik{N�� M�����}��������.�TdHxwb�?H)ګ�mj�,s���z�)��Wn�Z��ܭ"���6A���	m�uq�1���i�V-\��6<u���X��Ma�Ӆ�-lTҡ>e��%�o�x�λ�Ex�{��g�K���1����/=�v�H᪚B�ԛۤz��^�5�Q�=zM��鲘|v�[�<ϯ�YZ�U!���Mj�����Q$���˵w�ҝ
�����W���3'�,^���}&���$�@"�8 s�qޤ��M(A�A��o��A�?�-��L�����
u���Y��H��XN���׈�C6��q��Z��g{�z�0/�̥���pp}v�I�ׄB�%y�$�6�E�����=m��1]H>���h@�*�CܦL�ظ���M�.�1d���k�r�:�l� D=���:ǢՏ�9��14��&,�t*MYS�^��ʛw����Q�0M��y�7o�0��8��	I��\�'�t�>�Ν H��#���Pq��i�I�6)T^���'!�����E���j�%��n�E`å�΅e�l��mҒW�q#�Pf��d���}^�SoA���
��B� �0�`���9D�;�#Pq1��a�H?ȼ�9Fh���0�'c���z�f��%�@�����Э�*ަ<�1-U=n�î�z�*����DĄ�Q�ڣ��l��2�HWD�� *���蒤�+����fW��}��M(��Mmi��4���$�@"�A��$􁁁����*YqU�^Hxύ���=���͠�Fߐ�:dj$.6��jx�}��;��%��(��n$�'y��p}i�k��k�:�.�i����Iq�f(�ʣ�[cy|f����k��o-|z�{��,Lna���Xg�^�O(O��g����o?9�%sy����֨�yp��\"�AE?�蝪h'o�O�]m�8�۶l�8�%���[~�͏�
N�D �#p@:c��C�~Q<��Q��K&:�zA�箭ל8�D���KF���䡒_ǋ-��ȉ{�����K�&�R1��m�B�cQa��^����5A�/z�M����+�9�a^�oJ��o�4vo���Z����-������j�{�"2Hs���<��.rv^�Nx#����0X,wN%=ߝ^׮��vS��ϸ@��o���Jr�w{��o��������D H�cHBW5���Fr;Q�Y�� �h�
O�HE�_'vJ��������;F=ͺ���x�"�AʋaM��J� n��7����x]�L#��y�Dd<�RZAڎVAn=�z�Ye]�y�JҲ1L%�ۊ����9y�5#r�}�.Eq.��E}�-F>�gg
8���f����e�x}�*�]��+�=���Z�9FK)X��P�D�j9Gr�=�`u�}�~��3N��?��w��_���D HۯDD�YXxC;���+=�4)BQ��o:�3�">�{��O��[������.�O��s�n,D��C󑿏�"e4kDC�����P��(���Y��bލ�Ѭ%�O�[�ɏ���s/_���"@ΐ|6�GDz"�)^��10tJ�?���g�V�@}�*f����9��1r��͙�mQ�~�j��;~x��_������lFu��D H~:HB���{xdDN�k�GkZx�x�Ѷ�z�(��.Z�PS[�F���t��:�F�x�婽
=���ժ�=̯i�5=�P���~�r=��U�h��9�;p�P{䟣h���X�R5�J�tU�s��7���щ  .C�����u!G����az�_t>�Ð'.�O�J��z�+�`���F�G����0�=�rǹ����iV|�]{G��1�s�°����{�aG���[[e$�}xۭ�8�����[������7��$�@"��./zLĦ�A���$��� �c�#��O���*m<�1y��x�&�
kފE��甽��g�I�}u���.���z>:zν�܏M����!ߨ���xLE�}}�//��}LmmV�^"��N7�v��G(���1ˍ�|���e:�:�L��s�\�5�1�U�M(��\b����@��\��9s��}�r���i��ιE���v����#��eD�}F��������}��{�9��<�D H���}��1���5l�Z�O%-�,z�!?y�^G�R��}���evO\D�:�uR���Z��ApEw�1B�3�Y�ޏ��8�B�E�=�(���n2
�|u'�_��im��%_��d�@��6��������77�?�� dޣIaoZ� ��ŏ�y>�@]��Qy�I�:31��y��l֪�s����u�}��f+��gX���n�~���&���p�"H�@��$���:jT��A���*$�8J!=��	oV�)��fUU�F�G�>�P;�b<Fo��7�6��,��s�WSOo7���7O��{A$�,շ��V�{���F䠱r�/�r�F��Ň�T��C����g.]��0)� Ow�^U��'�a��)l�W[���=��� ҥIQ�7�+�#� �t=�*R��^���P�B����z�����{_�+x��9Ȝ$w�;kf}f��$���R%�����n}��;�+9�9�� ��$I�*��u(T��ѻd��Wm���;�r��,\�!���ÀCٷ��/eלƾ(��q��F1�r��!��i�?����_יܰK�u �*j ��.�wԧ�0�RC��zQ��*o�G`��!2�B�ݞ��d��[꥘���2�dZ��N����,D��Z1��_��÷�V˸E�����f�q`�s��ln�����Co/?�<��<����ƫ�O/D)[�G!��>h���33��)+���'�g9ܩ�3@u�O��6���H�*����6Gl�G�P�Ҫ��Tg�W0nf�IXd9�"��9�h�YY��}9�cq6�E�7~���W��IY �����E4��ͣ��C����L�1u�V�d��.��"7�i�8$c�b3���n�<����$S�;�F�RV��m�h`|=����Ǖ�8`κ��So�/�aO�@�9em��y	�3��g���\��٣uw��R��yBN��^AJNh�Dlޣ�ӟ�>B�$".�.��Nj�xG~AaLX�TR�q�8 �jyd9�H `��#��c#v�`�sH���?���G�?��$�֐D��r�z�*�����ۈ{F�$�S_��#&�50�������ư�w6j�F�>�p�mp86o/��pw��E>��)l����K�����Q�I~Wg�Z1a�6�n��~g����V�ttr�B�`[&B���|�`��e����ޢ�@qˇr7�8k#����]6{'Ŭ���q�vti��������,��L�_\w1΂��7݉mPe�\� �Y�+�t�n��fw{�<Q;e;}��	���Sc�Hd�]�f�y=�=�^U j6r�%1�^�Yۛ�3^��9y��Ý���7��SGkO�а�s��NjZ@�q'4+��[��q�S��f����C�Y�VfF����//>v�S�]Iu�}��R��;!���]o���a�.�C,s���s�4��C��F�;�Б�v����2Շ|�gѧ��aڳ.�!o��k��0B���1�O�����f�S��Ry)�VE��Qrc����INiގ��Ϛ*����fY�%$^ݒ��w9#�ݟ�Lsd�B����u���-F�㥀Z׏��f�~z�1!P�L^O��`�,Ss�B��<<��|�t�j�
��7m���'��ď�	�#��9~� ;ѐ��x��|g'�e!3to""�����B�{p������@����a���q���w?��h؎���A���C!_����_�^r��s���މ��2�w�D�ۀ���	�H�q��Lr���b}��|�>�`���&R����P�!��g��r��y!���\g/p!�L-��Q����J�5+w;�m���\|�(�a�s��M��jhD��0�*k >ȷ~+!h�e{��z�7mh�!E���\�s��z�o����R}N������!}6����
���sF،�+�,%�Q�]yKA���Oq����e�e-N�2/�����f_�~�p�5_I�Z�N��j΋�X�ش8,\5t2C3>���X���^[oD���
�R�V�U �����U�D�NZq��Yğ/��ZЍ���-~c�CV�N�P$�Ч�������Vc�g_�S��G
:��KĜ'u�'�k=���H@F���L7=�&�0��*rs��C?Ʀfǎ�e�Y��ف��9��P��fŁ���T��U����`�-K�ȱ�_ �}�)�2��Cw�Wi������0�[���&���
�j�!�J�(�A���Ѫ���ќ�9���Z�V�,��M��&t��A�ye�i-A�r�8�49�[4#\�}FED�<a^wܸ�hZ�!a�sJ�xSQQ<Ѱ��W���c�E��>!=7W��(���|��=�L�Nm{�}�5�M>��{�`3f�wͻ[��[%bNӜ�,�+?�1���o[l�ejY��7�����a_�����#wS�s"�vt1��A��r���z%��Jh����� ���Q}�n��0�w�!)��^�{wQ`��S�xa^�	�E
���7��R����{Y���g,)!���R�=�e{���l2\�۷��?�%�?��ut�-��AUJ��o��%�5>G�| 7�}>����(�:M�*Î��^��Em�4�Nَ>C���=��=i�WkSŝ� F�V-�};���<�ſ���}T�y����#�0z^=c<�����y�i��S�P��Ε�ay��׶�e7b��0�]Ȯr��BЩ��y��&�����2d�Rg�-�:�]��p���P1N���`�O����F��]K/g��yyCa���!��lnܰ�S�.M����FDR�O"q�bK��o��.�s'���)z�s��G���rf�����df�E�ЌMY���cb_8�#��������֏�4݌�|�iW���@9��c1Б~eW����%����Hg�y�H�QeN$������En�� �ᜃ��#�N� �������&�H��66�!�5�g��g�1)�-_�я���ɝ�o�f�(ԯ�)}lx�hU1��.Y��V�Y.tB(�* ��+Kc\�㐐�����ڄp�f&����?�����E����M���Q��P�*�Z��u��$��y��nL=��w? n"�8����������x��ᴊ�tCx�;yGu���ތ館x!LgH5qS7o+�SI,��6ݻ��U�xGx�e��ǃ'K���(����.����2�_���[ƙ��ެ�-����_������x/C�!n����m���7�ua��x��E�n߇��{�J�7)���py`l ��L�c�)�l��/�=D" }GY?�}�C��]GJs�C�#�,y��	��^0G"g�4���>U��D]u�Z�����&�Fǈi�	��-KG�9RȁDH��&tQ��k�m�LH1���O���3�P,Ş�h��nоA@���c'�`i����# ��:\�6���t���!��T��u�O�ܒp�!wC��O�����)Yk����n�h1=��kz��Y�7�*�Xĉ�7g�d7�����7�%_�a-����o���oe=�[쿻z��Ô�$�E�o�Nagb�i�C[�٩�ޢΓ��:^L��h�K�c�)�d@�Ǯ��O|ҏGH��Ľ~;'�`k����C_UyԷ�+fr���v�����vU�ٳ��X���ܽ
����T�#�u�.�2�̗4� �{(.'gXt�����uvX�z�z �����ޚ�ԧ�����n��+��FA^Lٹ;A�����2�rѰ$��Y4Ѩ�b{�7�I�pg���>D�eZYq�ܓ�C�Zz�n=�[�}�Ȁ������?}����aB�5]E�nO$��g��9�  ���4��lV���7�4݊I3 {��MO�~�(^�-� ���.�ۉ���pԖ��G�6�E�()��
l�S�{5/}��fFA�v�Ynm{��[�r�0�jH$��f�֑��ﻗx��#st]��Ry��+�F7#����w����Q�j<�j:�
|,��	M���r����%�������G�*��74���1��˼Y�Uc���;��n"�-�GEʛ�_�E�OO��ʢ������S��?^��"0����Ϧ�Z��9�x�~��A����&�@�E�BR��3��+d�+(_�L�}7GP�t�#{���y�<_
6�E��6-�yO��9k�C;�,P�d�U�{�QM64�m�`� �G��~s\�<j%orYeh<�b��a51x�Β�OIP��t�~Wޱ.0�OT�*+-��`�K�p�zЪ�g��4\M�5�JEy�$3�n�j ��@Jp�7$�ǖ#sz��BO�w�C,8�qX~��@.��^q	���g*$uD-�� B� ��xK��1P�pS�pB�^A@[�m:�|�ǲ���� f����QUY�EUg�7����c�}�7Y��4Sd��~�C�ݼ�]�M���*X�������r����}��oX�r��&"-A�
�Vy3��3�	Ƴm�"jL<}Cƻ,��=���Q�5*im7�3c�������y������gseh�0$�5���jS;�-��y6/�l�y2}��|}��62|����e>8�켰��V!-
;H�c���'ҫv�+l�n���A�@o��V�b�x������NU(����8��ͱ��,C*�ݢ�1������l�Mq����C�)D����.x�,�0p�0���当�'�j�̐�b�<`�V�����zK5kDuD5��A0n��6�D=��E��S�0QG�0��I�0GW��æ�4��b�E]�S����s� |m�T���؞��tw��x����G-_�ƨ�kX�\���&�4��\P|�R���t�iW�%u�K�뭝�����Q*��êt	�+�S{�_�d������.��+C�%�K�{�ٔ�����B�Rθ�T��*Ko�Am�&ݠ1��i������+�,���`q���y;�S���*OM˨�Q~��Y��ԝ~��RTᨰH��)���h��3B̂ ��A1Wm �6�tE�]�y�B6����3������a�ZXj��8���CP�#�����!��:��fN=���:¦��j��>c�:󝉫�n&	l���b%W׫�恬�1����~g����+D�nU�^���O�=�����n"J���P(��’�S���r�{��܏���z��A�2�����44=:˩ٳ��J�dzSJ���U�r���Gf�p6$�
5�2�~�d#�)8ѩ��8�|tΔV^���-s���3	��RYbW��Y��`�"p��]��,ٔ�Z���^�E.����Y������=r6�Np(��FԀ�!�Ϡep���v��#����-(�'PA�|�B'nIN=m�Ndq���"�h���:1��2�#w���loBeWS�M뚠�s�������	��D� g`Md�e���R���H�9��ӌ�z�Ӎ�m|%�g����oBmT��K�Fٹ��Z��RX�H��#>aρ�&�>�:]yߚ�W/U�Q̒(W��{���4YŚ�����|�M�VO�ʐ;;����ެ�(�R֊8��� �"�Kg���T7]�bUڤ��Ї��R\�����5x����	���t��)K��.���}��:`�q�ƣ�&��,ߕb�'Y�?{-��4��������$� �jy�a���S���Z�C�xS醒|ثd���:2�ѮPq� x_��&�d^�*���C�ԍW�j��y {u���'�o&��^���\Ts�d0�ܲ����e���/�E�����@�y��)�P�k>�c�~���`X��w��0�'�Lְ��^Z�'��'��gf����z|:��/�Ԭ��ߒ�D�2\FyL}���s(fn$���ZAe���U�n��k	�55�c�R�n�Cʀk֐���4��LrtT�����ih��߅U� Dn%�~<N�N�G��px\/���1X��)(�h��}�|�!�Z�W-�ӯ�]a��6�7���C���3,:��?�Fٛ2d��5�z�o�e�~bZ|����'6#̫�����^;^���5���N�:/BM�:�4@�����?{�<K6���rf�T��lY�l���h�$��;^h��`h�?XT�2X�608���`�;/�� ��忎��\O�V}�ۇt�����y�*��mo_AZ��Z��#}j���$������ƙ��Z����m����s#*��FQ��ǹ��e���7���ߑͦ�~�h0?M���	W�.;�Z� *m���P#'L-M��-e~��k%��/��W�Ċ�q���l,�qZqd�j�Q�mm*C�3'�6��m�����I���ބ����M�|���/53�����͹7�����<�<Z<@}Nu���g���]|iށ�a?��I�����-�9�c�N��I�
�i\s�2�6+����"]nw�(�����c�%&���6LQq/q���Ffǁ�8y|�G��t��w�X��z���C�G�$ݭ��W�7���U��G+�N�,�C��fB��oݲ_���H>
S(�m�IH��ˬ [��e���{y7�[���l�S+C��A�e�4�a���duh�%י�fB��Cߌ4ܡ���a�b�A�$��*.�O�^�c>�xPnAU+�JP��;��@��7@��8z;E#�����.m����o�{Z+u^.�(��L���(�k*B��tL[)nh+ݳζ��axJ_�����;��.4!�ջ��W����S��0ɀ��.���©+�E����Ka���M�k��i
_Cs���3+���)6	x��͒b���'yRM��eu+�×�%��gv[�߃�[5�c�z�wn�a��6�I�fr?ۋg^�|�:�Ϫ?��	��-���a�
�Y&22(=�󛡟4L����P��L�bh�a;�f��Y�eot����U�:��x3���E���o�Ө�/��K�U�����tPٕ�c~f�X����5�������b�@�d�B�i��23il�r������9 ��!�p�9ԟ�N��F�9Ż�%�R�S��-BC l���u)8G�J�v��$���~�ML˔�N�V6XYR9꣜2@���r	Y���5�c������������st�"�����He
Bʞ�w����� ����p���<C�hB�-�hG������H��r"c��˭..!��5�Pޣ|�Xx�R;C�b���W��6lM���:��6���0#�~&�1$�o���ȴ��9�uj�#+b�_f��[�;��P&����8	�������(]�+o;�l��S���y��[ڣה�MLϔ��a������Tj���,��������� v��� ��P�FgnlI#ad���O.�E!.ڮ�ɛ���	�t�)�?�K��MH�AKxx�׻:*��M�~�@TF�-���Ր;l�����2�f޷��y�mKeG��/�Vl�|2�e.�)]���=�j?і����5�F�=y��8�)+�����np3š\U���Ϯ���x�	4}��񌦳Y�Η~��{nC���,�"ө���Hl�sQ��c_@،�f��u�Z�g�"R�������㍤#���I�Ġ�����`b
Yz�1�l6%���-u��Z�����$2>;�R$ts�	�o���t�%9<V�)����|�oޯ֣�laJ��ud-b�?���|)[��C�$"��6Q�w�s,x��ҫA�a�EU��d� �b�e�����޺Q: �"wW����T�{��劢���|%���עY2�q��*�nw+����JRN�2[���?���-r�%�!{뿓�[Z��js��g�������/h)a��E���e�M_I>Ҷ���\��,�\>]�xtµ	�y�j,$u�M^��nq��O�u��k?f� �Y���Ǚ���-�9���5�,�|Rw�� d��lۖ��g��C̦l�{�E�A���;��1��R�qd1ɖ�/T0F,*���P�����w#�_�����gxN��˚��hm��~=d��f���w�����f�����ĔKm���>��b6Qb������zq���hױd���t�w3<B����#8�;��}�S�*��%S����IS�J����uO���9�Tm���ʍ�������!��4Q�wT9����1"I�lŝ�]�2���`�	�|���p����f�̣���蒕˳%�$t��j�NDdw��.V�������q[�����)�1�����Si�����;אmk�k��� �׽��E�r�
�-?Ô�A�V�<�-�lP��wjƗ�{�µ���xP���I ����;���߿�y�ٹ��fo��-�s��y��p�U��2${.�����1\�m7��
M>��el4���'���_���j��&@g\��T����%�g�9�ߊ��'���[3S����J?!�m��f>���/s��2�|5$�jxR��}$B���f�0�����$��i�����Ex�:x�v�=����DVJp��kD�����Q�o���հ�y"d�_hc��0C;*C�|/���	�E7�6��I��Jw\�s^��)��E�W�"]s�,��K?l)��C�e��i���,zy��qf��Xi8����y��6������[��P��:���nr�%⪘����u�G������\��uL8��	��"�&�H�����4j5|l�kۜj]X����!+��5�2v|5�W�S{I�jLe��0�+{��@&���=×"g�j�-��d�Es�T������>=�i��)���k�0ɬ��n���4n�/�*c�|��R�ؑx\��ԛ��t@ǯ����ۻ�c�DV��Ãm1��(��g�=��e�W�",�F����a�;���ڛlx[���w��U�ňڟ�[��"sW+��K}�=5��?*�y�MƠa�\ �x�J3q�Ayc�
jG��1hѵP�2ȼ�~/&VY��R�J�v��v�L�C��f
@�ƅ����}���s<:��e�t��W���1	R����X�t�������g�JQҥXzx�4he��c()���(��~���$]iȧ�˖5���t�`�����ފ��q���Y�J��[���a�Z�K�;�_��U4�7е��?�u�x����������N�q��83��7AW��r~=<��A�7�S�4�$�A3���J����\cw55�E:�B-�Ut|�u�G�x������<C�S�����$�]������v�B�qY��԰���Tæ�3���zn��F�2����Q�N�h�f���L�78 2n���(��X��M�][��R�_F��D��h�����q={8�鱆��ҮG�d��
qS���U\z2���ި�>ݦ��RI� `9"nģK�0w,�2�
����f͵��J_?Y˸8�,��LO�9���}Q.#�&C����[�NҔi������)�wN�r���ѿS3b��B���Z���!VP#��|Z�[�5^\��E�EL7�jW]v�O������y߾2�X�*0i3ؤ}$w�����=a`n�.z-�t�ʿ�ȓy��%���N��^UY舀��rAY�m��#�[wx	��bv��~�{��%Q7ӟޛ62I���U���w-8o�j��e�z8�
����z��ۚu���fݰr!�|�'�U���p���I۱'~���9y��"�C�>4H�%�ֿ	xykK�!V�U�'*K��n����D	�U4]F5M���!��ܫfr�O;}a�K��K��8yo���ط�\�\++�{�l�b�D�Չ�A?L�ѓ;�C#��Ҹz �_���3Uc�������e�SD[�)+�Fy�§�;]���;�o��>�t�R����by��ą�h��_Ǒ���G�S��V.�@���c���isl;�����*9���<R�(S��?v�`��g����dku,��9���!�c��Ox�M��̽�����s,;��<�
J�i��\
:�����+�7f3w�/�x51w�<0*ס�G�Sy���Qs�� P�Q� ��ڟ�ܼ����S�����VATw��ϒ�<0g�PR�<Y[&c�ƮK�a�D�T�E�G�^=��I	�C�}���B�"�}ŋ�Q�9�1�d�Bf�:�[�;yE�b3JXEe�E�����:t�L��L���ä���vj��r��CW1���!x�4HC�ĭ���׿`	�$BB���|^Q�����z�Q�3�I9��$����$~Ւ[׎�ۈ��N	m;d]�͙ ]��ǋ�ë�������?��%���h�",������Dq�j�{�zQ��1�a�.��>�3��c��n]$qt_��O 3��7:S�
�:��Y{��"7��i�����g}�^����r=K��i%eI٭q�p������+J�F��p���SC��O5�y}��Ee�K0)�ԛ�-F*�1����"M2o`�o����U�N�Z��Aڃ���S/h]&��L<�nQ����׀{I�V"�M���Ի�ָ\^�o�v���K�4moUX�4�l�]�":�Q������_�S�U�q�w� ��;��%�{r(eI�'�EW� �ؘY�[���[�"��yM��J�7+R5�*	
����� �3�cU��XH@��nF���/"�z/mt	Hke��f0g�� .\h��"�z9[�ns�D�[�pي�*5S܉�,�b/1�l���kG��t'����Ǡ��xd~e؀(]�W ;P�@��,E�C��g�Z�q��@X�Oo�/)'c����'B.��/O���p����R�U��(���9]D_���؈1��l"�5I��&� YR��mu��]��!���?�W�ǳ?�U�S[��$C�@+�ݻ�Bi
��;�v���j��l�&AX��`��L<���#i�m���c����v�����U'7?6�����̨�Omu\��ޱ���x�p����e@���a�	�qk�f����C=���=�)n���|��@��vT OX�㏏"v}�C��,zU
�n�M�Nj�r�\@j3��/'�D��OT��@$���d�v�Q��m
���C2.���2�ˣ�f�2p����r��[G�fd1L�΁^F���\n��Y�@�=������3�Y��1�ES#��C���'�S9�0���/{��~��s�^�Qb*�AwҦ�O`N��Bk�>#�&�D4S����E�EP�_˥���� #B�E�д �?�;D�e)@t�\�-*�51Jyp���(7�8���"����z��'%�;��@} ��&�&�R�����]��F�o�_ז{>�G�a��#�8������q���b낓��������/�=��[rq+�9wR�<������u��q�>E�']��[�]��g�gYBd�U�\5�B�1��E!ˡσջ�w?v,�R�
����<�}�b�$�f�K���b���q�d�OsH`
�WX��$@҆=�}{��K��)2��h}����d� =�� �gv�r�����L`��^��o�gZc߷w	��P��~X���&�R:���jˍD�MK�2�b�B��n��o8?�XH�&z�?Y��3#�d�YH;!vy���9��|��:&�šw-�@��t��[�Cc����6�+�T-��t�}d�o��O_�>��Bi�G*}�LA�@���ێ�~{� �Y^	�5��pp��;w>�D�x*�׮�(PS0%�Γ�wR���-5̰"YA��-��[�QfՉ��9��,kŴ�������4x5�e>��q<�>�G
�M�3 6�u�z�?;����HuiV�Js(����e�ڻL8��^���xL?�F,$ZV�,��y��pxpRG?��B*v'}d�����䉀Ap�O�rѧJ�����~���z��m�S��X̝%����˻�b��go�m��M��|Rlt,[������5a�R/�Z�{�j`2e�cK�|����nJ��l�\��,!ˀ����s�{�fQAdӍ3�U��+/I�D@c���~���&�J���968\�[wH�P`�2���e �(C;�/4�y/ń�i`)�o����6�D�ঔ:Y߅6�j�����c�;I�j��z`oPJ�����2��~����o�L]Mԯ����,.Ba�K��?]H;��tH��H�����µ��?�n[k(������|B����!�dUvuC�õ�S��{�5F��>��6��<&��$�����uo�]ؾ���&9�Ɲ�����U$e�KN��T���W�RS��R�AV��Ƨ�c
�y2\����b�����6'8�s�4	��ڗ�Cc� A����ߵs�����T%�ֺ*�u�pF�D�6~�￶Z:�l��6�W�C�����%��?������K������m�G�+1uV%vT`�ژۢG��f%7�?I�'Z��7*5��~̶�������=�ru4X��;���}�˺���{������'���ޒ((ΰ��1Ӱ�C-/�i?R0?�J���8���AR��|�]5�B�0�s<x{�ǒ��j��Ke�O�ܹ�]?j UV�����Del�k��[ `���q1x]Ⱥ��`o���LIP�ej�w�c�2a1अ],��%�Kݴ����nqL�3�^�>%�l��u�6cH��ږ����=&�.�c�,cD���ҁ��9bZ���i�Y!�� �%!�\�f�&�>kc~��hF����0-|�nS�+�������>ld�0�h�mO�Lc'����۲�R���ZM���9dR�I���c^���"��,�&7�
�\��i���Ò���U��GA�&J�����Մw��8��m65��a�	��|П0ʇb��6w4,>w��r��񔤫x��5gV5�}dJXR�� �ղڗ^��y��S&�\3�Iޣ�o��I?�B��W3�!jP�m5�J�Sq"W�xy�x�Ub����{����MCAn�d��HPo�J�m#�1㲷�4��	23��}�[�a�DV7H���(����a���^3�8��?%�I�����9ۉ?i�c�d�a��+]�0���V>e[1��]�� ��R�W���y(\��@���Ԗ�����(27�����|����>cYFa��}�P|lO�Ӥ�-bW�}~h2p�4֏�,���H�����Ѫ���e�I��|0�|-1�Q%��YƧk���E�Nz��5v"�O��?��K�sN�2�Pg:�CW�$�uaS/����|D�Q��#;;;�H0D=����;���?G�關0��l}
��-�j�~��;�lG��3ǅ�$v��"LUX�}�=IK(�]�b�Y^/��G,����W�TGH/���k(�YR֞�Og%��:m[@��b�*���J�6J�v�3�ƣ��#C���.�ux�^�mO(:�l��qϢyT�	 �`=�Φ8��1�6��טF�rA��� �w.�1��*/�Pz�e3�{�������Igm"��iZ�n�0����C�$�=�P@�Ȼ4�?�˿��'1L,�!��lR쵑g�����LXɃ���V���hd���Q��A䠥rVT>#��?�J5K���V@�_ۼ�����i!?˭��]��W�e:�䳶�3���K!2cV���U/��|_���ت*���R�埙"��s*�i��]9o߉I�Bϣ�g�Ň)��}�M��K�y��k���U�<�d�<]���HW�&���N��V�J���/͞Y��3�l2�\eIf��l�~E���F~�ζ=US�z�/���s�|?�?���w[b+i��0,�˃��ǌW��F��4�dl#�u�@��I����	/փC�\��D@����'�Kl\�v��!���I�vuًIqǒ`r`���;�{f�s���#:�=1�*��)L<��,�*����?d0l�[���ݚz����̖�i:2:�H�<�K��Z��P�R�:�Q^LU^�z1���i��$�g�����+�u]�ǈ�޾�����3^�l�u_�2Ugz1�ɠ�r�)�� �{:�_�J*�͢:Sf0�v���g\H�7L7S�4&�U%Z����A���N���'Lj�c��dkP���l��1��yx��xd8�K��Z�_cXBs{�*���s���ܜ���q�&ڐ�RS�|�x�*6☓���{�i��	�,Z�ە�60����U��l��.��X�b��m�T~��|����'�"�o٦t��!�,�A'��~en�?�読��+�SVd %��(s³���T� \�B.W�,�P�����$̗��)�i��v���z]]�G�Qd\�V��&�tG}��P�vʐ^�Z���x���ʯ���Bv��Zh��{�zD�Y\5�>-%Uqg0p��/��į�Ǉ����"j���y��d"�P�n�M�U'PS�9��#����t���5N
Q�S��y�����T��23ƺL�Z��pO+��s�[���`L��5\O%2i�^��,(�%4��;����[���yH�/���4Z���#���u}��3�"Ѷ�4�:�+��I�N	5�ʱ�����d��J���hM��s=lQ��$Xgk.����y$�I�q��H��Z�t�� �W�/�fݓ*�8]�����Q���ɯь#�Rt����)�:�:�����PZ;���κ�  :u� ���Z����X�٤�E�}g�Hs���H�e��5�:��8=���gt�M�k�(��Ջ��Kۯ��!h���v�����vQ��t�Y�1�V����钼;��!��1��S.}/��)�i��˱��#�3h̃Q����> Ѩ��J�?*6F\&[����_,�ɨ��)�|F��������u�Stp��9v�N_��q���=R��8�!���v���"�E����P�jʨO粡��%"�����fa�v��FDW'ǵ�Z��"�TB���'pm���CJ�ut-�&dPr�&��$�[�������7�49=�1C�dM`ρD��'3��������x��i)4����������3LD��~�klDv��\����⾢�ʶ�dTb2�e�Y?�o��츁9BY.�����,�%���Yc��pkH(TSm[3�P0m�\���_�V��ޣmh��d&�W�d�["�t���=�Ǻ��O����l�'��RK��[<��<��; @4@�}@�8�6̜;GM`�s7���6�b�co����:�Izު(du�l~�V>r��I%�^�� ���:�*�1͡�\�2�sc��w�3���6� ��!k�d3��kv���W��/�n�D�{nI�]l��\��o@5��<��W���Q�ۮ��o��=�Оqߨ��M���P�+�xB{u�$$�=`H�ZI:��'�P{��n�㲸�ꡬ��O���g�M*�~T�nuJ�uT1��p�E�͐Q�F���ћCɟn�����ߙ���`o��K�f�|�S@;}��a%��+`���Y�>���	J��{�=&]��>ۛ
7����2G[�wcʘ���\���E&�;�H^�Ԕ��ᐪ�FN��Y�����i�;a����	Rl&�Et¬n9�ٹ����388�z�C�N:l���-�6+"#�&���,�4��o��q�q�>�-���S�/�J8�-�}�6��K�/�S��|0e����;�hsQY0]khJ4�9���NY�]���(A�����"̬Q��+���u�{>������tP�鄏�9��w �a��+��n����_u�*�>V,�x��QMY-��a���E�I�����W��l��*�2�������@cɕq�QL��ԻӰ?o�_�_�_�_�_�_��5Ȁ�N��[,ԝi$9�^���JYK�L���PK   �cW�>|�2� � /   images/2cacff52-a01f-447b-a47f-67011eb49dd1.png̘Sw%
ӭWl۶��m۶m�cul�c�c�F�x�����+�M]�]�s�3+FEI	   ��H� �  X,�i�4D  ��V\\EV\�T������ ��KτQQ��	��!������:���/������������[��������2��vb���ҶK6��!5G�^�FN}��u���r{�=��?︃v8܉����QU �h��0���Nj' j�-��B&Ө��D���q w�أcͭ���gl�H�, ^�G5iv^䅇��j��ҍ�}��p���B!��|�cn2U��\F<4�P�a�`R�������uR���{��,T&��t>>^lH�K< ��W@�ᶛg28.�w��!��F�3����������^J2s��0$���	O�f2ǅ�4�V#���)f$�F9B|�YMP,������/�z���ߑE�N���Ҍ˨�����ҙ���*�lRMta&:�hW�)�z^>6��հ�Fy��䗘k��ß��^k��c4m6n*v�&�]�/16>+�Zr�Ѕu�-���[�Z*Y��e̧����#1�y$�<SzZ�X0�00�pR�>�l�Q�sx*�.=U��L\�۞����.Xȭ_~�3�',[��6;3�zV���m+�+	`VP�TО]FB̩���^�9�d�����ـ��΄`5���@�B��RFC ���� Rޏ��� Ŋ�m���ɩ =�A����ҹ��(��@�-����ǋ����EEZ
 5�@o��I�9��9P!LP���@3E�����i�]���.��¯@���+=Ez����B��nD�	�ta%�c	I=`�Aa_�rA
�u
�^��n$��U�7+zPբŎ�	/9Z����"�WM���N���O�C�m�?��8ۆ����(⤴e�a�b!��ڃ����`�Wd�I+[.7"F�����[[FV\VwVЌ?#��@��ac�����M;�?�v��p��b�N�ၛ�d�U�xgK�~gЎ� \CT�����Y Xa0j0t0�p	�
�$�����܆Ȇ����T��z	[J���b-)*:	�^�%D
�-����fRbs��l�D�{�@!#E���b���\���YN�*��@M�K�W����z��?z�4-:M:N��j~�
*\ZV,s���B��rE9*�ĞTm�~)~��J�ԛ��4'Ut+�T�c��5�c��E�T<ΡV��c�d^Z9[[�Z��2��K�g��Jo�9�9�z�[�m�m�vnб�C��Kx��x�����<����~�1=��s���ǧ�O����g������ۖ�^hM�^�fvU��M��dm�����#qΧ�^�&ʞey�&��_BZ�FD���6��,��ϭ�w��WT0���@�9nW�G��:7{�֤�#���������QI��� I7R6Rq1*�!ފ������D��
�י�����ݼy�l�*�n��|��C2���4�t��e"�Z�e�U��G�ÁE�����0z�G;��u�eNL���@�Չ C3�6�z�n�z�)����_�ϩ�	�]�TŨYn}�m���v�+���K�K��������K�
��o+O�W�&ߵۥk	ﬗ���������ξ���Q�~��1q��y����h�[g�������&����m�k�k�k������Tym�Z�Q�0�濢vRϲ���կ�A��շ~玧L7���&�-�Q�eB4B.;<<� �>�>����� ՠ� ����ϋ�(�<��<�Hh'���Ճ�.ϝ��",ѫ�������J2l����͛ˢ�\k�si�J^�p7q�(!d�i�wOf/���������(o�rlI�x�3�.�;�4�4�j&=^� Ç(ܽ�f\�Z���{W=ג�� � Ǐ	�~_}��w��~�г0*�z������c��qtV868��1_Ξd	��#�BQ�	�j�L丘~����Ĳ���)�4(>�i��1<%r�++�+(�Ŷ��cK�K7xpx4���~��W8���0ǔ�ɐϻMo�p2"e�Y�o"4뻝ʘ{ZQ����^d맿��>�3��Ȉ�40�kj�9)ޝ�^�~��ʸ`1����-H_�Iw�A�ƪ?�G�n���s|t�j�������2��Ͱ\���G�����.��]��K|Ӿ5�l���v��N��m/�-�\�\�Y<��*�_��y;��6�Sx���?S7(�LiL�M�q���Ft�[Lw�ŵ�y36�J�PoS7�V�l:�>��ӥ{�T�{ۀhwoM+M�u����՞��5� ��M��ʪ��� /��]���gϏ���z���֧��۠���+OfOO�6��Q��?�NH��n<����.��2?Cs��:e��� A����=輽%�����)�(W������̨O�������a�y��VY�T����Sq3����B�F�����W�n�.#��ܷ�Y��{&��"���7��3�]����/��9�������/�g�s���N�;��[�53L�@���>�(��_^��?���g�i@h��Aߏ?w`JQ�IL��*���K>�N������{�z��7�A���O$�o���(�H+��Av�7'q�,o�rF��X�Uw�Dm�������ǃ�����us��Հ��������d�� ��߯�4k���l�0R8���U/v_m��7��x���i܋�EI`4T`7V4�7�\�e%d�L�M�O3� ��T A�N���F���;�͠]"@F�e[}Wz8;�������Z���C�!N������>T%~���A\��~>�  Y	Q��OK���8�6�_�oİ�d��F[,�|3%Nׄ�+�9M�9�҇�:���u:՜��J��L�\S&�q�,j����s����9o�Q��� ��8`|���6�FlO����u���@�'(\� ?Vc*��&�Ư��;Bڭ����xQc�0��8_������:���K����Mw�����c$n7_��a��B�ڵ��x��S �6��T���.���q��n���Y�����O8�?�{@�������<�Ń���yS��	�&�
��n|�vg�(�:p�����t�	�Qo�U�)%��d�����9X�ʦq
ڄk�`�<��#!�����+M�F���D5%�zV.��c�zр�M|]�.,P��R�K�v����f�x��EG����|ؿ6���>���qh2Fs�F�y@�7{�vm:�j��ZuZ�1��:��F/֕/w�<)��a>@�5�^%'h:�3N�3s�����1�3 ��Av�����HM���k���*?��xݝG�مY�bt\�!��|�y�Q_�M;��qۿ��>��Sd���1���ɨD@G���~'�����hi�H�OuQ����u.��|x��5��pA�Y�Q-,�2��{����Ռ�jb"b|�QH���u'�����D�UI���Z|�M8�sgiR�t�-h�i�N�S���y�����tV6 Pv
�A}0���,�
&Ѓ� �C	�2`Oyp��Y17��yB�_���4���oF��z��᪬+%Eۿ���[��<����ب�<Bz�|(����/�?g��)��BU@��Rs�_� 66~�Y鑊�����R���̷w����&������ݣ7����k�:��L¦Gu�Q���%Y3>���Y� �?3m��c �bȘ��
��!w �#	�3~��y�א��.p$PB1�s��r��2,��-I����.�o쏸,���� �s��9
�
��� �}l�3��:�x[0�����=��y�K
D�I����α����	X��`܎,:p�k��ԗ?J�y�q]krj�#{9BU���6�t�ܥ��p��,��'�Z>!S�6��֗�cI P��P�l�aC��o}���ڝ��Y��ez�5�f�����g������-�)��s&Q���)5S�~&c��&..�e�NQ�A<|Mr�į�h��^ϒb�S�F���a�\y{��C�Q5�a۟�����w�@%1�����$�		�!�5� �|V�΋�1���0�eA1pxI`�3G�D&b��4O��G���;�kż1���"`��h)�?y�F����,��w& ���(�f�]7�3���=���;��٭�e]�PN��p,���I�s>��>lx~�2�%O3\hf�;�F2|�(@ymh]2d��ˆM�&�0璋 cҢ;��9fw�;�@H�+<#�j����u2q7��aj�/����u�!(ȩig� W��?sb���m�ԚG-��J>d.�?�eG�M}��ߖ5��.3������cޝ�Jift��W�^9,�d�=�:V_C��R*�1tZ��@6Ȟ��6���P��h"k���x�C��4a�<� #&?��˂bi=�Q��6��d!�B�������=�kך� ���W=ؔd9Xg/��nYP�2��	na3�0m8�u���;�h���#L���N!���+]d��k�7�z�Yk"�ՆI��ےDx�������+�=�@ iA��0A��Z���)�검d5�^�ɑo.X�q��p����y'��BA/umO��ސW��|�U>|�
�p���ׯ�r�8g��=XB���7�������(�xo�k��LY�ে�N�4�/_5 ��jl��h�9&]Y����ǀ)��[��	Zn��}Xn'`���:{	v��?��6��Ћ��e�����P��	. b&�b�#pw4�� qO��!��\��n�����j>���O�V��^��	�~�hPU�ø B����� �:x�a�������VH�mY%�C1x�߉�z�ox�z �,��ӄ/x@ڰ���A5��ˀ�����O��T�j�=.���fwe��Kt�=��!�A�������w�joV��`����,ؤI�������n�8��:�ߕ7�;ɢn,)a�)ן���ܻK2��a	h���
Y҅��c��*%�� �:�^R��|����T0RH�����|�+b�ԯ`aLw��~�Dp����y��~TLh�V��T#F��8�sn�|�zG�����r	�t�8Ɇ;ϫ�?�R�L�:���\�<Xo� �Iǰ�����S|im�0��WQ\�@2�)����.Z�f�O�z� �
B��9&A�6�#:^u@����6�l���������.1�w���L�����-�D
TV�.j�qJ:G�)]��=�g����%}5���a��z�"�0��$ΧY��1��7����D�(���6>���!��q�dp������H"�<e��Jυ�XLKhη�]Z�wP�!�n� ��t\���q3�������̜�$md�
1��e|�&���������8��=%�Y��T��/�IA�����Z�7����ap��dA�b]b��w�|�Bهj.30$O��V��XJ����/(��˩�_6Mc^x�Q� =&Ћ��.f+W�����3'z�1#;o�ŷ��p�i4$�W��WF�E�D�DqZ�d*�����tE4ᙕX�,�����쨇{fq��xBauI:�I���L�ġ�������-&8}�ѓ�������3�������X�:Yq�9H�̷����+�H���&�Q�^\31~��M�42K��` ����J��t,���xZZ97���蛪��:hH���D���#�p�a��`��(.	�G��R��P�)i0�a`:~4��l�2B¹���L1��[JA�fKt�c3s�}��S�Y	d� �C�3�f�d�p�:�z�����c�d�x^�7@%d��g\͖<9�2��kS�h��
��C������4���6O������jZ:�e��&eb����侺� �EO�\$^���%�M�®�f���`�6M���q���0�-����=��O OS��wC�>�pW��ǲ��K8���?���;��c KA c���{|�l�i��g����#vBkJ���Z~���ƪ�`�j����[���#D=�n{��j�7(X�%����n�����\�2�_�GC�mj���0Fp+�ͽ��k��j?Þ
iF������35b21���c�(!sYxA	������*�!LAR� Ȝw���u����r-�F��.�i�,`�~���/�� ���|1�{S&(
����G@�ń?��D�
�2o�~�1�kC����2Z���3*kM`l�S�B�&�/W�*0n5k�m�p�Ԟ�%>?����_���]���;�F�tZ7e�y��[r�wy	�+N5r�_����|d8�U�<������u(�Wк��	�7�瞃+Jl.�pW���3;֕8���|�u�2�#}Dx���D`����&2�Lz��+����������[�$<����h\p�_XѮH�z����j!�qe���pRI�ж���KԂl]��)�6��l
}�IfVzƟ���?*~�k�6�pY�2�-**�?'T�Y�n㻠��Dl�:����K<����G�2�U�΋k�|���:&O'��,6����������1é��e瓦`�:r�#d��U�O�3�2��<ȟ�r��K|�QV0��R1:`"`����������5��33������d��J`7�
����A��]ir��#S�v!����i�ݏIsLm!A%��_zj@�Z�'���o@Ȟ��BDIf����g)�
��q����1�65��>T��veA��j�(���-ll��|�����VN�'&>)ϋh>�i�����7��R����s�1�>���3.�}UO���%�!�x���P�)�Uu����iM��?�?�\e�1�c�݈�[	��I�W�F�d����P֑�!�}F< ␐�!�GbE�!!��\��WWC|�bj����x��iͦ˛�H�B_c�=��\�q�҇�f��M�[���b��4¶f�p11Lf8��A��/���N���jة�G-��U��,73����<eW���7�Or4�V�	x��bЄi�#	]w���@��5�W2�+�a����z �x�f�͆�u��Wk�=�.���c+e���nir�,�S�CQ���'-����J6�WEj�gj| �e<�� �r@�x�b! B��=T|ٲmnnv/}�zH�u�ӛ��I]��M�s�Є.�������yp��%ˍ��D�T��8����Ә�
n}�.C��/�՝�����<q��1u�I�V�������b����a��y���g�EI��_��4w��#�f���8��K��b6�ݠ��غ�À��u��Q�R���e�P��������b�}r$���J��+�R^I��au`�N�g�i{LO׶컚(��ٸ�n��F�znPu�y�U�<��^��`}��jc`�z�v`j�D����F!5�����f�.���,}��u�,`���+h��j�8ظ*��{��;b����D���'c)�k�0}�d'L*^S_!��v���%�6��C�Q�C�4��5P�g������I֍���`*Tر����/�������{��6+v�R����_�372)�����G#pun� 4��Ĝ�~�ي�r��7��\���W��C����^�����-�(R&��;�}��X�JD�܆�L��ϙjmii�:Z �n{oΌ�zcy�hVG�̐
e�����ߛ���o�R�e-� �=B{���kph��{� �˷�=5�;g��.�/�e���)8@���&s���f8̮��q��N$l���w�<;���Z7VM��\e|��������M�� �-*��ڑr�7.���t�m�{В�_M��A������KA�r&0T7 P�x��ͧ���@8���VΑM��1�k�!WC�Q���sXߴ�N�u��[���E����@���T�R5����P�#��(û���b��Y����ҁ,�ȋ�*t�6HS���\4�8	�_���ߛ���C�K�����)e�⢅��)8�0�0�xZ�OO5��]�{Vu�x�F�ț;B׉m?��"�~��z���B�ک;^���\���'6�Nފ[�- �|�N���8ŬVY�r ���H�^+L@{~���p=�>�Q�(�=W������p����/��Ֆlᳫ�����@��S�c�!��i�*T�Z"�9�Q�w).>�1��L�%��~�m�K��ri@ݼ��ԔT!C�� ���}�}��Z�:�/��u��r��>zwf����j��7Fo}=+�5→����]l����aV3o�Ugґ�\���l��:<��;��s�^@� n�)����0PB!����}J�G�����	��&繽��Lz3�R �A�sϩ$��u�SXysf����_ӂ1�}�2����2S|�k���?@��1��v@��@��H�z����*�����iM�P(�	u�Ǧ'][' ���0-W~��>f�涴5��8u1�v׆�r߳�N�d�-1#
Cu^|z�ţ���׻;��Ş��s���N��H��oB?��#>���Z,�\�9��p�w���;�W��>lK���Y����������K�P��e�S}_�:�</2X�����������J��j�n�J
��o�u���/�_��"��p෈�sG �TWb5,T����|�3fZ�/�(�t��F�Cp��g)�F��"�Ԍ�<~XJjpʐ�ML��^�B���^��X L�կ謼�Ib"��U���ɒ�Y�u���+ #����ǂ��%G&�s5��J'�W��0F��5c��a}wӉ����oP'��*82�
A��������ƺ��}F����z�~\���H8;��a�.����m0k/l<&���A"P���1����.5u�W=�Pӑ�)8v�*�~�x֭o���ӈ��yu'�q���К�3�.�<ɳ��t<���J�e@�E�X�Ҟ*���3����A��=�O�i��=#�0�`��ݠ�]�j[3j�M�Q��\�\l��6>�Gm�1�Z�~=���uTz������?l��C'�F����K�b���i��L�&��]\u(��ʬ[F�ך�l�����Cpp�����e��H�Uo;H-^�a�$Z|���Ay�^�kW!��++A�Z��FD�9M1=.��sr۬k7��+�}6��,��	[[�E3Y�\��M쭲KY�LL[-��b�~��I?Qc��F/X`"@�\�N�=�A(AS���1��w�h��~
V�$���nȏ5�5��H|�$X_��Q�KT����n蝞�sz�~�t4^:ϰg=�uڼ�8ݘ���e�U:���b���0���۬���r��v���y��Б�/��	)���8dRc=㚝�[7+�_D��.h��t��O��Y���tCt[3z<;ڶ<"c�-,F�� l7���u����Z�L*���#�ұ��}�n��tX�����J��'Y �̿~��ε^����P�
kmtd�K�&"/b��ְ���Ȑ�����~����dø��f�پ���=b޵�<�ߦq!����L�B�!��Q�N���W�$lwS�^z�U�G��o������T�wL�Q���g��r�}�L�@鋈�+>�DQ5,��ϲ@�EX��D�6v?���ɲ+������ �8�����	�:6�NCb��6PR_R"ï@:ښ%�ޤ�H4;��5��(�13V�%Eܽ���/	s_�L���������tՒmP����Ud�e �E�ZAKCy�Ц�h�E�2I��Tn��9%���a��<��E_>]�N� � 0�1��4�✘�օc���b8�@*@��0f0�,�����xp��[H6����u$i�o�q��t�|D��O:a2��ATY�Ńˍֶ��-�0��͢��	q:�8u�~�9g������Fu.�����s	:��H�v����8yE���+p����|�&a�fX!*���(#�� B�c���ZW����d�N�;68)��T�zzR���r��ڳ؁!��_�r���
|~^�oDY'�VT�1�t�=q��O:u�#��m�k�i���\�S�7�ͱ�j��ĕ�u3����n���$׊=jX��ύ�k��J�8�]O@'�ά�X���	Im������C	�YgS�%�u����jM$R͕��/�<_2��ܯD�km�|���t��*��E���H��+}��!��m�H B�N6�2+�1�b�.��Pl|q>d���e����W�i�<�^�?�@1��,�3�ƪE�~� �����Puh���+�HL���-�X,l����%���vӭ�g�}��@������}�OZ(7!�E'GYQ!��#[1�c�O~y"���HD�/��,���OH�TNm��l+��n��'�\R[2HӴo�Q?{%27�
mCއ�)�<&�K��|xB���f"22�q8R��/�`�!2��E`���MD�(g��}���zN��v��>��\y����o���	��Z�K������$*$�1��hYђ�x�sU2�
��@��R�nd���8L�v���&�o�&S�ݚ!�
_1���x3�鑱Jt,yn�ǃ��l+i}�͌�zm��I�9�*��1��5�6_�r�k(�A;��Ǒ#���F�>��P["�MMf��j���#��YpE����~iw�'���M�L����E�G�@+� �u:Z�M�EbZq��-�ʡBB��®W�o�/=4Ys�C�V��9��B�3�Xs�����.�?��j#t���䔯�Ɏ�@_fĭ%]n"S�h[�#O�Ǒ)�0"���k9�F$ϺuUW�3l�qN�A5*y%N��`��.�I.�{�ߏ��W��=i��ʗm�Z�~e̗����X��B�,Wǁ�����C�����W�:U,%1EJ�2�/]��z�q�D��y>���GT&d"�O���:�u:�H�y:dp��F��ѯ�b<<�Vb�D���dՀ���ZOo������?�?�~1H-��gi�',B`�����alP.�������_V�:��K�l��8/�l�BB��ݥC�����TU��J�U_ڙ��:����1ϡ�EQ[�Gr�S𢺊GW�D�B~a��nF���``Θ ͍⯖4[�="�AJ{6uq�6�SqLNc�J(��H�箼ťK��ӊ���q��F�:��x>���1����Ǩ��>)�em�IF
mt�@e@���ҋ�%>�M�M</��o6��1�˟~jԒ%�Qg)�Tl*8��=A;on�	����̷7�5e�[��Zk�lԫײ=�G@���z���C�Ka��s: �hy�¨��z�������}���:3����q#itӂ�=?07�����t��L��I����{>�hB���6i=�"��O:� h����J�#��/�D�[XXxl�dc�����}��8E��ݚ�z�۷DqҖ�:�8i�?�,]\���%���m^����!4#�:��v�����8���]35��%B�+�ܜY���U�:B�L�]�� ����v;D0k��pk&	���gh��XK����OX�صbW)�]&�o7Ȭ�_5���ợ<^���b��b`�{|�g�)��o�IE.�:&:���]z	���f�,�F���շ�.�׺{uW,lr���x9{���
`v�9<d,��\����ȁM0��׉_`g��PĿ�]����&-	�����\ ���\f䀜B�#=�O��1�s�yˮb�_{��f�g}�����\NP�M&�M.Kzn I"�>I����9)>��\��Y�<��Ⲓ-M��a@A�u�����{�S�f�/�U�T�lڣ*���"|x�Y�P2yR�%v�>���?����J\���� ��G������"�]����k�T������/^�/�W����KOTP@����lvJ��lr�ɏ���XWl���v��e��a��\G���ng�[_�%��k��>����c�"o��<sE��h\��w��7�(��6��L�ڂ�F���kx[��ؚH��s��L<	~\�?sR�Q?QJ��$4�H��"t���[�l�w}���z�g=2W������r��m5���Q��L�N?r�
�"��$��Vb���TO?Q�VҨ�8M���yT�*��a�I�k6�׷�,��C@�Ц�9����J��=%���!���!QyĆ'��Ӹ��LYPP�=��������5���;+2m<�A�n� G���D1Z����q}��r�ͻb���P���V7@�O(o6�W�"���˻�:��´��ܵW��̰�p�6��ۥ�zPNGXPK��'�/�Z)���gV����us��Q�(��>o�E��c�Rh�~|�QZ��<����k�\�������uV}�n�Jv.�;�;��B�<"�`ٜ
�ĕ�C��}48J��e}/�X���+�P?��h@����YSǇ)�H%�\�MG��i���t>G����d�Ol������+#BO�Ҝ�H�����!;�N]^ qŸA�b�I~7�6Ǎ��[�sJQ��R����|������[7]⍍J<���s�5��JC��x��K'�ۢiC:t�h��!�3d�Y%M��E�!T�ꗋ��Z*A�	d�"E
ͶC���?M������&����c��e��S	�{��sx� \X{.��uG�Q�w��4j�jw�s7G��]5��d�ڜRJ&�db +>�҅쪸fjӘY�>#t�><�AҤ�jYjm:A���Α�G��7Fv��ⱐ5�7m�����x~ӻ¸���\�I͙���@��_�G?�zO�z��vK�[�>=��ݭ[��P]{�o�4<*S	�k���Ś5q-�Q6C�:��Ix
�������D�&�y��Y�^�zK=���5+G{��m�C��?5��L�aq}�}R�ׯ�"��zxGCϋM%��]j�晝?�t�)9$�6���k֨�
�^-�t���H�� �1��$�4*�Ku���������`.�2��8��dM�j�У=���a���9�}wa � .g��|5,(���j��TE'�<�`lX��I��M�����Or0�j��Z�,��ON ���rW�
�.���m�Z��Z)_u�6H��e�z��'v��LTkO}�����(5�X9��G��z���r�f��ur��ܵb��ޅ�2�GLMe�L�(��Ny�L�r�f5.@0.|�[vT=͐��dZ��B��|l5��wor�BcZƍ3���X��[<Ba�q:y�(�=E4��r�_���TPj������Շ����FmB�ܼ�S���#3Cl1Jr!'�����}G:8
uB���Qg��78��K�y��E4L����h�q�S)8�����i�{U��P�}.$7up
w���U�5�mW��wR��s�U�:c�� [��UI�Ch�W.Arb*�޽�ѪZ�h ���{�ev�L�2��f�����/�"�a��z�����?�u����W�p��p��?�\���Z��ڎ�z�E2X�L�ٌ���_7ZJ-{<�a�f#E2�eh�lGiqG;m�ؽ$��W(��Hk����K�������jZ\��T���t�j�3=	���f"Gƻ媴��v���..�F}�����ł�-x��u��j�X�T%m�U-���d����۬7�����?\O�0��)���Ϗ�S��F)'_M�Ѽ�U�^g\��v�[L��^ռѱ��1���u}��nY�&lKaw *�x#+��kҸsDtq�52r;��E}�Rg���(��^�(���b�N�	Z��V�R���7u\��)U��e��U�qd������ۦ+�0چ�.�����>�Gx��]}��m-&�]�ٵ�Y�R�T�����������u��#�ǔ��l�h������P�MV�W�}��6����!�]�Rۃ�ۑf&=x��$OC�SqlC4y�N?eaBi��P�������N]8�_�Ӂ�Y�������(x�t�t9����,Ga���qu��'�þ�n�:�84��d��1π��[6�@����h:J�o@���<�!7
.��V���F�jx���j�J'~���{J`v��2sS�����֢��h)Vt����,폍�N���zy�v�;�M}@��'��2��m��gn�%TB�a��7,B=����� fj����Wd��/|Q�pzj�PE^S�|L��k�K�)6Pv'o9���v(��H�
p��`TU>A}�^P�<�Ԓ[Vk� [K���>Gh󪾸?�:R���=!�-W�c(��Ҵ�Y����z@p`��Z��l����K��v4/ö��&P� xal02缱����`$$�<�$�4�J�n�;<tm��2�aKX���)�p-:\<`\Na�A��(s�����O�_~)���٦�!=ުè�».��IО�z0��
p�h��e�-�9�ɯ��0D�<�XsX�4��ə�U�8�k�/`&��8G=��#�z �(�����hV/MĬ���kTrt�d~��|�/Sp.�sl�{��:$���,�g�����ٚ�q3�����2'�I'ߊ�P��~hՏ�x�Ժ���weW�)Z���MZf_�}���n�(��/���z9N_n��z�c���n2xp��u��j�O�F�Y�����Y3�e8���i�9����lń�LP0m0�K���p��?��a�~��4w��=[�7�9�	[�6*���q�w�������w�+��f_F�=��՚m= R��+�>���aY�H1�UL�3�9�ӑ�ٟ2	ѯ�br����á.FgM�I6N)�UW�)6���Y��	}��ۥ8Dv�B��my��`gg��F�{��#~��`}�=ВZ�G�y��gq|����+Uk����o�@����!3�����}��a��f��{�zA[�*���Y��v�	s�t�ۍb�ΤG7rM�	 ���:�CH�Uid;m�Ř�y�@I\y@���b���\��k�!��C(Ɔ�B�*�	�jJS�2
+��#3�e���,C��Ŧ����
��N�ghD�AX��<�zU��4�R|%��.^gw���� �J��9��D�	�-�_�G=S:T*崁"��ު=\��!�`D驓)�>]>��Ò�!?���|>.�w�R�6d4oc2����O���lTس��B�:N�Ai���<8��H2��<��PZ�Z�w^�$�]���}��!s�-�'s�1�F����ܨRݎ��0�%ִ&�y��nĹ�8Սm���~/���F��z�W�]�*0l�C"p�3���Hw�v��c�hגo�TO5Չ���Y�1᳚�@2��:�u^C#��T �`,���L)c�*CӯM儨Q�>,|>o?��h��GP��e��k�r�ŵU{�؊DVXoA��mn��d.S�(���v�x�ٖ���-{�0 �5V7��+�OB����Շ�>F�zf�upLgu��bC��s�N��g���?�h�� e;ݍ�����j�E�9�eH��)�T��,�M���y�+O
��q��)gj��s[)����3B8�Qӻ��$���d� $�՘��Nq'1�?0�R&۷��b�5��EE��+[uʣ��E[��0E��˱}ն�s�^-����&W���L�V�!k���c	`����0�,7����aC���5��@�y��vɦV4���D�{�6c�H�qU�Ln�;oFe7��D���2�M:�C�
�����?����x������v���,�J	��!��N� �ͅ�DP�u�Hn��b�s�H��N���`��i��(�Q��-^�G��&n�6`���^�ȕn/�>�(W=ӯC�p�֛xrC�����T�sdBc������,���mu7��g֑k�	O��+�Yxa�6ǭ�o7g�������+<=�t�6;��$OeC#�YiB}�1^+%�B�w����ȶ��*�$�5c�pT�ڀ¨AgJ���!�����lXO��^s��/[�<��EfF�Hֳ����>�9@v�� z��˕ߜ�Ět$pP�!�H�������T�Ń�p��S*���H�����jɘ �7��Ol����2��A���z�x!"�N<�B"Dt)�M���JK���ݑ��5xW�i��bwsϾ�֓$np��h��E��0&�,�5���vrgj��#~}}�ⳁ�%� ��Ed:��h��g��8�1��Q�T��\��� y�A���-�m�ij�9��j�=��t��ԇG/-�<�IINA_*����=`zf��Q�:����s�~��	@�����7>v������$��*�B�f�`Y�ߦ��� �y�`r-��V�.��e�kk<W�X0߂��bI�Sc���c��&��(0�����	� �T�:�����cC�M�U�%���,BY*(��8�k�@�mQL��~�G�D@I��'-���c�1��~޳��  �~і���2�}Sھ�nج;��A{��q,'fmrh�5aX8H�e��粙�҅t+,ٛo&s �ϷÄ�8��f"`Y���xx+�+^�?Q�;7�յ�x��?Y��"4+n� �5G|���$�RU"�)z]a>� xoo�� ��;WX4 P�#v��M��7#�S��&LgQF�R�`S�Z7����XK��̂���k��^k����usy�4��˱�<�U���1Fi��Њ����>��Ƹ�yx�9��%��[�Pe2V�-"v,�sӔ�ޫ��t�ĄEi��g���{�ZHA�`ːy�Ř�Q��^���Y��p�j�Q�Wt�e�X,r,��xWH�v)�͵̻��U
��n�X^�N��=���j�� �M �4�k�7K��X������֓l�m��n��`�`	�������9�n���k�N�vϦ�<�l>xE,�VL�3���͖�-f��px�#w�O�}<߾}!ӑ����7LL���iu��ji���h��I���b}��ݲ�w�c��L��IR\�O���̨�a��B��dڙhY�e�E����/�_9DO����lqz�*v4^���_(��j��
z�7�sU'L1]�&lX[g�R��]z�N���?�5���l���$�67d����D7đPD;��1�
b������ L�B�[j���[�w]�_��7�2,l���ҫV�JG��N� �m�.𬹡��Y� ��#�i�!��3����CG�+,_�|w��rd������:/8�V����' �����
6��B���A�=����5�sґIJ���SI�Z;C!��2s��-g�]�=x˃v��	
0Ho���`��Ƭ/۰�|��5�퓟��m޼�6]���|�4;gfJ��J,r��)��Z�g����esG'|3���7 X�7�,�5s��C���36�Wb6��cR��#%���/�kO<��FNYoGsU�-����T,pE6r��9�`m1���)@~�,�V���t�	�w�́ 5�4�B����8�����o�(5m�����);��q�+��d~X���ykIU��4=EJrѺ{�Se�;�Xwi/�"��ˆ�Às���y���gH���,y�4c��+��Č
k��e�vG��e�>��&�ӳ����`�����+I�L��>Jg`�r��W��g�������|y���m�� �q�"$mBC�0@�Vk�Yb�2�����α)���bb�;�)���f��4�V�Y�0?`�"!~�v\iˣk�Ҧ���p�Er���J�]̚�Ėi�pD ,(տ�1)`�	�y~��wbp�~���<Lnr�c����p����J}�
�4	�+�hq���lt�lso�m�ke���(���-��)I�)O���A�"��\3m#�j�/�Q�'��V�R ������K���vo-5s=c�S[F>�}�����*5����_�d�;}o}7>�%a�f�C�˿qz���;�Vߴi�h�y Q�>d�]>�.hr.|�.Z�m[7w۶��m�����<I�ry����͙0d��I�8���V�'��$�J'O�4d\�M�`��"w:����+� �����6�����p�����3���O��av��+�	��	l3������Z)�g�\/�X��oQZ�o\1}
$Q5�LMZ���¥�%��"���>oVMp#RMT �p�5&�#Gڒ�WV�����92+���J��( F�RuA%1/�R����5��Z6��@�ω�t%�	l�~ L��o�}DM�#��=T�0h���EA߃��[ k%E���#`a:r�#H�Z
�-,Z�d�q��k#�Ibn9n][vY����FNQ�_����v�>�M麋�/?�����1�u�N�Y3��%��V#9}�h��Nt8*'a9X�U����;�VD|�A[�Kf ��s���K��
�.�;I�Y Ȣk�vl� ؘ%��,
'IzL�R#��Z���M�;��l��+L)?�f�&���f_�W�1�I��� �Y���9mG�q�\`��;�+6Ĵ<R�&4aq�N���6lz���O��nX�*)ܚ,*t�k>+L�@���"���`�Ɗ���ϑo�6g	X΅3����f� ��ş�%ɐ>���ASjO��3S>q��l�X���ʜ[���R��`I�iЉ'$؏;Q�nx�[�(�?1pv��;{��ftʲ}�=Ҵ1Ǹu� y5`4�beˀז1��g��t�l f`������]��N��Y�Tw�[�`5c���n"����_ω [�9��!����ƺ���cv~�.\
" Ư�0�ӧ���&#�X=��*>0�����}Nfg��M����mB�sɖVX������)/�9!}b�V�KpҲd�C�q�WH�{6��{��؀����?}�2����ԓ�o�����[�zR�����8�-�K��/��9Ƃ	��/	;�l���]������L����Ge�3y��yl"k�<�G��?[�+��`�7v!�L[Gs�r�S�=mMv�Y�m�G3#���g���aO�����-y�F;����:4hw;mOOX�}�-��hM2g��3�s=�XLO���4���	��jKG:X�]�z���]'��u�hc�����1k%���}�C��OO'��- ��hW�� ��|q��T�tJbJT�"V^����# RIXN�X���hoUi)�S# ��[�����N���	:������.O�6��@<O�� ���!� K�9p�^	�����N��(S�����'� ��;?C�K$��J������dV��Wl��S�!�K�y�g�q7zv�uؒ��ՆOYl�e;;��Z��eo��nl%�8g��˿b�?��n����lG2pdq�����Iq��$X�[H)5�'����! �,�R'a�h
*��G��u��*������њ��
����o�K��	�aai�0EtB�@�R���/�o����S����P���Y&B�3�	�W�����<s�n��m���|m��ܲT(q�*��5w+ ��b�-�R�Us\αk
L��j�5Ү��oC����`�B@J9ש��I��&Y�Ҥ%��P�IJ�VP^c- �
BLI��B����.�c-�]F��������^����K/�'��S��V���k�{bq�����s-��KM�O���U�1��"e���p��+tQ=���;T`�e�E��"����W)	��L�P� �F<���342����	��9���R�����\��B�@���乩J�V��2���)��oQ� Y��"5��+����Q�F��v>��~�����l<�'Yr
FrN�jƶ�l߶V��Ѱ�������+Y�^XF��{���V�I��I��4��L���oP���~�Ik�r���k�e7_�������c�*�q��{�
� �����,^��������ټ�11��񒀰#�z�C���?1q�tv`}���u	��@�[����}�:�q�V�e���;A��n�NzHdZ���X���[��N�@�7���z�ܓ����٥.����-����������k1�\���.�DJ.�U;�豚��8	\���d���XXS��4�_��MV'7�iڅ7x78
���)4�4/u�_�v�M��p0yf9@cA̐fVM`�J��zt�y�h��1���QIwqf����P�e�|AX۽��:-��%��@�#�=�]0^4�-Rp���� -"az.�8<���e)g	< A8zɧ�]�벶��%x/i]��q�Tf���9��u\���s>���N9*����|w~-���8:-i�#�ٶ<�d:�vR[�G�d��a�6X���}��v���c�����ٿ�-���>x�}V_lZ{��$R�Ӱ5l�ַXO�4 �-�\é��)�\���� ���d�<"���Ɓ{��e��wx1���b�fY�� fm;/"]�U��4lI	w��4F<??��S��6<.�=���99%0b���t������>��r/�g�����KW���k�7��y �FCU�`����z�F�u�v+�����a'H��#��$hH>��Ot `� ��aP&���l��� ��=�+��+��6kb��{KWL�Ǎ�D4o����yJ�*�8�X��T)�y��l2�΀V�g?�/m�&8s�N~��M����}���\b?��7�_���-� %�&��Y���*U.�]iRR�e�AQ,�|���'��(-؝��a��OX�[^#��iv�CN���(F��O�-(�#��� �q�1T��|��x�G��@K�{(Ћ���窪U�B՗O�8=�xK.�P������i�fEZ�g�%K��4)
���@zF��x��S�E]j������ϭ�?�y2"�DF0�9{a�VF���c��l�]�-o���I�̈́�z��S�-��Mr�v޳0��}�a���-��%�&-&l�`vS{�fj'��mf����/��j;84k��Q�s;7���s6�O�l��^y��S�޳k�����+��W��E��Ga��u���{�>qs�}�6�U���v5[,��@r�~���#��.�NO����r�b�j�$�XC�T�"kU2���4T��7��Ti7����MIƍ��v��=�����+w��k����ì�����䩹�I5A�Yc����C�k��j�֢�$K��4��,U�R��[�=�ѱ���N�A�\`scm,�&�-�q�m��4���� # ��+�&&V���e��+�����'���C	,�i��k�όk�Yh���I�|�L�9�a5>�D�Z΋�K��]^0'��ka	�0�\P��E���S�˯W��|{�c���E�ѯ��4r�o11�sV���̫`�{��@�/��8tx�	G:)����9aէ0������E��G��Jo#0�!u��`����׊�c�h'��/�֚��z�)[z�ꋮ���o����
<���a[l!�%IK�|3Y�Q+mn��Xl��6�/�7͹8���M�C2��ոO�Jl�*]�Ņ���/�I6E ,�a�̸�u�(����q`�,�r�8���ͦa��$��f���П��`���*�"��8�ӿ+��2�
 �}D@L��X���u��;k���Rբ-��/��r�s���ܾ��6�GՈ�6N�L_��-�juk��tFi�<��u�bn��l�*8hC� �( V��%~��+%�,�����$�Sb҉aF �ҭk�0T�z�8��� ��9�AJU�>?��_�����?������'��۾l|�K����F�ۨ�C�]�nAY�j�,�T�JK��1ǯu��;@
�7>I;�!{��iۻ}��dA����I��/���!�6I9�:3h���V:��t��jGW���}�G��+=��Q�YJ]� �%��fEշ��Y?t)n0v�Zid��
�I'ɃҋF�\�ϴ�Ybs����И}��>�$l4ǭ����I��u��{��NU�RDXz�g�p��t70���@�ⴶ( �5�����:��Z3��+a[�aQ~� �挭Gj��Y�,(*�3C"[F:�0�k�����ŵh��U1�mI���Tg!su��i��S�����:�����G+S��t��
+$�m��f��m���7?p�н{.�o�@m�>^4�Ġ���ԍ#���T6���+����659h��i��w�ho�b�Fp�X�B
LN~ҋ5�p��%�t��K"s��`�Ӽڼi'�Ő �E��\�YPx�~����&�[�z��'-��j�ڶ"�ﰱ�_@��J�b5\Z�A�T�;�;�s<61�T�0�ɝ��C�S�B$��]�����mq
�;F�ҙ�6���@�6'\��a,���%6pEHR�RKڞ�J)�: +`N�j�4v� ,��h̷�<���-����۽Kx?=O� :>f�����y���/͜gy����|�s����Jt��Ҵ��	_�Ŋ1Y)�U?�t�:���ZT]=��8�R���V[�z˰��]qd�������u;:�<:m���?kɞ$ҁ������������A۳�ͤ�𞘰��]��'�6�\��.���.�e'����:>?����4��y�H��2�r0:�0�&�'&g�P�:z�n�ta��Y4I�c���la����н� 	�e^�|��.�C?�=�/d.����q�=�h�{��v�Aڰ�O��Nf���h���h�K��!�owc��X-�b��w�L�Bh���_"��g��(���;���f��F�(~) &�� �XJ�g���x*�̀��oH��?������n�����#�O��?B����e�Z��&�'��飏[P�)�	����&�q��ڭ�M�:����l�.���FF�̝���Xw�FC�85��A�r`���?�3� �vu�'�Cc���Ͼ���C"`V��c�=��"�=��}��i�5&��*`o���{���#�;cW*7�%��;��<��D;spKq˺���L[mF2���
��J���m��v���T�NO��Q�.�����(�Ybt�vl�l;;����Ha��6<��#����uJ�Wg�W6�&�a*A�u戻��3�,Ud�'ӫ+qQ�iXe�]�g��'��ѻ��v_���kv�?y�(�6�m�e�1 l(6cW@��=C�)tpe��N&���rAs���b�v����^n�m�F�8l1vf�L�@0��� 6�C �q�ĂT.K߮(�{*Qt�ʁ��e���A(�n9��$ϢosC���}�͝���?b;��J���i��?�)���/Eh�n�G�5.{ �2˨���ҋ���br���Un��҈,F���z|7<=2b=hI�\g�`=����a+��5e*��o
�҇�׬���q`�Ұ����i�hã#�m}��<6e
-�.Z���j��8T���D���E�2~���΍@$��E�}�rvl	�sZ��e6F���O��'�SS����т|�v�}��o�x�)�"`XY��ӶHzd���ޛ���z��wN�����E�h#��B�K���,S`	 ��9�渪ռ�R�Zq+`,˼�����Yi1��}���`�&`c� i��}��SŘ����K�Z �`���QV��+8���K�Ͼ�Q�+��^E��� ���o+a?ÊƄk5��[�����81� ���/��>Ue(L� � �t��f�;���j�h�x*�P!�!=��� Æ��Ul�5���+�(��;}z�«y$'���Qv�.����>e���u���~����rl���I� �Fg���&��=:��0f�H��sg���.�w��56��<����T���6|�(�Ț�^A�;��-b�1�N�Uv��)��)nUI�	�g yn��@+�NNz����]������P�/���H�M@�cb̦��a#���s�6�(��t�^�>R����C�޻�Tz����h�Rd)td;�@^{6}�1�1 >*s7)����IkM��;�Zg�)����ؘ����])Hz��$i�!�
�"ѹ�b�9�Hg{:��]�e2!�R�&���z�ҋ}gw*�͕�=��u��aڄm��h�mvjh�����l��i����3,�	P�-�],�����e�E9|h���x�LwVf�n}ն�T�����0i[����k�c<�u��~P�^�ׅ ���F�oob�Y���K^<jN$͍Ojsϙ���@!�4���OB�Vn�S�'ܶ�O��Z�R��;�]t�^|L�6��
 �������5F����z�8�����p{op/��+��w��-�Lr�����d Pu�<��@���+1���v��i{�}�w��,Y�+%��<x��&O��K&A�~G������)��|��`ǐ��
�ܵˁ���d'����q��rFBm1e\�����>+A-���<�/��+��j����Y�|�}���H f9������K�,���u�03I������7���z�G�+�݅�%�ױX��򜁝[캋_�:m'єm�������d�������q���:9ȫ�&X�M�~����Z�<��.z �-�nQ�/���v,��������1bP��ӬM��ټ�>i���M�l>�M)v.��k���Z��l�1y���ͪ���M0�{68�*��d��)�*�$�i�w�Tr�ʶ-��,�s�M���p7�:]�y!@���`]'�B���*�A	�I�k��E����R���b��`]J��17~����au~�7�=q�d�������m]���?� i���X�L�&�b���l�`�f
1;x��n����~��v���w܀�mʆ�9�!�Ե���1���c���cSV`fIbdanJdL *���|W�Ȼ+`���J�`nD�u��ױy���*��mӵ�]
~ƞ�T{�ٲR���lq��R��u��O7<�۴,����8���*j����{ׇ���4�� Ș��ȃz[�Ҷ;?K�z�݃y�v���sh����m��Dz~�R?B���;��ܽi]����m3����z�_^��J������87y���Юx��3W.�o�&Z6�f(��U�V~^H�b�Q{��k���y;D����Ik��WN-V�}�F�R���x� ��+Sl$����;��ۄ���{7؛X���U�+s0�3�T���hox�m�K3e�ڭI�	���c"�?P{`�WQ���Y�Ey�����S��}뮶�[.�o�y��F��:�vZ�Q�6�ދ�4B���4U�{*x��	p͌?��4�/������2�L2>�z��o}��8r�6�뷏����n�;gH ��T�=� ,�Z���&}�tc���Q�@��u����u!�m�Xo��p��s�m���8�����~�gPSb�ଞ��G+�xUw�y��߿�~��'��u����;;+BZ�U� �)��.VF�΢P!�4�����_a׾�F;F���߇Їl�]�c�	�D��aS�m�t��˰{�����٧p�&e�K�(��=!��L=�Ar��S���9	�éү��&�Yx0��TY����'��H:\���[����,~�C60��v\t�}��� .,Z�Hx/wEW��{Y��%���3 ���E��l�)�|���Ҧ) ��	��'�	 KQD����-8X�+��ť۷�6l���4h���yW�zG��sO! !U�� ��M���pҠj*�jc@%@@ `�k��Ha4߀}�[w��u�����llj��!e_��v���K��o�m_�����Ƌ�پK�b��Z���m�nǇ�DKh�ߝ��2�;��ݡ��X�"�I4���"iɲ!�F_�T�ړh�Rt�����a�E��ɵP�]��5В�=S� �hc��~�(�`����d�V8��O��yգ��!ʤ�y��s_�R�s�S��Fs#���@�P���e��0y>3ՄW6�\���v��=:�t�L�c�vP��ל�omX'U�pjӓ�����C��>ٻ����6l;���3�k��,mHq���F��ii���_w{�m�46|�O�:��;7����(�� jggG��C�Z�o�U�f�G^������ǎXۺ}6˜�)a�Z��d?^4�2�z��P�c�Lآ]���^��J��)f�Y@�CGOx�ʺ=�Jt�ր1ɱ��`"��v2����uu�
EZ&�Jՙ1��rq�󤪒�:�UU�H_���T�m@H� ~�ν֕���?|�F+
n���/]ʕ��w�p�S
^�`u�Q`+]�d���5�R�i(�!��������g.�k�#�������tZ�2�ڇ��4��e.-���������������yAee X"�C�Y�z((L�P�O��D�`�E\�[��%E`��������|֮��*۷�R������kL�K9���:�t~i��8,,���؁��A۹i��u��6�8��~	���v�5f���?���h}���NqO������}Ǖv��S6�+�}=�{�Wx��+E�6��+;@�8�� ��B�jJ���3�S/n���]lB��F����niV�Cs�d(Y-��6����T�Ν;4�ݶ*�!����M�~��br���ї��#LQ���d��@o�.�����R�Ki�X���ZvPT0?�s���.�B҇16R�[�w[�}+�LR��@� />%ӳ�����r�5��a(���p���f��r��g��[%V'�
W��e%�קh>}�c��	���K��q�`w}�^;��!�Es���e#���S��g�v�[�Aŷ��f�Y�� {�[���C۴�3|�˕�fM�H���j�h씚�@�X@_��&!h���h��>~�7��w�n�8��SI:�j����2&0��S����j	�120t�Z�m�UHc�4�6dA�.���@�~�wsm1������..�4A.Gqv���(m�u�W� 9�R����u��&� JZ�Ә���bs"6���4:���B��M��u�k�~��?|�BS:��]�ST���鹓7�颫'�mǎy�C���},*��
vT�r�����p���}��fCΞ8�' Y
Ĳ�:Ƞ����鏗���N��a���c�F&]id�Y�L�M�����Q;cx��`�Z@�����D4O�8U�a(���M;�-T#�:������	!�Q�B�lVJx�{R�����,RyQ�&[+���+�H�v7��{��^	)`�JN��րq���%ӼU�
2]l��v���tw�8@�N/�����YZ�y�$ƨ.���E��H�%͈hU���O�+��� �I�4P��~S��]O ��Փ�Ư.��e�,Y̘�NL���!E�N��HkȧȘ13�-O0�ͅ_��w|V���tS ��j]ŵ�>��e�&��##g�-�_n��g�kg�:i����.��
�����o����
㓶k�evx��v��M��w^nS��6?5l,�	��a�b)�����	 O�t
*���S�{���8�Q���f/��;�utѥ��K�کx���V��Y���]��E+a_�ۿ����,쁳��,��PZ�_�F��Wg_��t�˳nD��:���_U�`�ĕ�����GJml汩P �ڸ��HC. �[ �*�Ѫ�~��{N~S*�q#P1.*�;`.���X1�-��S���FLU~���:ڑ�P4>�F�����\��#�) GU�īN�~g�'��PE/:���7�M'���>E��������=z�Q���>o�������Πm}J�$��	� .6)�����$I�yAP��@���[:`��O�t���]6>>n'O��.w��HU����.+���w��B�ϞzQ�V L�2Ǣ�J��sP*bP�T���wN��t����6��c��Q{�����3�5����b��Ȍm�S� �L ���g\���9��`9��=�F��3A!W˒љ�������Ow��/�ֿ����h��C��~�H[���u�6�:pϷ~�83|�����Q�a6F���oޮ��C���v{pbֶC�W�O���<��x<�E��&F\1��)�Rn@aͶuvՎ>+�<aٶ9��MXW�i�<C9<2M���;.!hSq����15�z��Z�=�� ��yzOOR\a��nÐ�r�S�q�.�n��(7��	���"�ZI>Tq��P�a�����;Y�[ֈ�
��yQ��7-�̂��6��pZ;"���b~�Nnz	O[��?���'��.޵���	��JE��fm�mv�= ���uW^�(W|�TգpjF�oëU���E���D�i�ܵC�����{/񳪢T'CMi-�3�;R���T�4Hҽ�[!y.[�j��/�q_�)��}ٻ�ɹ']���!�T�	�h�����8x���?�E���v����~���*�)�"�N��wݏ��0E���#���/����<4-	7]e� |��H����J�+�i<=��C�::���h�n�4��Z��(�Ҵ�Q��EW\i�l�iT�'����yQ"���� Z���#z�Rbd���<��z��0%A&(��ڸ�'r���y;~�t�[�PI.s\�����h�%m��~��܋��y��)��4lR��j���D��x��`t6㺄��$���4Ϝ����$w=`��CR0z��%C�ɪ�K�]�����a���;�p\`�6ı(�VA��`~MpM���O¸^uݵT�a�S�3ڨ�؟ܷ��-�����Ω�B�XJ�%p���^�
�=t��XM	�U���掝;���ڭ_�6�v�kv�k�����5P����P0�X� )F���xD)��Z�Qt�\��G1L�$z�*�F^Re|�Bh� R����r��3��>�0�o��ZR��s�L�IY�tv���V{�����9��#�ѷ3O+��.����$s��P\�Y�Y;Y��������k/��o���]_���y�h�l����C?u2��Ҽ��?v�7��6��r�ց�"�es�N��")�=��y��r�{��[Y�z鱞x_�U�xQ �yGw_jY,57BafA�7`Țm�6(FeN���N�<�<����1w�u�mBHȎ7�A�PQ�Ґ	���Y�=�x�c�Rۋ`��΀�5�ze�:@~�I[�ẝ��(A׎����M���&h��ޫ��_`+ ��"��g,	�v�	.���ts�����T0��듇�?����������cv��o�i�<��Mz�%s������ԗ�E�*��E>c���u�Q�RԽ��JM����V �ݨv��tJ�d�Ǐ���YS?7�PG���	@t��ޫ������t+�-�3��O��������_�B�����q�� ��w�c��o����G�f�-^�4D��i�Q�]�u;����<e���ztHDW��Lh�x�(7n�Cw x^�<S�;LK�˟ˋ�X!Ff�y�mYRl%<̔:K�ɜ\�B%�����<`���6a�GF���k��_��u�7��w�= S����d�����C�1朔䋻l�}u$��i�	o`�=�K���[�����o�n?�S?em����(�'.&��d�3x�4�5�)����,�#��j�h� �{i�Y���Ő��R�#�6�x��]��Q{�A@D+)be�Q��(.���)6���n���a��R5��X���dڏ�ȏ�?�������������iKo�k]�lVv"�KV���!̖�ǢWDz��^��:���	���?��-��~�~�#A�Ά@,��+1���������i)�@�w�Vp���=�i�PB��J��HN��N)� LzFܾ���w��>�����Y�FA�T�s���I6�y�^�q#�Aa��60��œcnl� 9�ߋn�Lm�T����xk�Z6?�q���o��� �hG��.�@}����3��]r�M_�<�3zztG?����u,@�Gۺ���^2X�c3�؎q���f����@X�V����zbv2��)� ��{i]#�R�ʮ��M���+P�'غ�R�IG�ٍ���?�qn��y��/�kP��븂�t_U���<���sq/9N���LV,+h1
�3��R���vUAPў/��Ip���A�"/6` �����[_�"v=p�����>�$�9��0ڇ�}�aRYE�0 +�O�_�Bb�l��)�:p��O�Kv��e��J;C1p�%J�  ��y����s �+��]|����JДV������芮Lɬ�������r���sAn�����'+�k�u.�6�}ى>�s��<ړE�ɏ~��684i��`s�kjse�9��
8
f1Ɯ$E��T���dY�*,4�nH����t�1��=.6#̏	j~K�ߊޫ&�,7~<�Js�;��*��t�1Q�g&XYG-�s0F[�m����(�˩s�
T}��	�P�˟9��׹�}v�~z��n��3�#�g���I�4�}H �%��dW,�,��<���D�� �B�/ 	@�*م\Ч2����v��I��̙U�,r�+9��(5u�}���[��N��۶�[�}<S}(7��qF:��w�l����G?h��1k���B��
`���B��Q�ta�Nc�Z�l��ՙ���'����4`Q��!�=+��88Cl�'9=3��d�n.2�t�˝)��ʥq�g�e�~(�_Q��r�W�Ӿ28X�̑e�[�2��K�k��7���I� �&0+=������q��W}M��l�7��B�Q3���L��|�+�Dv�+n�\��+�����u���<�ؗO�n��U ���OljiG��`t�sq<3��w�.�|ۀ�}�D5�%%Zz�?^K�3�E�\K�+'�\�{�$��)GJ��Un�h�.f��цmd��r�%�Щ�1U;�@T��P���_��z��w'�y���q�,�G|�"t:څf�E���� Pkm���%�x�^Р�<X�����&���6v�J)��S�BU�I���6�Z����.
�� g�A?t�C��NE���,�*�v�>	[QN������,�A(��T�|�sS`Jw��'	��V�k�O�>8�
�v	MeU��V�$g?�ґ�>���)�.���E�%J�d]�b�t^��r�H.R�����T �u�-��j���?�+���Š���66�Fk}�i��w�{v#M���k�˵֩�� �y��d�T�:%�|�;P0�x!�V�{�/7�T5 @`�� Y ��}`�mصϚ�BP�C:��{zz-�i[�cV����Hѱ��Mi&9�k��c���	��H���mޗؒ0�,������i�A�ĩ�v
�g���!i<�m����3�LMچ���;� ��",B������Y6��1G�Rp�:P��ݟR�٠��,����`Ǥ!U��Zi��^��~��ٶm��	�z��O��}��/c��;v��8
���1��In�vo�>���hM�G�����������؎NF;=+R�휢*rt���kM�E�sUi�|���І9���0���P�]UKVd&�e���̹NA�H��H���YM�`m<*/�O �V�GK�%�5!TYx��ñ �f(� ���5d�B�r�(0���\�xH��HbɤN��(lT�����.��e�aª����Y����tѦ
�X"�Z̶�mܾ�d�u�Kf��wٻ��|i�g`�c����S�����ʤ��h;����[�������B5��U�xQ �%����.v���T:�Ksζ�aA�i� +��Zb?�+���fs����K�!�m����=�A(�t��� ����՘T�uX���3�2Ŭ�c�J���k�
�	�J�k��Nai�����n2_,�����3�W�)%�O�ӋP�V���<�=�IS����0��$�(���"7u����i�깞�tF�C�W���^� SzD� ���*0i�H�������T�)}AB�4�\�s���J��"�b���k��ct%�ذg��Ѯ��ό�<O�k�5�R`�g�+ձHZQ�fC�\wb'm<I
������o�Ύ;f�6���~����~�n��#�ӂ(�U�`.��4g޽�fǋ6�&�XR�,*j}j�M�I��x6��e��>_�HP�R���^�S�o!��/҄=v�1�OCv�u�696e�X h�ڼf�����}�_��	6(��H6Pa��I�.�y\��@+�nɸ�ٯ�yF�;7%/�Z�bv�>v��`C���˿����~��C�۰�PU];�ɩ�O�&���5���2$UZX�b�J�e����Ĝxxw&L�GY��"�g�hy�C�U*�y{��\/1\mu�lR�?��߷�����:������q�v�7o�ߪi?��w�T������O����Iw�����7�F��(&j�٤J�L�q�^�G�8f{1�ڴ�v?Ka�2�}5X '@ؿ)�ϊGb���K
�����h���^����5XUŢ�>�:����8hj�������@�	|���S����>T}Kq�;����}�<���)V�G+�DU<�if�Đ���+/�UUd��	yCjq�/[�B�ʕ���};�G�g/j���'�~Ѷ�q��U�/H�Ls��d6q����S����G�9�^H���q����䚍��f���f�?^c#�\��S�D�d�7wR�>����WZޙ4�2��L���0}��I7`*C��*)�PW�@s�-����O0���S�F�DQȌ�Ȥ�����r!�)}O��뤜��9Ⱥ!Ji���lĵ��i�Y�k��><P�\���i��zJSW�*a��nJN�b�<$[�`š�{��m��0�'(h�����b�H�Y�#���cռ�cɪa-LZ]U0|o%`���qcF��
 gP�	;X��Iz	��*(h�y^1)��&��Qpo����Li��xݟ�9=[�B9�=W�i$2�ec�4�7��� _�,*-�m��}+%�\ϱ�Ql"��������>�X��Ԙ65��]}�6K�יqv����p�˲�q�\�4�JfAs< �?��%�0�ʴ�:J"F��G�}��g?6t4�!Y�������}61;n�1����{��T�QE(��ԊޝB��1�22b��=��F�z��e ���Yk��p�4�pSޅ>���cT�aE#G|4_S\�\F����]�t��"f���޸qӒ��i-ñ�����
o��uo�Ƙ��G���3����)�m�=�����X3 ���9~�~�W���"5����0@�`KPL�����:����a���׾�t�$�� 	��Z1�LR|:|���8��v�*�q̢���c���Zֽ��*�^�Y��X����]]�}�A� K�����J��}�"=�)�&�ޠ;��X`�����WF`>JT*�b탱l�c+�ʏ�7<���t{U�Ĳ:8��e�}�T��["#MҰ*NЭ�1���'y�}�"��=[�K�	�y�
�J��r��lY�s��̀���l[�B�B��d|2��֬eZ�_����A�Y{���@w[�PZ���{�+@j��њ�o,�IP�eq�ס�h��(�@��/'��Ï���6���A(�
�47iQ}$D��\��_���/�7[P�ЩUZ%%�F���,�+�l��4h��y�f��$=�X�Eˮz�O�Z�ɭ��f�+G�!7o� [l�3�)����C=o h9 n+�άu�\YϑƔi�v�������U �������#��KI�2�`G�]��ΊV�3r|&@�W]^z3����R��xV�ɯi��l ����=S+G�ґ�Y{�g�-�t�cy �	�R�b���c��؛E����kJ��v���-����Q]�Q����TD��e�n��?j���׬c�$,�(��ӧ�m#i��m�G���C8��w��L�y�Z�?�o�'gQ�2: ��ԩ�/���a5�W�����0
0�G+�ۙ��i��GK�kΜ�fϩ>L�3�af���*:g/�N 8J�9�"=�k*��� +T�y�:lj��ƥ���� �cG�0�	�Mcrb���ea���&R�^U��9[������ݳ��ܐ�����sfR�F-��;��s�	�����GR���tYti��F����,<qP��Y{Wͳ�����>����?������F��8�2Qs��b � ?Ata��b��C���o�g;��@�Rp�+:�|k��aє�-�{j4�(jӘ�5�"l�\��I��sTP��^=.cki�6��� �9�V�B��� s�4���<SQ�6U X����M0��(?7�w��̗ޏcѭQQ�Q�@��c4�N�K��G�����l�hu3��4+S��[Pf!8�V�,6;�r�X�pY����\[1����:CI!��>>�Y�:~��Uٝ�4��j���(��q�9�O%�WS�X5>@��T�	\��Ŝ�Bz)�C_�ۘ���QŘVI1���)�"q��z��	�R,���H�L���2j�Шl�NөQzK�"U��c˪��t����4�Iwa'�JQ�3�h��0����klh�TW1�e��K6K�IC�a��5�
B�E"S�h#B.�XCg-�N�nv�-XTd�I+K���f��Պ���n�e_��խ�t��@����@<�4p�͜���!K��)� �R����u~���h�ݧ�,rx���sFO����(�!hJ�*������ ��J1���e��,�禲Z)��Ѽ�w���>��V}m���8�՗������ظU��qt)�T�Γ�N�a����:�*��N����G�m'��������_��Q �8�2ٝ�ǟ�����5n��'()�~E�殔
	6v�PO��d���BsC�����$2gƳتt�Y��R�bt�,V%��D��T��Zle� �����QB>Q���'*4fب���}y��孿},Z7�Iz��(�1�d��R�9E���7��s�@�Ͻ0�t����F�XG� �<�9�`�h����tn\��(�?)�������#I�
1y��n�w��U/FY�:O]6bb��	-�xS��[J_�)�H���PP�����
�� �|K'ڴ1;t���\��qy�Lqi�1O�-�>zu�\1;666��fF<z��3���^szªOaT*�1� ���J��L��O�,�@�폞����;��G���z�X �ʹ��,�~�J9ֹf%�N���wXPzV3� �S/ͫ��?��m#~.G�u��*Ƨ5�^mbu�U��-�����GƘ�Vk��
EXS�0�U	�pƘ�u�z� ����(NJށ�R;�� `��q��܏��O�.�X�k\�,s �/+�ױ�!��_��oE �%�s��Y�,Ȃ2$9i$�"�/�#�wM��O��%h���ʐV1���`H�tl��t����ƪ�V��t$�h=V/&H���L0%���v)�J��8�j�1�*�*a�u�6du�>;a�1\�o���9P{{j��5_P�s����K�^�xT��fT�����tx�/�b���jǦ�$�aT�k�pN,7���2��s���]��R=9�D1��Y����ևE*���g&��gIM�)cy�B� ��%[�����>����A��_����[���p�k[6�ӳ��
tDE�����qi�J�l�t,� �]ū����#j�|'n������Z�UV�f����w(`n%��@\�7�_g��s?g�<9L��שP�/G�c獞������v�������n���3�q4��wm�/|��GE�����;O�Sv%�n��
�uYC�7)i#y�����s	�x:\����P�kb'>�*�WjI$F�E �f5�&���VS�=�/�ʦ 1�mX)�*���2)��������j�^�ez��qϠڴq;X���A�V���oR�n����q׷	�G_���`��@&0K{&�uI�଴@�3]\��e����wIA<NOv�д��l��/��w�yX�:�j��#5В,�x� #�}h�>�w�����6�\�S�~��_w�5̕>��]�ѩ�S^ء���m]�V�D��Qjݶ~�v����v���k���~��?3��-��yR�b��Ӈ�l^Uv(�,��6
�a��4����D?9���	�+IW�j( �w^Rc¼��B/n�à�/Qթ_	����W�4y]hrs��2�H��7?w�,X��\��3S1R�@�a6��>�ז�.� j핡9�!���-A?�M�d��@G�Ldc�z\��٧�xF����w|a��P��B*{.3�4�0�9�~g�F��Vk��/�S_�/yQ 2�N�wZ�+���<����2jpé�C �&g�M~,j]�����%����gM�`au�;;�"��*0��`��>S5u	 �Z���I�'o�6
���C4͕��{kQ"��e-��X7��F�.����TU�)S�%	���j�b�w����m?���Tor��2�JY?�U��e���p@�� gӈ+�v)��fe��v[SP�s��Zl��Q7L�LZ
�e��>s�>Uՙr��v�s��ɣ4A��B��|=_�s�0p����M�y�*�s��H�nْhi�\����R,��:q��*a�{��؝��o���]��2�C�ɐ���)�ld���{���M���>�)�؂m�o�-�;���|��:�R����W,�^�D^��N�S�Ԛ�X����Q��eWbй��Gyf(� �<��un� =�661#��.JӞO��|�%z���Ξ.��fBZ8��z(����K��ܮ�[w�g �UVAf��&q@i6��bC&_*i�CZ�pW�qgg��@�|!6�(*�J�$`�4��QI�4�Q2vָK,��0IC�G���3=��ʗ��*���#5���w�4P;�쳭��v�=����f�B����l�Mh��z���g������o�o�v��s�>�b�%���D:��#�7/��U␀���@�:(����n��F'�BL�ȯ�ۑ�(�^\*b)E�̈́�]�}[G�8U:*晇Iҩ��jc�=$��2'F�yF1~d,R7�#���WQ��	�tæ�ؐ�<t�~�[�{Iw����1V$K�����2�^,U��ǲ�ex0��B��Rӱ
h#�E  �K�gP��{��U�_㾍Ad�x\}����v.���,9�B+�vD5��&7�RB��j"�7��]�*k��'� ��<z_w	�$2c����@�<ǪJ����]��tK����K�6)n$��4������@)������yiq����q�X�E��7QM7ڌD�զ(��k�&Q����f�^c\��ܔ;_�ʌ���P�������6۽����;IsL#
�X[�J�/#Y9f�1�ǝ����9�5�]���M�R!|�4�?������w�Ԃ�ֻ/(�� /�a�:d�������*�g1UJH���0.��,~ێ�7�x _%ᤜ��n��,��~~��}�H���'?�7��+vۏ�л��K�q��Nt�x�E�e@�:��	[����vl ���PJ�}�*�{
Ff۶�P>�q���Zl��o������z�.1DbcC��g� �Y,8-�6WW\q:��l�:�9�߰P�B<`���sd�	�ߕt��\n��<� ��4-e��~k�^x#���p����� ��Q�!-�J�i>�3��>���R� �4]�F��Y��E�D� iV�{(7{�ғta|���������7tۆ�8���s�� �y�ZO�4v#�-
��.�a�K��ti�s�1��\�^���A*����"%�ALR;8�E5� Rё�u~�x^�f.��B���c3��lR���*�,�}�*e!�ƽ���8��s��\��1��.C�ՙ��F֬�%|�Zi1Ձs~�ۃ�`�ڨ>ªe�������*�r�7�:'�I9�, 3! �!c�F#;;W��A�, L)\e�[������Y)1O��ֵnB��j�����4)�U�t�}Q ��Q"]NfڪsT�hw٪�/ˁ:���ė\���HhӃ7�W�8��	��&�2��;{��3<�`nb*�P�\"~�+��$g���Հ�Z�^�^,��yK�����]�(m̤�`�W� ��8�1�����%�{���Rf�\�B���X��p��_���T���[l��A��&i�k�2UqM������ZZ�b��.�7�fJpI��A���5-���Ot��i�4fA�@�1�p9��NCSCU�b��j �}*������P���㙗��҅�.~��AA�rF���V�/�	�%hZ�Βݾ��>�\H�Y�I*�׳��H�m޾�S}�C�l ֱIn��C���(0�d��h�������-r�ؽ'�)��ZZ���q��L�rd�!"aޙAƛ��M�|n�8�V���n7N$!U#���`��3ԉ�������! �]K��p��s�.^�s>�4�*ι����Dgw�?�������>/��f�CUu\rU�js��Oߺ0�t�5 Hw��Q{��âk ��`�,��5����Oym&�1��S���W��_ !����T7
�LQ��F�- ���:HUE���f[�lG(�h��[����u�[�y�!��ڼi ��8���B���t镗�� �iR������LTo��*���"��4Ũ�I��ܚ��V�p������^</�O�������`y��a�`��?W�Y�f�kK��E�d����}\f�hq; �6X�����r��~�=��P?]���X4�ҡUYݛ�Ul!�+i�۝�3d1*������k\[��It`q��iέ��]�T�3��*��<~t,�w�Kڴ�Y,f��~`a.�u��g���Ǝh�F��>shb�ߚF˹�W���Eur��|{ubv�S�F�1��	,���؍y酜r��y�  �J�W�o�,E��]X��M.0�tdP1T��wZ���R" ez;׈qqS��%�(���p���A�9�9�&����0�B����}���R�Z$��Ƕ�@1_�&��qn޺;Zm�@��x���Vf�ͯ��r���Wo��N"��b�����H͠5S��
��aD����_�Μ�V�[�y��E��b=�fةj7t6P)HIF���R,r4��A��(<�����
�Lg.��� S�~/B�B&�]TJ;8
(_�nט�247S�ǭ0y���|��?򑟥�1o�#���d�l���* �0ԁ3���,�����T�.���կ������S�|yE�c�o�ߞo0"&L� _Tx#V��ƶ����g��-� �0so�Y�tv��b:E����_�����6���<�����:#��3���L�٘�#�?��a6�#خ�{�����ϓr;��⚦̶ZJ����j��-�nŸV�v=T�*}� ����Z(Ȳ!��[9W"n,h��ۑK��E�P�cMV3>�X0���E�T���:��M��7\��{`���^��8+n���V����D�"5+&Jn���5#���" ��~�~����a�:�ݻ7���ת�:~�u^�bҔ�5�I���&A|t���ɪ"��`��V`�t�b����g�U<�����O}��a���o~�}����B}��5bcB=%k1oY��4�mn�bߺ��v��YoO��p�o����N���F	��T�`�IZ��P(/�4Ǧc<)pm�vs������q(�L'�Ʋh�vp�e'@��`_@ֽ�`�����m�:szo��]'y��K|'����Wf��H�+�sXV��˅-I6 �N��������>��/�R��K�>/
������T�2H�ع2�JP��T3Lp���	^�<��7��/���Z"#B�j?��#Pv��p�d�?W��I�AJq�����7�p�C�����\7([9��d�/ɸ����G�5a��Mz������axZ%oB�24�
 �*�Nc��4S\��:	n�VE���p�P����6�n���;�ŰC��;U�3!��"� =������]Ə�x-X���\���I[�گ��7i]G�ࢋv�s� �L9��q
�
R��p���v����7Ζ�_e�:w���b�t���l�уy&@�`z�LXtda�-�q��0r�:�{�{��^s�5���}��oٕW_��73Op�����u�� }�fY4�)�Bxm'Z%~�l^K�X�t�F�0 D�b��<F��g���U���	0	�w`��K�n�f���?��o�jbjw��g�4y
MNg� z�d���Q�O,�4Kz_=�Jx
Ӟ�ы�&���/Hv��m;vl�/{�A���|�co�\�*���I��~���[7@��6j�ݳ�������IG�ꧩ_k�1�.+ 6kV��c	��]�P���3g�kH�����V�j�#�Bk�Zb�v�vsM�a����\:`�����Do�3 ��o���|j���o��s�NA8�n�Y|ɤ�V�U�ʜUw��$���	g�Ka@	-���߿���X�b1G��4�Kl0O?c[�nu}�<U�J��R��L�b�#$vV�aa�׉��|��:Yy��>�����#���q��S� ���������7�UW]	��)-Մ��f�y)��[�yE�b%�Sf�"9Y���G���X�^@�Z� osb��RcMOM��:qMw��������Х�cC�[r����"�\���Z��&�6DQO)���&��@xu?^SW��l,�YK��ۣG�l�U{Ѫ����U]��  e���T�e��o	��{�EX;�8���u�ܹ篹��9|RJ�xL�v�<e��(��R��t+Pó�PSп�2�vv+-)V��:7�t_�	3P�J!i��<���H�]�
ŽH �Se����)J�y�zI*EX�0���O��=u��+��.1��z��l�NR9l�tcg.+�J(*����V�T��{~9�{.��Twg�.��=(W\� �.�o\d5�
iW������������<c����
�
B]�]4\�w��>������3�m�l��k����i�Њ*�eլ��Γz��׫���p�y6e[6�#u�j/t�0/ӓ�Ss�qR\̑ǟ|��_��-��R*׼�5 �i1���9[��$JE)-]i���f�A���Y�%[�0�������+xM%�+�nH7�E��IP)����]o�Ԑ��SW5o�9����//
�Y�u�?߼z陮�S��}����U�){�Ji~�"}c���9�2cĵ�I���K��a�
t�$1b5�/0�̣��QemT�!m���<J�y�M~VH$L����s���v �s�5{��wTy)��
�
AW��Ȭ��)M�/R`R�`�>iMi�8���D|�����[�BK*����N��׿���:겟��`]�]�;0ZҨ)[@��656�y��<�w7�,C��|�q���oZ��=�"v����q�Ӹ�K1�]��"t3��+b@�>��iv�U�6�Y��@����<{�	�Q���O����T����fk�
P5���T�N61���k��|��s�-�d+@Z���u�f��L�Sg����Yy�-�k@�{p�Z���~힘���o�S����/ڸ�>y4S�8���#���Z8�y��H�V]�'%^�=�,�I��b�-]�eȉ�ґϴhit���$.�[m��Q{�e�#��'�2�A��$HW���X�yjslȲ}"��4��Φx�� ��*�[��Բ���
"�27o���!�م9���	�Z1�)8���+#=F�ͨ�r%3�,��W�"�q����>bܤ
ʢ؇��l��Z��A�F,0�de[}>C��j��Н���]��7��Ӻ_��6���G���bRJ��������#(��N� wߞ~k���*�fp�^`wM���N�`�k_f��;�pٗ�U;Z19v�I�������N���	�hy5�m�� �޺���/p"���1��*�$HF��|�т~d���0c��y����E�g��[�t̻vL�Q�״�S��P���˶@�e�kp����+�N�P:穨��CT��C-���?.G@,�C�o�������ao%�Vi�&�jzȩ B,������@�_	�-�����3^�`���=�P�Aj-pd'����?f佦����;���r˯�:U(e�"��9�h~T�'���N�3`�V�	[q����5���O� mj�k� �6��VZ�&���ڨ��`�n�Ң�>�f��+�x ��2���ٌ��_~��Qˡ�z�Wm߾}�ۿ���$ͷe�*(���}��*g�\�,)G+��9"@�tc�m�$z�ёQ�dߥ^�q��Sv�%��<�لl���OM�u���ZU��I���*O�q+i�	#��}�GZêC�X�{���؈�o��i��M��+�*���]����K�x��Ҹeyқ�Eҷɔ�"������_�U��Bj�j�c(�X'{���S��3Tӎ���͗�)<r�}w}�#׿���<1x2ӻ�'
������?Q��⊽[�=cC�C���:�_ �l�͎P��kKVb�TM��U�xQL��z��_�'�sͼ=E����g#w���L�4i$��Ȩ�5��8cݹ.7�KC�O7�b�DY�*�%HƵSQ���VH� S:�kg�-E|��4t�li⧠��e�8C��%S�O2��$��}��� FiH����bM@khd��/;X&p�ηR���@�Vت�����_��_�����ncC����!���������isC��c�����PY�����Utb�r}�%[[�61�i����R�<m�Wl�v�a����\ �O��V��|�	��ځ�F�bRUѥߢ���q�&Z��bE¥`�o�^�������6xc	���� Ua�S"�f���}�V�fﾽ\S�wl�X���Dx�䚍�`ˤW�����G��][����L�"�^^)$�����\�[.�V�@F<ĺ��RpB�p<�W!�xQc���ԗ��\�r�H��=�?�#����4����R6j>>�Pj�����/�Ur �|'zş�κ�Jݪ���#�x/]Z�L�"ґ�R��D�T�&�� L�'0���T�ֳ�3ތ;��N�ecS���5����e�������-���}�nz����Mg<w�n��m����І�W	���ݚK������ov�졇��{;�i�$s�V�e��񷽣˖A�+Ҥ"8��
ڮE�_UWvPU.&�Z�.��롺��������5�ϒ�DM���@�p��:a�z`����V�&眼�9�n����k�"�4��m18�A���A{�V�6�dh�hǆ
��ciq�t���R�H�i#�D��{Oo�;.���k㧆�}[VZ�=��]\Lg�3�N��������X�.I��)�f�Q6�ebA���g�vd�k��?�]�ٰ��|�Q�.H�%�?ٮG�9o���wp���@﯌���*7�n����,�
�	&�L݋XFy��잞�蠝i�7�M Ef�fY�KcxW����g)s� p���K:�iR	#�h!��a�ӌy�>I�ި�,Ɇ˘�V75����~�����p.ǥ:Ǯr�=����0;�;���������nw��E��Ҕ��/�����)�7c\r-]�ōKp��y`��Ѝ=����?vvb7Cp����.R��2�1 M�����)`K܂��H��~���&�/?�I��_�g�C�&�F��;�N���ДH�����ʟ_����s���/�-�b</ 1_T��C���[��g���!��Kl�{��hZ��]Ү��&}�o�#&�924<l�뺼:-ᛈ ,�}��P�Ҧ�<,�e�:r/|���c��^ܢ8��e����^9������L�Z��N�ۈit(�y�V��!�
�H�d�XiW�,S��B�c�f�!#���U#��x�YBr]р��uU�4L)�<�~bn��,Τ��ʙ��q�����	�*��O%֯��֭�/}��|�_��������W~Ӿ��/Ж���,Ɯ��e|r�\I^Kl�ڵ3J #��eVZt���>���ƛ�Mo��w�����l���jg�nztv �X�1?~�nz�5*�i� ���;���	Tʜ������?l߸�Kl<{�4ޢ]�?z���	ۉ�����/����dlt�(rZ������@�]���y�6��9�#����'��X���Z�"=���u��f�7[��R�4����z����m�������BjӦ��ٜ;v2־5�s{4�#���S;�[9��{6��v�2��8i���s@-һ���mأ'&m���4]?� ]ӄ=�H��uˣ;�Ɍ���l��<j�o�^&NzjKR|Mf���d����[q�*�RT�HA��ւzdҀ�ň���J��s)�d)�����O��8I�;�p*�̭��]m�h=J`�11�A�^K�6X�`7��*Ev:_Ő^����@Uau���/��Qs7�Q��5[��W�������Oُ�؏�O�����ܨ]�������,���.=�x?��҇۔�T�j�9*'1���B,mD��u���Q�J���`z���>f�[T��y�պ���/�����h��?����O���dt]�T#�ԃ���;�h�^2$]͓�%?��JaZFt�,���؁O�;��}�N<A��D���x1�b�,�*���F���;,�u�g�ۛT
����Yzz�K�M �����{s���7Jc�K��� `٪C�������
����)�+��=j�(��~ӄ�PbuBrTu�C��px��!=�鿏F=Hl�zPJS�dm������T�����)�K6�SK���,��.�,mta���-[6[o7�w��@P��${;�CU	
���*�?���g�ڟ�v�7�o~�}����F��T�!��:#++�-�\�4P�P  zu&̒4[2�.�c�N\�u��{��_땐J
]u��^-)-���\K���H�eUoJ��B1Wڜԩ���HW�}��v��{)��i�Y�wn�a{vch�a������8�~�u�O��������������{ ��<�O��M�E�Q��y@l.O[#�)GGa�`î���9 #E:�۰��=k��mN�<u��ۿ�W��kϥ���w��Vg~,����v�Ξ�h,G,To��7�<���}��5*3W^�m`���iҭMیEe^����0&���q{��`f;�J3U�{�*��t$mJ�-9�F)FJv������'m{'�3:z��(QY=�&�83!��P��J�,�-C��5�zV����"HO*`�UJX)��L��<�t'z3��Ra���k�|�c�������F��C���aa�!p�Q<Tk����uwon>1T4�����b,���$����:���&����cbw�y���`��uw�}��b\���Z;L��Z��c�<v�.�<�w�<�CO� Օ4K.��@�#��s���u�^�ƎU4�RU ��yGw�}��>`���۝��a�}��\�p�@��ҽ,��{lW����b�r��9 'd)��_����R�*��"5s��������o=UN�ټWU�0�B��N��~���F�ނȝg >LVI�#��2��>ǃ�_b��=�zF���U��ރi(����� -);b�)&�U,I	y�%V�����x�Rt�r�*Dm�ܖI��ǆ?qM�4����Ër[���t��;\��a�V���Z�UVՏ҂DX���Q]�����>�����{��c�gl���a;�2bl���*U������Э"IAs|���S�h��h��+$�}dh�UoG��)��_̮�2�[�2��BƣR=�^��.ڹ����5�\��B2��}ލn~�y�E{�;�i_��ۺu�Wg�a��
c��`;~쐛��溫���tLr~:�Rt�d��'���|�CEI�GF(N����Z,iܕ�#�!c��j1a;� �i�ḟG���Ǒ�[����#IK*�`�h�ǭ���.��ag;m�=�üw�M����c6�P\�9>�h����K7�}æ=�(��},�i�l���:������-�zh����ޱ3O�qh�ȞXla������X��a��L)�zZ7�t��c�v�������Q�[j�RR2�rb��s$/
����h$�d�ͣ�`"giWr뽏ۮަ��֑F:L�0���L�%�vߕqR�\��TJ6��ͤ��O���Z��*��-BCi�)�^��]E��4eX.q���"�Nm"�����GO��kv[Y=�=p%��|h��bSU�hG)A2�+K�O	m��	�P�b�bR(�橈,��ɡ�$�$@w�`u3e�~�[���������y���8�meש�����Gg����	x�|ZM�Q8.��(j�J��b�����GHt� �]�D���+��@�*�����w�m}�u������m��&v�{۪J�����B6��ė���XbE4@����%��Z	�����!����C���T����G��'�(��+���haR5���j�E�+ �؏�ƻU�q��L܍A��%��˹t��Z��2aYܨ���J�G�i�F�"}$�׿}N)IF,��i��F��b����3� #�*!���~/�)�K�2`���r���t�1�B����Q�%0�_JO: ��M4���b�kW�I,��+&U��5��Х�ut�ӄ� ��%�-��N�ꓭ�������D�b�$kP5�*�e߰���!�';�c'N؁ǟt�Ť��{dnl��I�QZ=��C6N�( ��ߌ�JwY���
�q�F4�P�k.E�� �G{�������ԯW)Tyj���:��V�����o?Ie$�f��;ˆ�ГObgq������_�$U�y�\�P�8��1��˾B�vdOҡB�� ��6�p_��t`g��~s�K���.Γ��Ep����+��Z'=9G)�I��W����ǟ:jO�E�↝�Ë�1��������M �u��(Uk]���5ݻ��'�����xoo��\����Gyo;3�{vbj#��+�ӓm�ۻHS�(F.N���՘/y~n��`'��w=j'�a���$x9�����1�p#4�/4L�y-~�j�ݳ�ݤ}�'���lW�5\�m[�<�I1��͡���V�q��/�yrx�T�w9����hH�3���_[HtK���a��*ä�&hu��&�	�_f_{l��Ϸ��,���4����V^�Ff�X�B�}-��qҎ5^��yh�`���L;oЬfI���d�"�b\�������?d?�#?lS���_��}���9�{�~MП-�ƕ'�Vi�"���Pc�蓈[7oক�lE򔎓V���$V%*�������3-+��S�&������J��
�"i>�o4&-���o��|���'>a����][��<jA�9�Cq��x��p=��yU��/�AF���
B.];g�BAv�8i!g��JUjJ�4���Oq��%��o��J�F۲w�foi�}�:*b�Щ�R��KZ��>	7 e��^b;2̉XE�,��L���HS|����E�B��4P�~��zo�UC�(CO��ݥ�shg�Ϊ������_��Yeyb��]�P�Mb|��lI���_�`�
X���h�VVJ�T�蹾υ�HV��(c�XH�V����M�[1�_�驥��%+�������4�{b��C,��M�@C�t����Wc �E	 P��
g�0��+�2�@�%�$�:gmXc�d�P\���o�.sO`�P� E���j��D�j=}}���p֎��H_�>�c������f�=��m���4��{/����Cﷻp�/@<qb���Ϯ��b��/���V�T��N�_�[�r5�R��~�Z��F�'ح�}��ٕW^C�t�m߾ݎ=h���h���^��k 3}4�~a3֒?=��N �XOA�Cl&�H7����*#h_��� n�׽���.,w�����;z�)�`J��*b��M�ҽ;0������S6:5aW��|����ufz��Rc��6�z<C��zR�\�Y���f�0�H�ƞd��osm���lhh?��#��ߓ���b�"D
`,���5�g
��3ӣ���#Ult��9�o��Y���-R��,ܯU�����8�q�
e̺{Ȁum��3y���#h��&CV�^�M�*�g#ɝ�ꓑ/�m��FO�Yl�5
5�ՙQ�����m�5v�m_����_���=�א��A+,N�Ӥ���������k����ib����MD����@�x��2m�1���K�n�iJRy%��vtJ_~x�������M�}yP�����q���5#�5�����,���5ѥlQ ��y*��EHM>�9Ҳ������3�ځjgZ@�Z�lY-ôx���}v�_���T���7[/;�3���-;�����9.�Gї�`+�/Y5�O��Q����Gtz��>���T�6�/"PbʪW=��$P;@��dUz��y�-�y��w���I��"�w݅���u$P���;����3^�Y�T2��ϙT�`�J��!O�:�̓�꥗����ߌ�Z� @�q{��;��Ճ���`K�	Z��F]c%�t-!�=��S���4T�W�\��� Z�4S�,xy������a YI�.a>����fq��_.����A�|������,
��X��@����P��#�s&�hν|W���|!�g�5���`tV � ���"H�p�j{��R��K���$������O��'�{B�9@����v��,m�G�\�dj�^cC�M�X�&1C�w���e��{�Ŀ�0��I�1�D�ێ�U��Y�K�j� �W$��°��<,�6�>c����a�������g���&N��N�s��M�x]ԁ��O�Ⱥ�^���2{�[�h;Nڬ�J�V�X������׷��#���}�[�L���\fO��|�+���~���o���Hk�U{��c��o�A*�j?�#?f��D��w�i��연�ً�S�:c_�­����kw���S����v�7��������^�,C�G���l��Ŧb �s�E�a�E���?����`��݉[��'�=��>o�^����k_koy����l�ٙ&�_�O��͓Y�}���!T�����*v�/��^����NEs�#���xg��R�δ�s���*k8�5��f��c�/��c,���̝�K�&�p�6Wid7�����,�T��J}f�+��a�?1dzW}�~Q���\59.zb���\��"���~;�؁����G��h�~�ï�+�q��vh�	[�������$zl�'��h�3)R�n4��
3��������aļ�\+�����~�ߋ�a�o_�z�>��C6\��
%���*$��2$ȯ懨i���F%�MQ�h�Z�P�ٹ
���H�-45v��U��D��+Ѧf���'��f�I1�4݂?���h�����G��e#�=��.z�gi_CO�"�Ⱥ���c�����:�AO�No���.���iw�V��) �T�v�Iy��X���v�@��l�#�s�uR��=�5�WN��^�w���K�Kڠ�F�؞�)���Z��jxk���w"f>�V����GI��Є=��a��!��Mzi�B�t?�<�Cg;i��幚�Z�\P�P�Q��d�����jy�D�������a|%�Ν�9�q��r�G,Κے�)%�e�&�ꚫl��{wX�y�����[>c6g��Gc嘽z�����]��%?+1b2N���^8`�b�:�}+@&��[��`��l� �*\���D��������V,�ܑ�3����]�L�	9�c �]�;��I�:�Wo��O=���t5̍��,j3�M&󰭳���:}�[;EYw?������s���ڇ~o��=��}�/��ކ�4�|J���㧇Њ�rX���5���"��o���"}��G�Y�����M�3�!y7�IUP�"�FsTⳣ�C�	��	tX'�>l[6L{{��~���/q/թ�����p��y�1,(6�]�.�<2��@'V�N�ˮ���Qֻv���V�͕�Б���7������ֵ~���z���q||Jk@�J�n����1�f_���h�v��~���S�k�����=����[��ã6H����2{χ��=r��m��v�u˓��I��8��m�)�`�\��Q�u!��c���C�^f���P�?G{� s>c�>9d����j���q=].��<��҃��ǋa���g�::���,@��a�7��q����z�Rݓ�/~�!���}���O���eǎں����j^K�ɂUv>U��B���M�L�T
��
����[m]��ֱa�rI���g�_;f���i�5���ǭ�����|{`Z�����.��i"�-r]��`qv�
u	R��d�k��<��St�~q�4Z�3f�^���~��&����f���7���20�}[��9@`LX��X@�+Ju��������){��o�|�V�Y�30m��	ŅYR���fU�F��mB���/L�4��Vp� TR�MZ�H�Z���4�Uz:�Vi���O��-{����4d>�n��፶�r�T�VUM��i�X�����TI截�Pe���ܙEZ��,�J>z�FX������ �zJ�(ИA[�4	l�9uF�tz�V��e���#�!ڶ}�7��LU�/��2��a��unQK&���S�{�B�{�Ǿ��/�+������oj�T�b�홲 .iϺ�hN!���P5�6|I*�d�к�(�)D�@J�	�e��. �\Pe�4{�7m�*��.?57���������*���+��
[��q����,����{h����H]�#lGx�K�F���i����[�H����r�����S����������]�	����A-۾K��/|�v�������g�^�a�h���gao3�`r��d��?�7��4�Ҭ%��0s]h0rc�Զ���#�=�1���]~�5ץ���֋.�Sg&�$_��\ac���j���SvѮ��7�c�s������w|�3���=;`�:[�r]v���bw~�6�H�&x��Ư��߲�������?��ƝG-�N��r����v�]�����Gl��!��9kA*�E���S��㜋l����5 �5�B�̐�R/�&E[%֙Y���ݘ�v�ș�=qh����'=-�M���MX�: 2��ԓ2�[��tc�>R�V����ڥ{v%K���S=��n0q�n��7l��+�O>{��;R���7�����*��-, *�vv@cÆɵ�j�M�<�&�9n�u;�nd���v�Ԧ�����OY�s�M��T��ǩ�X��()�Q5S�t�>"-�7Pj� %�������5R����/ȕ�b�ԗ-pӯR,!qr����Mh�O~�iW�M���|��o�lo���>D����}� ԴY s@����|�L��Evg���]0	D��590��,*_*X�����^�^G�WZmL����4������V3*�Q9�v�j/�~C<ʴz7RC��9u����u�y'z����K�7��m�}[mQ�>ۊ~f���ԋ�����o#�q*�-KR�{IX��\c�ԗ�)�����f߳�蹐),��$�̖�v�t>d'G�d1O�����-��GO�^ȼSl�4K2�T!�t)ev�jV}��3����D@?`/�����?�^p1��[$,?��؍�#���$�d=�i҉\���>2U�F�UCrPD�ׅ�B"vU+��b�ޝ�f�m��>۵klٝ�IK8İ�X W����gKR!�k&ƻ�8������%ݴ6a������R��b��eh�B�H
z�����6���RL����CO���'�o��٩�i҂]�ҷ�lK�~��O�����o��S�㸷������_�_��� v��}�e��U%� �+�Z'�չ�z�:W����~R�o~�[�|�Ϳ���F���p�V��#T;�fg=�'c�7��2��7\����7����wv��q=(N�j��3z�6���n�����߄>�C�5�k�o��L�7]b�������O�������b�1cd/~�_�˴����O�e��࿰����x����<h�_<`���dW�C��S�8v�f۹����f�ul��-���D�1X$����9�`C58��o��$@�>��,ݿ�&c�d��NK�)�r�� �	�}�+����/
�a'�(Q]i;��B�����I��>y�<3,G�禎������#w�o����쪽�T�����Fu��J�Gl+���&�XU B���*M��^�22�k<V&-��=��(MN1�CCR�/Cs�����(mn������(��K�X�6R@�b��`TU.߽נ�]�N�!�l����_�]ņ�~o;3GE���\s�v@1��f(���+_����i��]l�>j��v��xN�x�ɂ���y��ϻl�>5>@,�l0��aZ;x��j�aۖM�Ys�	Ȟ6�ݾ�#�Ig��x���xZ���O�ғ��d�_��o�߳/���� �`0�,7�S@^��\�u��(�dR/�z�q�{T"���v�%lq� ��+؟�309��ۦ/��y�4�����h��y��3����3�ڈ��QU�ӕ����`U�i����X�T���Ob���%�����������̄i�ty����)*��1�m����r*	�{i;u�u�%���aõQ�����@��Ç\h�)�0�����S\ǘ*Tݜ7�6�|*%�z�f���'^�Ŝe��[
� GF�?��m����4� �E�s�0�Pǅ��<l#����3���?���ů~��p ��i �վ�`������=p�v�U�zǖ�Óv�#��񃇭m�E��`Î�ƭ�g�CI���y(�Ī/�0�ƶ�.�W;�`(u��Z(=	9��9����� L�~�{P���u�I
 6n�c{i���?�s۳s�s��گ�������6o]o]}��������%}?h[0I��?�c������CP���Ĕ�����[���8��Y��3�s5۸}�����������k��o{�}��w���w�����-����v�u�l�@¶�]b�$2�M���Ʒ���@]
@��يő�9��e��?���]�����lW���m�̠a�a�9�i��ʺP��zT��Iׂz��-��__m�Q �4��bOG[��;����_�_�������ц�`��N�2 [$����@�����d�j}G�U����rbO�����U�#�Fϴ���ȴ�M����c��6]��u$�?Q�>�Cﲞu�婧\��ww���[�B+�i��D^�V1�uT�O�AjA�q�5A$��ƽ�VQ�$�E+�$��X�� ���ڵU������������鶏��/�.��'u��gaE�YU9�t\|Lv�F;�u���n�i��C�����5�@�"����@���������*�xu�b��h@t����0{1�6�,�HۤE�/W�ȗ��xu�
����e$1�r��B����G��.�+/�1R33ӳ�O��w)��o��bda�J�&��,W��:��L\�҉)��5��M�k�����~��;�?u�$�HO{��R7n���݃�{���nk����/��S�h9~�l�m�AV��4��;��F�٘��UC��sC;��?G��V{�/��#w�Zq=�$x��14M������NZ�M�n��~���!�"�� 36.��$����j�T��$R�&6��3�BN�t>P�j�ɡR�IXS+lq,JG��Z,Y�Aj��'_�VR�U|F&ɦ/T�+IE@��b��zv�X�I^������
�h�Czz���Tðl�j���O[/�68}�kv�7�LP�\�-Q��|��!}�"��Ϋ ��v���M}��y
����p��67����[`#�%��{7�׉Ӄ>[v^�̇`��1��l$�T}��lG��@jn�� �?�����B���#m�H:�1��h�.�Ŋ��PԀи�5WY�LD����Ϳ���WoZG��Y@�\H�i�w\e�x�N^_�.6Oձ�����@���Ԃm��]vl�=�G�g}�.ݳ&��Z�v����C)$u)l�8��0�������v��~���+����?�cO���$&d�-�:=�{A��k Z5�#��퓲��rGl���i��/
�%�ԙ�E��ď|�G�b�9�_|����o|g\�f�]��@��	n��<�	�3ytd�:rϘ)n؎
�n��^sF|��-���Ҩu���#��-չ�n|�����3'�wg���={���Ĭ������pP��lb�;���.ԫJ��@H�;l\̼UI�MM��|��j���i�7Zq�=��Y5�V:����@|��w�����>�џDt�`G�I}��;���a�?;	j��.����9͎rvlԾ�[���EQ�� m��)���B��v�NUe��ZZ�Sh�ff�	�P��T%��`U��L��Ǳc����`r�V+�P��rܪ3�j;}��kԫ-J������#b圥{��3�f�g
�j똜����dY�S�w}��D辰]Ʌ-�!�y��-���>a?��#v۽��s�W$�gAL�"t�sI��h��v�fG�be�f�F�dU/k�t�#Ӣ��X�)�(�O�o@��B!.ׁ�WM��k�I@T%�sf��'�\�Ŭ�y�y�^XL������*��ͻ��ΎE(^������8Ν'��E�z:�9����Y*��3��	H����n��zo��f<�X��EMV7 ���?{oo�Ye������4I�&����/600�fg`�l𶔺[�[�v�����ߵ�s���(��������������g��^�N�v �1@Ş��	|��٣��;�'��s�
��Pq�@y`�ʚeM��\e%?C�ƃ<_K�FG���v-g�(�Fv#_a��� �N�U*iE�z�ka�${e�"�����1���,b�vqا��{`�"�$�҈T��c)e3m����D4��>�*J�Ʉ��<"�,�3����"]6o�L+��kmKga�XAQ��~�EE�x0SRr�X��2V3�J�V�Li�xK�j�Z�o6�3w�H	�X�ǎUۧ?�Q{���ȡ��C��^���ϭ~ҪfU��'۴���#�����wR����.��'?hu0Z�T�����hʝ�6�V��f?U���;�-϶d�Ә��e���h5� �SPf���h,Ͱ����a��v��ӊ�)��y��0/MxgCvN��nǮ;\��.��|����Lk���?���2�ρ{O*��$_Q�f�u�1�㸮kj�{�;P��p��_�{!ߞ��bf�>)2�RQcC�=��Z۽u��!z�����)K�p��#dh\cr�����FZ�t�������L+�i �t2�:���BIN, �Yb�T�>Zkl����g��-w�� \�N�ڢ��-�YZe#�O��/�~'�T��@�7Rr�a��B�b)d�	�k��G�`#���\	�X$�,/��,��x@4�R��eZVhĚ0�K�1�@�D����<;��3�G�.ĦGRM�tc�2����y�6r\�cV\��ڑD��4�r�dLb��X��T�]��T���8��$ )"�)���`&SЭ[�ڼ���Hi�Bݑ�u��b�NWxa���KC����3s������e^^���Ni�o����KH:@��00����u�K�k����`�+>ξ�gT�;$�VyI��JB�Ff�~泟��p���{� t�����a4!t�k�����	���+R�?���J�e��(������C���h����l���r2�>��9���t5�=#�����K��T�v@�2�[5����*	?������/2�����8�/a������*�u�����~��e�~+�V�+�4�4�U6Ax�r!=`�$i������� VF`�?3
z�*��B����ňt�����/��7n�i���̢}����䒏B0S�uɐ�ݕ@�OHN��#G)G��o��R�� �g�����u�x����>
-��<�3�0�0P�'Q�2@�zX��]�ed�rt����a�4J-�N�����;��z|�ˈUe���>�-8��`|�lμ�1��be�=Һb�A��W_�>v7�z/�)�ev�Y������q�N�M�1�.`m�fږ]��㺥Y<���ԣk� ى���2&�+h*-�k����Kf��0۱�vQ��E���2��P���Y�ط��[v�5W�%�a���Aܿ����>��9#�� �m
݉Ka�uﷱ���(f3��92�.V-/��bѰ������w"S��T�: �z�%�f���S����|�Kv�U����Ҭ���n�W�Ǌ���r�%è����(��:�%JS�yמke%̓�E��&���>`Bl�āC��1ILo�E�M�V�ZG�[,�����:(Ȭ�&>��O9�fdd�N�T2v2�)��E�o�{��M�$Ēe�h��@Q���r����Z��"R�ǯ�fS�VX���^���]v�Ёg�������ܒ�V�p�2->|p�,�4ϖh6� B�H�I�5��L�DPrf��a��N~�O`��U�[�����ϲ��Vƒ���\��=�݇M®��J�����#�C0�?21��Q����l�>��e�X/Ծ:�Uj��\����VD�0]���b&�N�Iehx4��� �%�s"L]��*9���tx*X�Ӄr��%p �scIξ��ɇl�����nT�����$+��17��K���L�F��C��_*�����THץ߇�9+h��3�v	h	`��C�w�2��Sׯ?�Xu�jXs��K�����% �` ��:`'8�U6��j-Hz~)kH2�	˞Ract�I�%��(�QsJ	�f�!�}��"Z68��t���
�K�8�u���e��`M'"���Ќ���lo�p��.@�L�a_Ōi���k�)c��-<�R����Od�N\��u����`�v ��(�
��K��K�2����Q��2�߅�3x/��Jz�8�U��VYQ�@Yk%ʯE�([i������nt�61����-oy�}�[��F�p�S�7XA����!���5XQ��aJsz@ΑtXv���?o%{�ǵWݔ���q�����YX���,�"��ON%h��ڛ�g�i�nK5�$#����x�7�1�YS�^D2�c�sk�=�5NG� ^%Ñ�>[�f��ݻ�^k���@\�i�]y��<!ya�&�meě����ɻ��{�byϻnbp}��@� �`O�o��Ohl��-���S\��וt�'ۏ�~�Ӯ{�hƊ�8�a���m�c��*��|X��~�q�����}��J�v�Wۣ��Ԣ:�-���� �Nuu���g��m]���#�����Ʈ�ɒ��6!�G(?6N����o����t�d4z���a�i?�s�j�N.���Z���>��n����VfE[$���E6c�<b7�,�F`䈭i�[+�37���V0%�.*�TV��i�C����x�~��S+t3����w������->�ι16���G<�'�h�VY��{�
bI�0�_t�s8��B�EwO����+l�)+�o�-[v���X<�I�bq����5��+*-�R��ϳ�l�H������ʋ�`sr(��Xb����ei��u�J{�w�	ܜC��'�?`���*,�\n����Pާ�4�q*�Z���S�a#%n�;���}�_m��-��x�Id�o 8%�0r?��>���M�7!���H�Ͼ����Y���[~g�d�q�	�u�9h���xUf��-m�17R>谦�f[�q=��2�N��A�:d�ӧ����4�S�ʘZE�*�y����e�֯0��p�]й'.E�˒�(�ټw����@
���Y��r�^�@I$ӏd��:�U$�J��z�P�T Lפ���/���>ZHe;�BI�b����	�7�Y���e�D^tՏ���Ƥe���!.g�k�jM�LY�y}�&i	�nAk%�q؂�J�<W�7�}LQ �R�C�Ԭ�	JCA�������p���bȚg9��C�Íu/X�*����G|���^��&�O|�0�z9���־f�g�|% 渶-̀��q�U���֋�� �����@���!�3y���G��i��ñ ���OL���u�I'e�ԩ��j��)]� �[%*�ٱ>�Q{E,�Qr�n[���n&`OU�T�r��ӈh�����
���q>��86*�n�Y�}�K_���~�X7�f��j�x�	�ߋP��zU��Dr� �f}>d�:.����8$��DX�	�o`RB��y�H7f4�S���)v�;�f�oڋ�!����}�^���W^���J�(��X�}HE�&��: ���ᥑmYX���v���/���ۼa1q%;�
?��O�<f[M�؅W�ۮ��V=��=��#�l�����d\�p��̕+�('��h�}�3������+.��v�;��.��f������H�G�)!���?��v��޵�>��DL`��\_����NR�]jްt^i��0��i.3����W4{`��D�k":���Gm�����#��W^n�S��E�``5��I��@~B������4~]������d3*�N�R^u*������@����˿��y� ���i�ڬ���%��,����M�<#AZ~Nb>�rT�U�)��G���a�� cl�9�g��G7�.Tg5��8�Jc�R��D��˷�.�[������f����Z�`�~�_��*ª�/��}�C��#����@�.�"Q�/�"'��]�V�:%^RPD���}U;�P���*�Cr�����k���Rn.���6k�����ˁt�� � `t0��	���ՙ����#�^?یe�&t�Y���e�8�!�2/�k)��"�쑮G&�G�̵����3����]�%��b�,�Q  ��u��X��Z�ct��6J��.�3d\@�w� �g���3Z�!��f�*�J{a�I��d���ןʂ���)&NC|G�����#?}������/���5��WY3���2]!�$��pW�3J!@��%�$�.`t� �uC��3�M����)Tf
�c0;7rI�%2+2	��@��^1f������!�CR�ѽ�5j+�l19��o�Y���: �8hG5�G�( N��	�G����j@k2��s_��,U��
�N_�i r�N����K�p%�ҩ��k�e��~�Y2U5��˟3��$���9�H�����P9Q݅ѱ����bU�/��5�f�$ћ#x���1��;Ar��G<��D�"��i�� �LyoAyi����h�m���Hg��mŢK�0���O���W�Zs+�`�X�}�/̶M��J纒�iI�Qg����{Y/�!<� &}윳�ه?p�:����S��F��<�"A����eM�V���xЖ���J����UO���>����Kм�r��3���k)�^����m�v߽���� Ʋ�z��ٖ'-Z�s$���ȳ�>Ͼ���pI�w��M;����w�����{�U��o}�rѢ}�_ᵖ#�i�t��,,E^�r�>����v�Z��d�*q �a�v�P��1m��[y��L���������ꧬ�V������j�4�Tak����=x�cVQZe�]x9��K�Бöx�"�9�D3F-�a��}������Jk�Ru��2�:�@ov����E7��e���������+�c#�*�q��an戧�P���NU�c+&���0N"�1^3.�#���V�����%������}�c؋����V6s�-[���:��������%9?�\��0.�]9-��DDJ-r��,LU�z�Y�t߸��V�(�F2k&Y�@$;�E���n�
�}3־@W.Yj{��~��U�ꨢD�n�<:M(I�� ]X$Ϣ����z�)����{�83�"(%Lp@���4��@tl��Cb�F�R p�4d�v��Yv����Npf6 ?��x,
䞰��' �Tn��WuQ����`��k`'2`��CR�������졕<��ob�t2������ >�gV���_{��.������~*`��ʴ���l ���ힺ�͛�I�a��K�;���A<yO/��� k�:`�q��4@�ِ� �� L��H�Օ6�O�~�#�x��'�j"��	1����y�Xрɕ���Κ�lǒ�Rr����.�'��d% ����7��L�~����m)`�$8�����:l_�*z���ď�Z8�|\BPb��륗���q�ud�D�M��K�/^wh�y�d���[�I����XE�nT��S)�=7@�j&S	W�z�ڂf�	�0��3;�!��LUl����Ҡ���T@������p�͙���O+��� |��1��ϝ;�mJ�`[�n�i���<B��.�hp��@Bf����D��C�4��n�}8˓,T��[�^e��"-Y7��i�	`��gPogV������'>m��ﱓ��ns�nj�������_5u��w޹�QE��fخ];m���K�Gg�wc �� !�$y�0~�%��!?+���.;���֍[9����9�1s��o���^��a��e4A��v���6�d�������a�=�]u�h�
I�iZc�fI~���W�w0p}汇l���6e�i�b,��b�{AF1;�tJ�4[�z�=��j�яnu�\6@qF��pVDL�@\�~�̻ଳ��nт����9�������M%���vҩ����W�-^���qO�]k7�^$1m�����4�qj�O�����5n�7��^3cYG&������#�R�a��1���"�G�=�ߗ�F�hc�'Q�,�@����CO����,�!�`b� b������ۊJ�u���m��Z3�ÁR4F%�'`qmﱝ6��8�~�ﭱc�6�m�ﵵ란��t��0a�0h��!�<���%U�s��r��� �)Xj��ōT�i~�x���L;��:1=���h�F6�'�H�L��Cg�y�zTfB&�4<V����h@�!����[�� �jI�	��&�%(��S�)��=L�R2>0Q�m����,7��!k$�t'�^�X#Ϙ�Ag�4ٸRd���E�	�A9��+c�a����J�-ʃ���>�(��*����P������(�ݠ��~�����b.x?q<Пvul�&!:W�J׭���o����^�ܿ|���ì�^Gס���1�}�q{��އH�,�a��3l���-�@@����AyR�D��ф�^F�t3�-���8���Ȍ>1
 *	@�� L�j�ײP������w�z@�z1Vb��(M�$��������K��) �h3@�~^v�܈в=�E�.~��Y�Y���}~���p`����B��׭�?���贈�?�^�\*��ʂ��A-M��A؉�*�����^�B��7u��~xS�u��"}���>7R�>E���h�ߢa��@��`I;�DY{���@l�֟J���JZ��,��9�أq�� �y��%#�bIJj�]v��ӧP���߫t4aq�18��2)#T��u�\{0?<H�T��(#�-iGe.�dN�/�et�M�O��*�5�x�v�X��$a~nSAzG��xW_�@k4��=�̅�M���g֮�h���8@h�v��n[p�bX����<l" ��>��e���%$v$oh\S`�b`�N_��54�ıAF��������}+�]�6�;)>h�7b��y��`�ێ�{)Q��T��.YN�a�m��2�E�9�\�V)�v״�3t3�K� 'ݖM-���9�:��[���N�E��� �� �G�gh�jj;m4:���~ކ�2,�$�b1��m9�&��ι�<�f5vڊS�;41Yz�(ʤ���c׿��u�a����X|��eE٦�kl����;�b�E͹3N�2��H��F ۃ	�L}U���z� � UZRֽ5>����,��gȆ�KG����>CJ4�6w�LYt&ug-��1Zb\���+�>�&T	A���$ ��	2���eΉ�~k����7�i�ηo|�; �N�����w�϶l\m�?���~�";���;7=�Fes�b�6�{�f'j�p�d�I0��@�G�ʼ���]��Ɇ�@Ip4�ܨ8{�H�~�kR�2�C�\��̈ �ea҄���B:c*`�F��3�N�L4c��h��(6,��#HL:�UK�X��x����o����hl ��G N�h��\��c�Ґ���xr�"�V{8�Dz����KL��J#��+RCz��?P���xP畂� �G�<�K ©�?�G�xP�ˍ���S����A�UW���
��Q�[���'hL����3�@7A��"����3z�"���������6DV�^򹛬_uv"jm��@zQ% ���QG�ھ={���� FL�N�C��^!���ʙȰ&,T�v�h��4r�WY�� �1#�N��+g�A��}:hd�+f͵`:��CD��<�!��p_'I�`���N��
U2�����D�a��#T��#44Z����F�,[v
"�
���@��s�K*}�>��mu�	 H;&��kJ���?��нS���%�_�������sFW�DĆ���W�z>��)� ���V̔�MeAS2U�O�D��ߧ��g=�r�^&(ǆ����XM�a�ϡ+��I�%#g=p���5�}*�;�U0�Y���С�v�m���[`d`wĶ
x��ң���|�(�I]�Q�h:��HT6�3~�m�>`��>��b������y�.��d��A�q�.����}��P@yM�z���V�R�83h�t�mP�:�D2~��~�9O��,��榣q���
83��ct�xW-�ۈ%j��G����Q'�A$2	iK��x�q�ٜ]��4|��X�����F�I�d�R�]���Wd��J�YԆ���hk�쵲"L\{����#�\!��?�
W�K�{��oVj>��T�F�<�D#��a��sg�k�}�+ߠ�j�ϣ���#�-�5�,�CW{R��1̢�����{��|��v��7C��70vtji��o��Wٷv�z�M���L�%׼�X��շq_��AbF3���ʰ�Xd���a_��/XSK�UV�s/"�ky�n���2A������ڷ�O~�}�f6����)�2] �E�=��Q!�)Wg4�0���F��a�ka}��44���O���h��� �k�nJ)=2z��h6t���	��H�)4�bfFYU"u�;~�_*�x��xW)x�O)�疱1"�u���c�1`E�7܉+������F{d����(��b�iv�?�G�D�^�c����\������|���I���g���B>2'���0���+�J�����쁙pj��G���I\߃�5	j_j���HF��Q\1�Z����q�8�`�ȡ�ȴ���8ˍ����v�ܚ:	|��b�;B[v�O�jc�۾/v �$H��д�9�96�2㦢�ddG���$�!��Y.��<hv��4�;$��EO�F���-^lrԠ^�g|�Ù4	�u	��9�l�,�$ �j�8�,��ы:tG\L*�y��6>�<�t���s��A�ׁ�R]G�
��RX�>�'?�W\N�th�/�?�A!�`j�\݃x4e����43���!VCl@�NH����Nґ��Kp����<3�*�Kx+�G�����;
���$6Cɕ�GS仔M����`����ǡ/�Fc����UVg�>����A�� � ��,�Y_o�u�`�~[T��>"8�[Yw�K���pw"a�Vy5�M/5y���X\�z�a�73co�e��a?A�^��8�f����tE�j�4K*_�]x�&���[BV��!�G�����8 :1�"�D� w�׿	���#�	�se�>Z,4���U��:HR��  b����x�ֿ�(�+�g.l����ܬ�W�%�)����5 K,�>�7)p?ӆ9��lu?���A�*�0��X��z5�V�w�
��bF����W뻫 3ZO9>MW,z�b:�Z�4� �	��d��@�FX��/��NԧX-dY.dϥ�A���K0�HM�c��٬%�p���҆uZ׶�&Hk�Y4q�����0>%Ɍd��P�ޟ�t6J7n�~�M��sJrY�}��R>�,�Z�� >W���~R�F�iIaH�`&gH��w���g�?}���� ��z������4��Ԏ����c?�Ńxg�!�I#�2K�͞{~ɨt�t6�٢�WX��fRr�lξk��60��d'�8�MJ�ґ<�ع�>R�H�k��+δ
��w�h�7h3+�a��7�����&��#��i\�v���Ѝ�%0����ԙ�Nu���@Oet쩵��
;�i	�l�c���6� 0�ςt(R�v�p���]���M:��J������}���bK����[f���!�;�A�6���3�J�b��
�(�{5��2�זI�
��KG������ lhb8�MLe�+��HF�u�Y�7n�|F/�M��Z���jC��Vu� �)Ss͆�LX� �x�����A%�۬ @�� e_���V�hD���@}_@��w=d����m���{���=x�!���vly-e8L_�5�G-�&�!@���yW���`з�!�˽�|����3y�7ԁ6	���%/��*	qP�"�� �D0�-&��u�0!Rm�47� �H�H(q����Ud+�Twߧ�����1OMmܨ���1T�w�Y'�kGe�J֗���#͐ӳF'�	l"s�&ȸz��ܥ_ϟ�붟��8v�";�h�U�[`G������!�z�R�1��r{W�EkV'��}a�t�c0�h�:C*{�ܿ+T��sW���v���3J �Jb&/9���C7d&6�P��g�@3&�U�r����˻0#��IB�4���l��¾cj����&���P�ȧ�ԃ@?��T��+JIH�P����XY���z1�L���ܗ��'&�}4o���<��O^��f���ێ��f�?�\�%��*VK`D�Ҋ����1������=�>}A�G]����(5�.���A*��M��D�I@:t?���=w �?��	�j@u���/�6��A��^`ܵwZ�f�J�*��.#�\9�Uc+4JG�ȯ�ɦ�N�h���W	��ǽ�d��	�o@,J�
��X��uj�Jf?�������DW#��>j��Pu6��������cl�LA�~��蝸�!y��3T]�� �3jӱ~� x� bF`��`/��b5Z�bɐG3�f�j̏��f4T� �%�
�oj�Z����͵�eT�� ����v����`�-��d)F�e��o���D^/������ו��|yV��e��3:����Z�F�_�٬�A��Q����b�3(��!��b.#�vn�bw߳ʪ�/������8��}�fͷ�THއ����ζ� V��3�.��R��?���ǚ���P�=��:[��F����~�U�k;ڲ��E��W���g)f�ľ��"ա�l�:oX�����U�L~��QsU0ǟ��h��������0��d�?��^�����n�wi�	�f5�k�< �̙v�i+)cγ��Z�{��޼J#ϧ�M�c3�] NUn5c��ϴK.<�d#371a�_� %��h5��m� 3+s�J�V�H5�����-v[qIפ��c��P��H�����
��5�+Ԩ�DO*c�	7p��ˤfJeEi��y�"�F(|��X&l$餸��=�T������Ťl����3A�}dÝ|b����0�����>w�O������t
])1��?���Ι��_�{Z-8y��U�
�����Q�KAS���B�;L��0%=	D8�2ᯈ	u]�	_���Y�h��(v�g��
]X�ִ�c������"�րdʐC��H'�úb�2@T�؃`������^nJa�񫻻���t5���H����E�A)�%��q����J��˷M A��se�
��a������N^I5Y��j�����{���k�( Y�b��������2/K��J�}�~o��!0���j��K���5���Ҩ�U�Խ��Ld��II�W�e�ƙ`9χ�}�~N,d�\��%e�Yj���-` ��A��)}A6��8�ab�	㰍����y������8��YfL)=Q)sd⸟��iM �(�W��"(eD���I� B��"��r���%�	؍DZ�`�SB8���e� �C�K���Y�~�>>M��x6����K�Mf�[n���qO)}/%/ٳxY���є���n��o qh���A���$�a�S�)��h�����R%0DxNt�<�)��   ���T	��]�?J`L�10�t�1Ht/FY�I�U_���aJ)f�+����C�6����J�U� U���G<�G[:S��"H�s_�A�R4~U��B��R"�&��q��0=l�����uo����֫�;��Oۈ�r݆��s�.�
��W�v,�ZI��r����sρ]�=};��L>�Rt+���@���ʘ�l朎H�.�dEt��R� �5��9�|Ԟ��"k)���A|�����R~M��Z�Z�F��gڂ��9F���W�6="�ZE��1������}X�dYi�T{�Χx�Ö���J��&J�Uhe:I�`�eC�����$<Iv������JDH�#�{l��*�m�*29���1�fȇ����'E��Esl�bƪ-�jȰ{�=�L���x���4l���щ���|
{\�F3�r,�>�A��K��V�k,ac�ui��|*7��0�V6B���ںzonr������|�u�죩��!���2��I{ϥ�0�r�4ERFv��[���a��M񭭭��7l�ƍ��*,'�d��'�)P�? ���	9'333>s7e��b��3�IwC���(?�����w�_Jg (��:1H��,	EiCW@��ͱ[�痶����&��E��W��������A�2$:��*f�=x�kش�=�ù��   IDAT(@�:,F�v�88�o����z����CW��.��q�.9�|[�lj���4B�3�#%�*f�LsB�hzu������y!�w����
KH-W<_tl2r.�:��(dC��bF�>#3B+��n�����(�,�zЁ��	����B��aӆ��� �ȫv�ń�����c��_M���t��OO�� E���A��x�I��\��*�y7�VYs�@��q'���3��`=&��dO�f
��'�N�{,��6��\���+�E?�݁?�!~Nz/�O����L¶�Ͽ�*/���e~���<���l/v�_R�v�5[���C{lae�͞^��t{�rV,?�����6�KI@��7:(߹���x"��&�[,��Q�c9�{8d{���������E��s5�~)>�|�(h&�?W��u���W��$kjDPÀtv��U�U��ͫ�N/� Y���#��_̤�@^V���a���W4a�9�!����˸�]Tft1��3uiZ{N-�c~�Z�c�<��i��>�$�h�����J�z�BV�貒�ϛ7ߵ���S2�r��7�9J~/�z�� Qye,Ppm�tʵ�6ڞ�۸�^�M<'���#�n��pw*�XXZc����~�������}7�4��=�kA��s�F��m%S�����nD�������;������iy���9��-�2��N��ˢ���`Ni)�1���B�ݕ4%	�΄�����x v&ݗ�^v	]���/_���Y!�.��\��ǳxfxh���ٳk�#h����#8�^���E�֋W��2eU8l�3����OL�������eM�VHpې�4И�_Zn�1�������F.��X��:�lf��b�@n�ƈ�n�X���!��lX�i�+��=�plƺw������ޏ���z��Z�LaTR4�+�S����)�0�l{�����E���{�Z)9H��/�i�Mń�Gp�:�dRJ#�J���&��\O�_U�#�����d��Vi�����5� �q�G=v�����vvw�Ǎ�e1��D,�3
F5���D����j��$`� >�N<d=8x,S~B��&q�6�~^�tc�����2���J��l,�$��o��ٳ�UO�����J��-;���[?�m��5����E�8% l��?��T"�D4�%�pv,,RUWj(�@���G� ;�v@���e� y�g�<8&��)��S� ���p��"Z��ccF`QQ�&���@��J6�a���H���4��5��`c���|�FdͱY�ڶM,#���������g��wPB��E$�.�q��Id�
�*�M�o��\�D���:	��g٢��6b,�t ��~��1�ߩ?�d��^���rY(?t&�+���OJZ���W5�����#u��j��3�^2s?�?�Rp�pG��S�3��{���4���ANM`]�Yb�1��,���HY[dӱ;V[���r�������z`�?x�p�% �FY#�����t K
~h!T~�{`= ���QA<�{��W�ݰ!G(}� >r��-6g�<��BO�L�%��^���5\*��|���zb��H@
����<��LE�Mӎ���L�7��Hz�.�a  &$i	�A�ӡ�k�{�J�b_���:��}�F/+c�^�E;I~��U9��A���� �@cHsZ���ku����|.���b��2����h^su���:�U# �4@���yt@�юQ� ��J��xV�����v 證 *5��yU��\7$��ֽ�Re����~+�͠�o���'�1[Bw]? U�\��S�WF`�b��x4 F�D_��G ɔg0�����j�'Ic�i��Ky����لb��1�5?�s+����C�1V���5��$:�(�v�)[����`�9e>5c��gw{3�#<�Į��*b�C�-�؃���y�y��� �d�y�I�� �,v?7���D�������c�۶;:L��&�⽗��"!�a�?�c�3v /طw�-D�`���l��8��yč]��H�j;b�f��L��1�/&���J��A�
����M-�#����H�����}�ف�k,.�؆+��0���CV���@SR�Z�����^�L�.@vNN�8��-�{rf������_�,�E�a#�I쎞|~���#`�L������?�~=��_�k�# e�I璱^���9�M��UL���n������W�� 
^��将Dt�!�P��'�0t8��+�{Ǔ��P*tM�*��f�[[�,����+��>(�3�9�)�C뭼��6l|�	�s���W��wԴY-�Ѱ<���}*-A����:�A���x�dE�&�G�����̓��������̀�����/�ܦ�ݽ�k�+͌�"k��R��`Xy|����nbc��i�*�-�@Gı���jR����gB��Uϡ�0v�Q�0
u�����׭�b5T$RcCd^T���de1*	��A9�@%i�$�>�d~9���M�U�����.1�*G��Q�އ�5�w���K�b&|��Tꋠ3��ch���(�Hd�����! zJ)�!�5�� v�<�:~������X��D��v�Hd� /0�E�&y�q^��&Jö)c�:h���*.˳��Ƣ�����"��,
 ��B,>�A��'q�B��O&Ѐw2�[g�$>����<54���|ػ�W�i���,�U=��s�ן�\��!�X�ϫX֍��( ��^%��>JkCr	��~/Y�7��z�3qdqܫT��d.�`�}�eD���\����ɢ *Ʃ���K��O�g��M��.�I�WIքʢ�M5a�N���OM�h(���/K�<:��c�N2v#�c�z���*�`��o��u>̓�@!�3����K ��Q�n���d�K &�91���3gL�z�e�]t�s��^�¾���ұ�M���BbϑC���Z�{Jݮ���"IS�p�ρuͣ<��a��������A+D������+�J1S����G�?h�~K�b����z� �*���b��k�N�2I��F�i����\�0�/
f����r�e����F���M�)+%�C�j�g6Z���izh�h5�����vٴ�və�l���v�oo�ːJ��^�����lƼ�6��w���SJ�thƒ�J ����v��'Y*>��1�I���XC�?y��w��v��J���Qt�K����~��P�oF�#���qr���4�hlS1�!^g���.�O�g�{�
X�Uť��f:�문���X[��$KĆc
��=-�VD�PE��P���~[�n��[����� ��m٥�]F	2�����;�u/v��:��@Z�L˥4�8�F�a��#h�z3���b�j����h�(g<-t$O��k.���7����*	ʨR��"Ĕ%��9��nziC�@)lH7����(����U�$BK��^����Fਫ�^ul��|���6�v�sϿG��X��k1�;
���tC��;�=<B�B&2�f�aUڑ�G��s�E�Wp�s�7z��Z ��H��R��X(�ƶZki��Yhi:�[@��P4�4F��=� �
����p��r�݈2��AK�P�ZNB�������L F�TVa�v�A��A�����_�lGq ��ʛC��yn�P �v{	�9����^M�J�oԳ
�\&@b�����
:�=��h_���8��"� 4xbė3�)�~d}�W����[h��C�D��X���`�}��x3�p�:�"�f�}d�C(��fD�EVQr4؀�co���,.*�����{��!�!���f��8�Ћ�( $"ݾ��%��'�,���;1U�*!/@���Ǟ�{�KŤ��\�E�8eJ�]pٕV�c�=��S^���p�~>̌ii��$��!;`#�8fQ
4�=��ܱ͟{%��E}�`�y�Fc�t�����8���8�=z\���94S����Qy�$��:u� l֬[o9y���C�%�����	���,�y�I�̚t�����]$��ᐕVJ^s�	�~�%��{�s�"��5+�LN����C�ni� ��$��I���Wc��V�`��a"�,�h�f0S�m�.ʬj�釅:dx���-0I��G���G�Ձ�Bu^���M�:Y�X_�耻H8��r  �Z�" �d\�u^͙���?�d�{��q���-��3O�F�[�+�*K���G�����.BsM)�PM��R�$I(�M:GFa��ܼ���;>�);��K�߿�%+�2ž��'��(S�|�\nN6eG�"<���l��V�mW]{!�i�6��D�J�ً�{�خ�}�n����.��p	D73�����l�>��=�8��1s���'�@�3N?�1�����@]c��s���9M��N�B�#���hb7uN󚭸�'s�R`��irh ���Zb��A:��G� ��k?�N�dF7e�i[�.LSRRh���SZ�H����߶�\�=�s�nSu��Yk�)��,-���*?O�����c�Z;��(�dk���o�~�y��MM^E�L[��^�@���U؅���f�icUj�{tC43�@���z����%��<�#�B������`gĤE�L����
�%r��z��wu@�;;h�O��}���0�˲��ȇ}�·����l�b�����!{����|�$J*����x�]
j��һ�d�p�|V#R�������(J���b>2�R]�p��N�����3��T��+�4��&2�xf?���;�v��Ю��S�XP�T�eԊ�@7��("�dD��������a�� p��u(?EB�kθ{����PP�N]��-��F ��Va�Ek$<^����c����������&0�NA?�#[ B��s�\�:ɴ��F������(a�����q�*���\�`�Z�Tx9_v���諒dϩ��ˬ�X� �M���BJ�BeW����xV"|��c/v���Pʖ��( b�Yq�y� ��xZ�ݙ���9o��,�}��R��{Er����^C����Ğ%��G܋��&4�d0�X�C���g���-�{���K!��Oo����ixR��~5��Pi�$k����a̡}.�kUt�D��_�YN𺷚� ��T�_�,�V�>�1@B2]��9l�=ES�X��a���Rg%W������ �J��|���{`�|���Y��������bfv���N皓3#�,p���x�OiT�S���G̒kp� �6⶚�rK`�H��P>t����Tm�91�Dw964��D�2�������d�N7%$��c-�(6s/t�:�8��D%O5C�p��<xn�V_�9�c��w�[n���̢��Yffq�ka��k�{�>��i#G�+ �8�YVI��}֙Xb�
hN�D���|�!�D�c;�P�����a���X�Zٱy�]|�J+�$���p���e�� .��ީt��Ql��v�F�8�u?��w���=�KXۀ9وd�a���F��9��O|�z����������a/����e�ͮ��ӟ�֞�ak�����F+��n�|�(-.����m�f{��5����(MR�D>�5��{;���c�<L����B�6�������8m�֕�k�F�fS�=��(����:�2�2� �Жm��?%�ą�ڣ��T�C�ǈ!ڿ0���d����O0x�6	v��n��{���b[��0��>�aE1U�]�[�B�|�z�L)�ةu6�/�u��A�?�F�K��Elޢ���ʑA��ñWXa�;$I�u)�t�;_�聉_�5�/g8{�
��k)S��j��j��m��U�M���f$A�����G�׿��L��v��csf�����O~Z���L�����񩣧��v�P�M ���a& x#�����a͌�^��_..� W[A5�hv^:e��&o뮨����,�9Vg�-<ǉ8;��k��g\��- ����Z�zQ	.��M���wA��Z�2��Z,E
�3F(�1cb2a�D��d�IP��ʈ�S�6&� QVdR�^��'�:':׿�������ax�Ý���*�{�����"&����3S��Xxo��D�P�Ah��WiE@1<V)��'M�[n8y��OL9_"#�������P�y?Z��d:#�� �
�̞)S>�bP�0RӋ�3��U�V
�������f; �j��d*#Ic� �T%�I�#A��� �,9��ڇo� {y�aЏ=�����RLpH��k����ZJ�U��܅v�qN�2���N�눡��:�2�/���KD$ۃ�o/�W��I0r3��,���`F8���
i� t��(d��1;��܏F��(if�7=�x�o"�G,���q�a
� �H�G%��Orv��4�P�-E��S@�}��s	�џ�C��s�F��h��yF��]��8�x�j�t|j�� `����9X�<�-Q�J�ka��3j�0eZ.���d�u���F�F���"��x�V:1��濣T=Ta a�'��=s�:��;�gU�� /�,�������O��7�2��lE�T+.-�m;w�O>�%���*�s�IV�s��wa ���R�������R�#%G�a�6oB�߅�N<�ܜb;�Z����＞�c`+� ����-�-�� ��5*�a��<�RFm����� �}��� Z0� �i6�t��fL��j�E��گo��BUzc^�G���
�L�5t\f[voB�UXNc}���Ƴ/<�J��XNa�� @�8e��G��nQ�3�ej�tf\.kF��L�\k/�~>K�P�����dq�}����VP�G�����yi�=9�:k')I��4��B���M⬑Se�>R�
�=y婶a�Ɖ�	�y�m�^H����Őv����fQ>r�(8�Ǟz��-����z��g����6o�nS��e0;#� �j&�P�&�o�� ��]_ߐ��Ը���9U#��-��6b
֣0>X���z_���"|8��|����p�@�#p�fX;$J�NL�T�ڡ��@/�3`�w��p�ͦP�.�/�o��y[O�if�W�Ԋ�d�قy����{+{MC2A9��y��C��7�&&�EO��K:��/��0�u`b(�_���`]."�,���&�W',�њf��4�,c����i5M!���cCX���n�>�0��#���%� #�T�=�i�ljX"h�!�"���7��V�BÐ�Χ���q��df�4�<��y��4��5@7T�9�y�̢�_����^`7�\�/��K�LI�����}�y��&�3E)���u����l����"��JK4{�j��-�Η!��[����K+��#�=�{���hR�+���v��f��&T�u�v)Њ��D����d���$L.��{$���BI6�Yz&5 �H;��=-�H���z;@i+A�?㹺{�,����_�׉B�r{"��	SaM�a{;ɺ���I$xZ�$��3��U��7��ϔ����J6�g���N��9#Ɉ�Æx�~� ���(��"�@uК�$��k���Q��@�(�������L�tX�J�ڏ#�@ԅ��>(J��k(`#epɾW��ZȭJR��Al�<m�0��CU�&�̅��l|�!\�hW�tS�ON�J���	���a��(��)���.$^V!�N�xȊC	�>�����`?x��0F	��`j��*�YD�x/++���ls謤��o�~�:c6	��i*�^q��Y� �*^���F-^�0n�"ue����=l����g�����яa�x�L���fG�w���{:�K`53� ��,u�&�����`Q�����3��e�����m%('��hꃚ�T�*�d�ת}�+ߢӴ�x����V>m���::��'���@c/6/b�c�wc����]<���4��P��d(v/4�*Yx��s�G��"�C�V�A��J30%~WB'm3DU�X��@�w'Z��ޅ�6�؄^Kc�J���%��H��CYU�J��`�/X�N�-ۋq�@sk�ǐ$$,�	�t�e�?N�@p��z�W� E���F�����Z�H�{�m��F�-d���_�1�c2	����Ғ��>V��Wֽ���xϽ�5#d q�u ){t*\%�PV�J埰��+�K�_�X0����W+:� �D?���]
PJɲl�J$�_yƙ��w�;���][���U0�+Ͷ�}�vo�j���gټ�����Vơ<�&��m�eĘt|A�������WȔ7�k�����k�����1Ds���9�Θ�c��B�5�9g�\u�m�q�N���Y:�䡄�^搃cd�h�8���XD���d����l�bqcxd'�0��A&�HV�L{��N�yg%p���%�ƹ�z�Fǧ�j]�4��&��z���_~��d@�G,IX|���W* 02���p+�`���p�+��ߋ���4�-��@E.i�B���o  dS �W��F������Hӿivg�+,lS�?��)^T�X�Y�.v��{����#��aX ��XH���(�7Gf}��G1	��G���(��t&t�%�=ǂ^�5RG~l:��麃�.*�⯻c�S :qg��5hk :c��,��ØT
X�s<�H���P*ϺQ�lqT;d�WeHV#��B,r]���C~�� ZI>���E�sm�n�>|OEy���d(--a��:��Ы5Sv�~,Q�Xy�͘� g��J6�0*�	H����`�3�����7�ϱ�*.mfw,�je�0C����Ĕ���t�R����Yͱ�^��}е�ع����t�im�� �z���z��w��w4�����qE<V���H�O2���q!u�z��ߍaI���3�9A��P��� �Ά�&�$��l���ۻ�ܳϵ��f9����C�d�'j:�d=�����u���rcW�nc-�Y�����f;��C����}�nt��b%�b��w�؜%+"[��i3q3Y��c�������ChĚ?r�g܎u��z�v4#�?��s�`[=V-v�G>be.����w>p��r��|�Z������H�溋a��H ����7���M�>�nz����R�3OmA��n{�V�n�Eͪ�b+����nU��Jx<�e���jq�T][}���I�<Al� ��x\ϭ��)A2��2�29�����F�q���JjQ��bݱF *��3y�Z��54�����(0�e�Q@_b h�[0��Ϧք֫�O�
2p��g>G�	�"���w:R�X%�h��ŋ��D�#u�!���ѿ�<�8l��� cZ�["ݨN��9B ,Є�`�7*��@?�_���X��}2[����*�F%}��0��9��2�(�8K��2 ���)>(���{�e�7��u{�����qK��p3���*������3C�o��+%����5xM�
E��Mm<�CC�S��<�T��+����tPyy#3� �@����Z	��릴�d�\�-]y��Z�F��{�JW���G�gkhmyE�����6���s�L�{,cb�ǁ��f�]���,�/.��}�/R:ӽ�!A��9kPZ������R���I��0��+��Z��H&}��޼{W|�Ƈ׸w�ʏ)�o|Ca��fD��Pף�$�N�p�T�q�������`���v��A�5؏�"�Į�����%^_e8ճuRn�h{�`D%F��1�KꞕI%5^�?�����;?'�Տ6i|SI5E0yh�Ko�=��}��1��iX7̲'�|��o�9�x`� c�	�t��r��ir�N�Kc�WPb��W���'/�M��C��JE��`D�s���e�K����2Xw���;��)0��q$.�����l3kF%����O�a+���4��A���{sW�y�,�:�k�@��V�_d��t ����P����'%�Z�-���K�ѱ��D��M3]N��ǚh���\��gPwD}6�[*�S� � 7;�\��2zG�ƈ��7�N�a*ېy�b�����#��xdf�E9B��xS�F�Kø��z��$�u�*�Qb@4�A:�D���6�"k|ƨ�wB�rLu�ʐ=������T���]M�(��S���X#ŕik�]흘e��!QI�����:p>1/К[VZ^e]ܯ���  4�%� �)��{�i��0<4�ʄ�)�E;	z#�ڱ�L��������XA�2;�`LV
�i�ސT�Z@��	�¦�ҳ����u�15�v��A7~���=��k�>��i����e6s�?���̴/<�t��/.��X[�!��YK�`d�S��+%���"0���Ab������(���d�ԀP����.��*{��g�̡1ĿKɤ�z#)��q�t���2��l��Mv.�W]u��uϝ���d�e�0�4b�	2(#f��,MC�OHW3
F���O��i�`�
	�F�EK�J,Z~��v�W{5"���>�D�(-ѿ�S��9�&�0���]M�0�ߗ�l���O�������s�,�6F�������1\���ta^ ��|N���wj��2n4F�|�@��5:�2�8���z��o!�6P������� ���8N�K������v���SK?�8uk��,۠��d0Ɛ��j�br$��)I��m��:LU�h�/��M��EK?f�����i��rt▬�ۥh��`���֟�=��,0���5��uFP�-���Z�#`
�K�7aЎ1���w��:�b�_�bq��	�=h�t�R}��K��"m)y&u��5F��No�r�3_���ɩ��Be�H����5����k��QݚF�Y���>	���a���g^����k��!�+��/S����=�g�yS����g����g�v#�K�,�|4ϝ?k=h����`�G����+�;��!`|���E�2B��P<������i4����Vb}�vF��w��rf:�@Z:z�h�^��`�����f�A�/,F��S:)��;jUY�U��\��v�3؂�%!r<�Ɯ��u�cʤ|�+���<�ٱ�t�͝1�r���h�� U��fY%!���`�R���5�ǉSYWc�wE��ԑ�c���`zfx��s L=�,X�l��v��]�m�iV�(�F���m>�Q�o? F��X�A�b�H�22-�C���	�+��P�m�}%�d^+����<f{�ֳ�Xغi��Y��V�RT��0	�I� `k��� #i*��^I���	��a�%�N��PU���[�U:�j:�u�ƍ��������Fݵ^��4���#�b�� Ƭ-��ʯ���ޖ�Xn�$�=����Oگo��]��욷\KcC��u�-���w�T��e ��OF��W"ޕ��3�Ցb�����s���R�~��D�g>B�^��4���1?*�j�st����O>��Il:����w��F)�%a��L��={l��B�Eg8�>DC��H@֊�ln� X~n�<��#{�(5Ʋ� �-_8�����Z�DkD�/-��F���3 k���LJ�T���t��7�!�GB@���Syy(�BI���T;�KLr2�A"�hTsD����/����W�m�Qe� �Eq)V<C�L"{~��J��	�g۽=������l�ؓEK�Ц�e�����ؿ�0h��	��jץ�؎�W�����q́�����o��Y\���U��t�)���+3T^58|�k���ô���z�EˬP�ygQ�$�&��*�Ze�M�ǘ��} �,.�ٴ���ف��tҜe�V�������p��6R~ d6���vn[Of��J�.Mڈ`xtp%;����C*5'���τjB᩿���	�O�t.`�fo�
�{���b�{��dBy��Wۼ�sِj���C��yR�qE)��{��I$ޤ���o��NZ���SY��7Z��12����gȾ������p��i"˝�J��I�g̜J��Z\e�)�H�)q<�$�['
���]�=�N ��w"H��^���/���� ���'L�Q8���Y1x9R+$T���?�#���ONz����_'l���TIz�0�%�E��Z#*�ʪ��)�Y����c���Nb(C���+
�.(��O&.���R�W�pT�E3��o�.����~Ձ��ȥ\���}ՠ9�cI,k<e�nͨ�":����"��P�2R�� ��P���t��R����A�+"Bc#v���)�.�U�=d� V��G\��������G?�awt���U2�YCC3l�t+�ٿ��gl#���[o&��C���l�Jw�y��}�9V	h������+��#ۥ �R���ؾu�m�Āq@�J��mB������wڴ��������}��|�m�>�k~������vժ�)_Ͱ3atP��P,�M7���͛6{�m���C<�ԁt5V�Z����o����Ĭ�%����n��V�(��s�?��[�}���s�\Զ�s�Չ���w��X��X,���h�`ۤ׊F�"�<@�;GS6��P��%��r�&����U���^��ʺ_��Wa���J��^���m��픀�1aP̥8�y��T�*�Q�LCQC�l񢹀�t��>�1�r��[���f46��m?��:�f+R���FI��A/�E�`�y"sm���$��j;�]��>���UTcZ ۱0|���43H�椴�X;��j{w�`s�W9��tF{%�܎��ˤlV���yU�?-0]�7�nC#��>�ۺ���#@s��^F��4�H��Lr��P�N�B0�LE�Dc��VG �j��%��;\�td�3�ְ�8=�&�ـ������8��W~u�����	J�&�4þT�^gϲ���1�5�M��%�g�;p�m*���l�B�RG�5�0�����$�Sa�Hh�<�f�50B�{�E|��R)�����������ڨ�=�ÉDu�ym�â�|���t1g"VI����|�J�	_�Āh����R��_����F�f
c4�X$CdO:;�Hӏl��lPv�#c�T��6� ������A��%qpT}��R�0 �<����f�0�� �KvX\2�}�w�r�Vw����	�P���̰���$�4A������b,H'%�XQ;��Uv��y9�[��@�YU�ՙ�6� e��c�HU�aD��P�W�c��0틾�E(4B�D ��59�T�O��x���������.2�6ڛ]����Z+m���y�1��|f���Զa+��jv���ϛ:�2ʧ3� @�$ �f�Ə�պۀF|���v��Lyp�DU,��T��e@W���d�̲�&d%�/���`?�Ú�p��x'�k�s'�8�Ǚ���֩�$$[!�֍5CZ	�������pi��s
,:<^ӗ���":��Az0_--F�@S��T ��85�'�z��E�q~�Y?�;������{,������C;��U�Q.�?�H����٢i��ko�� @�f��`F"�:T�՜9J4�]�p�u�:#[:���O&a�<�4���@�w�o��}G`z�1k��b1/%�a�KFH�Tv��������-���aC���SŅ^2�a�c�n6֨f�i�r��h��h�s+;�l�|�Z���c�EP��<�]ϼ'�/hn"v���X�0�E��K'�D�z>�P;3����g�MCc������+_�����9z�.+�qs�t����"�2a�v���B�4ʟڻ��&�u�44N&�q����c��d���(p�i8꣚�i:��YGr9�z��u#X��.��Xb�8]�(�,��������:�a}��^����S	�A�R�;���]~��8�S���D&��ċ��h:�8t���h��)U��"�Ɔb��� � �"(�Er��������M�A��x��bV(ck4��u�1Iٔi/����r{|�3.(�C'��V�c�8�r�/<z���s���f���7��NLzW�m7�l��Ey�ʥ���}�YHM$��\��9�!���K�4j��h�n\�c^�E�Y��)Sj�6�P�H�1����O}֛��2E2 b��*����~e�~�������>�O�4�t?�ٛH�=s%g`�z�_�)>K�LY� �X^i�,��g/��.��j�J�0�sF5�[9��2;y�a��@�fOf���~���\y�$W+�^o�veύZ>ݿ}��;���	�Y��I<b�%�^��HP`�s�kN��Y%���8�q��Bm�XBy�i�VB̐; �K���:�1���H�ȓٳ��ƕ5�Vu�����[����h�)Uv�@��&�z	�J�G��D_YYIb<p��G*��5R��õ�Cuq!X����-(P�$2��z����u�W�b-͐4�Fqؓ;�(T�������C� �?��C��16H4�J�'֯[M�{��L���wYe�t2b-� �`)v����i^i�����{�����sv�قE��ND��2�T��� �R�KUŸ́;Nb��Rۖ���d� �#��G�資���,���&��(XI�t�+4b&|�N���q<���-:�u�0֢���}ǭdT|�I�r"F�#ci��v��lBuT�.��FK�Bf4B�&=;߲(��<�h�n����
�)hO�ό�d�g�����Q�ᓄ�.A�[�x5S�Y�m���P �i��<a��o`C��C���_�o� �sv&2Ԕ"`�~b���|�~��^�+��y��}W��0YS*�����к���LJ�y���>���9���o(���\��
��ӽ'�(=[�Ie��?��]n8h�R����!���~y��+`~��k��4O�d��;��ٴ�'��;���];m��md̹t��f�31�A�  c*��e�"�u�dk~��F���)2�I��gO���xn:��=.PN$�H�u�ҘS��o}��X����s͕�a1^ZO<�4z��X`��g�F����@;?�g!�E��o����Q=mL��l��~&�u;&akq��z>2��I�o�D��������3H$�){�[̠���V=�]��t&������^��#)؋N�@�@��$��Bu&��RIV�������avż����ϯ	�%K4�$3�7�qfܳG{�d
�Β��+>��~&r�rKmf��x�>[����j�l:�t�=9&�*��R�# �- �]̞�BJr@��{)�{���{�}�^ �?�� �=�%������T!�{-0K��
#qo�*�s�$�yj���R��-���vꩧ lSm�ޝ��4+�ȷ�Iɬ��5�}��쫯o�D�0��x�Za�NB������v�y�t��<�<��?P��l��0{�9���I�d��t���l���������Տ��{0ƞJ�� �0u����ûl�Ք�l:HN9��i�%#�߾�5�b;7����r(C�sJ�A:�.@_��������F�Q��Y,� %��>�ieq�7C4R�.�+8���%AJI���h�d�Ғ�Qc�(열^�tn�!��`���n����gL{]�[�U��m��X[�����l��J�M�m<�HݿϭY�޳�\��р��<V�F�����a���wdTb���7p^��K|	C��SYY�i͚�vvuf���E&(�K�����Ԏ5�q*s̚l��LP��Ț�`R����-Ÿ�h�*I�M6��a�8��@��X�Y��	�*�d��ȓ�Y2y%A!� L���V=��}�kߴ��u�}�7��g� P5����������Xe�8 GQΌ��nh'�&+eqS;���iR�2�\p�q�WJ���| o7�{���3��SF5�4�p��R�5	ک����IZ��1�?��q�D�N�#A�l6�$����H�2�0�W��#�(%��%�㓖����]*����.u�#�4ʡp� ��=BX�L:��͚SDwL>��,��I��&���Ū\PF�kh��qὄ�3�Z��3�b��af����XYz(�R�`g���x���o����2��������U0�'�h*X��b�M]�*���i���`��0-@��%f�E���r����G����� ��n/i.�1&�9�1]�|�bb�m�w�a��*��Oz{��Kv�VVTfw���5���q�����zG��@}���8	�*�&ɛ�=q �q�~eo�\�a�z8�4�H#u�O>��SyM� �MQҩg��SI/̌��J���+��rK'�Ksu�a��e��&��;�S[��z=������J����uT�ݭj�Ƃ@פ�Vl��I�~vPk�]�0�����]��J\�w]�~F��3*)��m~鵂?�7�]��3Dpi�t�����EQ���a^�'�9Bl�y�?���f�;N�����4�j1uh�`�Fi����⑜{�� I��,y
�z�8p�Y+}�5/�D@r���z�_����t�ڹ\��ڶ�֯�`3��yV�"ma<P�몫��=�����\��n5�ri��F�{��������|a�eP(ih��T��h���@����g)0e#��,P�_|�uõ4/Ͷv:�y�1��%���m�J��i�Ls>� l��,��W7brJ��cㆭ�F�o_�k��t�r:V�ڃ=���p���5_v*���������?nE��>�Qc�� h��Du�E6H�:����n<0�'Afhb��#upk�,�Q�1Ja�R(�WM��F8��E�xUv���~i��+��}������o���t�n�T�\W0y"{��j��݈�m�������KX�<7�Xo����+l鲅����	�<�[��d��}w�n���͵�UN���s<!do��I����7��E���-��?uB��3-�(��dr�d�4�!��	p�����@���.�8,K� ��:�� W-��PѢY%�L�[j�yϕhX5Y'����uT���(��8�ڶ�"��I!�e�},-��P�w�u�-��[?��݂�a/AO�i�N�����W�a�=��S,���Z���eM��\g
"�NLNSa�o)�Ђ�@t���t����{ޙ�r�bͼ��H*�K����l^�|�1�sb��yȵ������,$�6Z#�����CV6��u*-�ǧ۪'���Fc ���~:8�I��Lqf���$;������S�P ���.�Xđ�`��t7hT4��%!�8���x]�~��¯�u^�o����)p�k9N� ��&���� ��p�k�� ��_���S��I��?��P�����:X]�O�T���^,h�|_��AÚ����#�����P�Kg�y������|?������0���L9
�A��M9����M&{��/���9�
J�qG�2�ih���}�6�}ե�ol����������d�X02��%��Z��h��9
��W毑fcн�*��6u��s강���d;%�����L E`E��X?�!غb�t I��d�xң{�{/`�%��*eʝ�����5ivrwpi��L$��`n�?|t`���Ө�'����W�G�P	A)�̰e�֝ q ΅{�0�q�4q-��j��}�{���kmk	��vL�� K�ߡ�أ�UL��'s�(���<��H��s`G�o20��̵�B�
dhKi+��B uT�mٴ�2�4:0���� )�nI��|!70z��K&��w��
��-_n��݃D�"���/�5���T 	��_e���.�k�a*��S�v�M�yBC�Y�퀱�g�m?���ط��m�(X4=o=�`ҋ�/&�po4�C�_2�VO����T���X��Q�~�gl��F �6@�x�uR�en�tO~���j���.�����;I6R?��� Pyv�mV:�b*�v�ϐG~���YDȧ�C�u�.�?$�}���ln &�s�{`��)W�#�"I &$�s�g�I5���Y�ҵt�vS���/��O�v�2�II�|�~z������4�ߗ2�rTC�9��պ�y�g���&f}r�M�a��u>��S�LM7�E��vcĘZ&2J1	|NM��PB�M��UW]�{�w�%te*����.���7sd��0�&q���?_���@�+d���	�O�^&���)cM͍��ELiqqd:�k@���	���_��f��tF}�ѕ��}og$N�=��c��OBYSJ#��Y�{��^�8w�S'&S�Z	zCvꊥ,�ݐn-C�O���	�JJE#VX��k��h�"������.+����r6q�2>��,�<���� ���:�Z�^��X������s�TC�Eo�Tx�0h�� )��2��x!M���h���K�^G̓,Dz�i��R��CH6q���ΝV6w���mcN�O�R����,�$��!�f&A(���5?�L'��tD�
;��{1��k�����h&�+��X�8���žs����#&-��MZN�|��u��p�/u�q�H��]�!߰�(_o���`��:��~���e�,�#MԀ�I?�@���}�?��]��B�G暩(/+uG]s�[�Y��D��X$����;#Q�4_���q�W7x�Et4�M�v:�������:�9H�Ӱ�I̴}G���n�4���pxEx��bQf��Bg4�y���X��.=����"�J	��@%p���=�H�`�# �E�K�dP-�%Й�9�������&�S^>��,VMLV�'N%_�5/��Zz�����$����?��Uτ�Ke
͵��C$����5�SN�ز ��9���q	ϒ�	+�`i�4���CkW��z]�� �� i6�E�V9��"���#��쪣9�1>��E��놦���c�����K���JT�h��a�sN.�lĐ���6{�?f��d���~zn?����C��Bl3�)Ge�����J�`�@���{]ɼ�wґ=���Ɨ��u�ća����Doxʲe���ØM���~�a���C�@���b��ַ}0���L����� ����ҺP��d#�,׮{��m�ŗ`ɂf ���k��᠈���$��t�T��n�����Y(+`���!j�Rl�\b[q�e��L{�5Hzv3N	�44������?B\�A'6څ�<6Bمxy� � u����q�[q ���.���}�`/l��5�Xݾ��nFP}�!��z�VJ�a3�s	t�>�(��g��L��	�����R�ҳ@�|%��ed����}9/��2�=gr�}>k�|<�V[��o����n�Ѯ�z�/ȴ�(_�ДE�U����3��>���6J�i�xM�$ʩ?�3.33m]��lo�?�<�:uj�ܹs�ܼyS;z��P&gڇ$�)�F��"b��1%sɒ%�����S��X�ޞ�[p2sߣ,%�r]���xm�d	ȏ=�2�^�Y��$<F �&��K16���t��1���wGЋ,Y<������w�!��O	���7Y�%\>i�L,,.%�!@d�P�.�s�����i�^G��L-~�\������@	�v�@����W�i�(�* a4m5g�XuM��8U6iM�>*�3�Cݡ��o�c��A�,�n4�3}xA�ZI�OW+#P2 MI�ki/��,[J-����)�
(oFh$�U0�i� �`���:&�#�xU<,����K��(A*�hJf�%�}�8���7����,�%&����������/������*y#�/?�e��
3�6T�qA���;&{�����G�OI�ˏQ��{�nsȅ��tU>^OH�D̮�����t8�����V�������@J5ߗ���a�mcƋ���" �Vhͣ�X����$v�2lX��s�[b��/�Զ��� l?ݶ�{e���%�W&ԏ�]@&FFB��X�_�y�QU{�Sk:ݙf���Ҋ��ϗ�� �C�u�?}}Op/���)J���b����~Vf�o�$���z�I�V���|�b���H�'p�À�+}�ط���C���.I�V�K�9�`zЕ��9�.u�=�g�F�(��,ZL �K�K�$:H��+>	���<����l+��|��1���u��;#��|<^F�{�#)�<*)Ǉ���R�������1
.a;���ٔ�
�D���E<Ӫ�
�S��m)GsCS(����9V�S��g6o�blC��0�یnt���r�b��jh��ΙmWRz�D�l���Z��K_r�� �Ϟ��J�B���#�?�3�O�$e�ALP�PBc<�����{��u��=��� �A,؇�Fv�����m�l�ιuɥT� ���(8cF�7��9"*�=4'`?[�[5��X��7"֏c���qεQ�ɰ��}L�m�}�����rz����I�L�䀸>$��=���s�>�Χd�N�� 1�\�im��@��m֪�V݆2U��Z�3�7��Ө�1~�����{���ϳEK�SP�� J�.8�<L�K�xڌ�F&��d�Z ���N=�T{��u!��6X��ߩ<����e�w.1��(vxU&���̢V@��G��g��fӍT��6I]�y�b����� �!�D/�ƌ�MdU	d� ��8c)�@O H�F,G��b�̙K�y�*�H9G����0��t���*��Rj��dâ�S�:2ș}�:^����}14��41�7��RiٳR��D6�x�ʺ��lգ��ٗ\�,�9��;���l�;n��.��B6m�=��Y��w~b{v�Ct	�Q�=�{���[6n��\2>S"�j��\�<~��(��@VAV�))���S^H߫|+&L F�-�<�v#D{�����C���6�i�}0� �?��]��^泥r�`1z��J����h�z�Ev#�����y�=�v��ߴ���I�#A��{9���X��K�[������B\O��Zڸ�5�M܁�����c?Z���#�GaC�y��G�� �L"����P��M�����%X"�4z��U@s�A%!+=G����L(�P4�VQ����坏!�NkS P���x/��\E�!x�qA���ϨQ�/���(��rA�W*;�	��]����WK�T1�O �)��� i��w\ƛ u���Og��˽� �M��d4յm6�0�j�%s�W��j ]V_��"�C���1bl�X��=��	�:Ŗ�'�>`F,�D/?��|�����B��$"z&L��;eW!=�J�)��p���J��`{��01	��В�� ܞ�{|�w�D��Oc^���f�z�Y	Щ�Y��P�"U��Z�
^_ݦ��!�����Д y}�Ñޫ!�JYb��̆�sm>`%�� ��-B�7�`Ų>�{�w�G%JE]�D�a�m�fl�k�<`� ��N�QN�T�>I<���N�?iw��]��a�,us�{���G�le1�h�Ć�"�覒!Q��]hj8���l;�;�a�ZU�L�tu=��T��K/�%J�_��c��>|�N�A�f���!�؅��+�t�\2a�'[�&���:�n��f�/�Md�50$<�D?�8/��و����4���j/#6�0E��DM����lF͞3�.��B���?������/��J�|�҈����D|��@�x7FS�ILK���K��tG��4if����I�cmւ�h��<��l�A1�w����Ⳋm��Sl���[�/���7�5�gN�}ܾa5F�v���n?�;��"ڰ����9ȯyNr��ǟ]�\e�eĒ؋ڧI�;J��(.��0T�m-�l�9X��s��<���Q:��d}Xo��Kf��������&�zڛ�5<lLX+�$"�&��g�������Z�=�~�=�݋��4�S��tvs��CC~<��q����^փ���ܧ�x�sJ���Q)E�f�d;���{������B�|5� ͕f����x�r*�&Z}��Ne��K�J��>��� � �6>}Tad�z� _��4ۑ��	��Y����s+Z&زSfU��9�0Q���Z��ܣ	�('��ȁ�ۚ&[�z-�6%o*PQ��$���\����6$���A�o�y����s���M�
� �+�E;*�V���ʗ�$�4�HG$�A�*jY&��[s��*4���ҁ�ț�B&���,%,V�����z
v�t��m��Oyx�(�ά�����*�,���(vo㥸wi���E��'X8�g��ˣ�=m��z������.�� �D�=h|Z��{���,�%��������L�,�A'/
Q�`�ɆD�@��CC�V��~.��~	X��%N��e�z��*��v�,^����~���Zp Π�b%Y�b����@G��i�^������B���2b��sG�}=Y����]��ӰKPp;������@�0v2A�@��!.+���?S���6�CG`E~x��S滰��u	�e��ÛsF:�*���e߫@��,�S"��ݚhOn�e%����T�k��ѣ���r��+���Q�%Wت����w�C���yV�eD&:�>��0&$qC��82}=/u=�'L��F�TVU�4F��~�J�ҡ���z���w�w�tVl�>��@��]���$��>}&c���O�:�ý�**-� �òSN�Ĳ�uWZU��Ѹ"�.�e)c�J�Z�ӦQ��<?�K A P@�-�b,�ĤM��O�?�͜9�Y9	��t%Q�*-�>� �`q�]�HX�YVY1�3თխ�C�@#��x��W2-R1���ISC�`��p.#Mn���x�Ф��t�^��z�]$�5v�{�eG��!��Ih]S��5z�����N܊���L#���I��M�l�杶e�AJ���{�� Vs�,�D�ZF�]ğ/b��I�M@��rt�9�g�XؖC���#�v�ށMBk�~�}�{�w3P1����a#"@l��-�uU<�����G�N��[9�"�؋��\�$�,�R�p_�]{�[Y�}�Q�x��(Қ:�#N[~�]~Յ���T(3����kv3)!�>��w�D��l>d՜K�Ҟ�j�Y�MV`�%�l�@��VM'��9#�kш��;�9�m%L<I@�)��y��Ώ��������o�ΞǟN�c*��9��f�o���|X����36=�
a1'X�mg=�8��芎J��KO�{J�m�l^��K�gP�O�堗���c�d �NEA%cX��OZ��63���qqQ�A&��?$.�rk�����2B#`��ׯA�q���V�ܹ���Q��&�T�խ�TY��ߔT�1���E{���R4[$J_�a%���0^���a����a�y�!��WC�U�0���cي"X �NAz�e�B�g��x��}8bѕ���y�ć?����� �s.��n��v{��'��6&9O��	8Vs� ��H��(��t&��^��T�a�&��if���-�%U0R���f
�?t�ڼ���)I#;++-p���x�Z*3������)���&��3)Ф�N�����o���.K����68���6nc�0Hڔ�ND�񘨖�S]/�E�c�ܹF̖�[F�\3�auE ����lھ�	��K.d<U��7��X�|����w9���u��ap(p9����i?�B%�0�
�����s�/!{ ��H�$�|�-�5�V��i�T��� /ߨ��;��t�x/�҄	�xI��r��;�j��O0�A���Z�'`���g!��׍;���Wl$@q4��k
�7��ȭg,�����x�[]�iC�~ysI'A����?v�!�?u����U�����W-�fX�t��{���%�t&���ع�y�@��7�C;sG)�H��1([y;
�I���r�t�������X���y�#aX�p��ga��y�b��m%р�b Z��4��*0<��8ү��do�"�h xAA6�S��Mڹ\����Q���N�}�%+����s*�������
�g��.�k)a���	�f3���3ϴ��9&7o�<b��,v���н�~����1k2��ܐV�M�����l���t�=�K�9��b\�����C|�)�1H=ߪt3�[gLĮ��K1�*ʷ�g�_�$a��z% pՈtc/ګk.9�V?v'�v����P�\��?M�HM֐�ty�����Vy
�z%e� =����x�Q7��8�ܦ@єc#���s�͵�wGa��������W�Q1�13U�����f�	K�l�milĥ���tX>�l����-Z���{�CM`{�����g�Wo���Hi���/7�95H�~�5��4Ð�mY) q�%�x��K���8�������J*���C��([�hݰ}�?�-[���^���k||�Kr:`�{a��`����I%0M�]�����D��1k�[j��Ts�w���>���b:�`��Y��r��s�zC�^�����d�^�(!ى���l����뷼@7,�"a��C�F�עٜ��m�z|�#d�q,{?�#���6�X��4���h�y�9�G����8��0>b�N;���
��lU�en��NaW���	�SAh�(F4�ee�ODG����@b�8���AN��Y1Y��21��mq�C��'Ws��?�Û7�n$���@�0���Q��K�B����"`�����r�S� ���E�^H�:g�(y��&�.�,�[6n�iU���w]@fB)LP��e��M��Z�Y����{�z�)�6|Z��x(�M����R���j�Ċp���jގ�����S�:�8Ą���N>�c�ۻ��r̖�z���**ěH%iՔYi��X/��i�� �
M�m�����%`�"i��f�P�G�1�L�bM�^�;--�lߦ�.{�M7��k|��������D~��~@ $��-��x�/�ԉ�َ��t�D�r�n�E��7h�-I�C*ƙ/q>�ʪ�H���/�B�Q�l=�PX� Ћ�� �}x���h��@{���v���݁�}i�g�$�z��¢lP/���w9t�w�uS�B�i�0"����%��H/�r�D PT�T	"x*��(d�gb��F�p�S̑����A��a��j̈́�m��"���$.jp��Sl@�Dk4�r�7�������9j
a���Ջ�}�Ƶ�췷���Y��x��'iJ�D�J�ٗ��&1��2Gd� m" A Q�0�G�gv�p�7��۰+�v�~_����cO��TiQ]�����m��2���w�~�����PJ��y�Y���<���]G)	�N8��1�J�Q �����gO�]����V=I��[������튅QS	S�6l���Q�e�����ˁ]��[/�&vtj�t[�탥;D�����v�>��@n��)O�5vzol<�c�Mh��M){�f�Qt��}'L�Zp4�
�U�5yӑ�5L?I�=���(�F;��Y��(���$��k圓9p7ڝ���5���G,�Ȗ�wrR�5�1;�̎�#�q:e_O^y�jb�y�s���y��k���g���y�lk��R!?/;�@��0�wmR-��|R��������q]yc%����N��H����s�i8���ᜳ/t���Q�� ���a�j*l����+K�@���>b$�>l���g�g/`OD�c��J���ڔ�D:Ks�
���S�ŗ\k���CX?h9��-�X_�h���)l6ֺJh����rO����fb{��{��YF��-�?:��O��0i���Z�a��%b]��&u$*�⌋$�Od-w�y&-���f�v��VX��[�r��/�[�Y-�O>R�:�s`L�)+�%1As4U�S���	�T9����ˋ�Ħ��~�L*�b'�?���%�ѣ�M]�ٙ5Gjk�f��I� H� �����9t,�D/٪��(nZNP(�k\������":a��JH��É�'hm�ڹf^�!(��������SB�
�	���A���ņ�.��Z��d!:2qt!l�Y:P�ZNƺd�B۰�(46� 80q����_��-e�r��X��cr�N$�'G�ƈ�8 ��)i��Ԉ�C�b`N�q��f��ٍ��WYt&�\	���7۶��^j��q�3�m���;�,+%��ƫfB^k�$�T�1� ؃t��A#�r�X3���yt*�jP�ʞd~�3�6m�Z�Ϸ�4yبT�j ��~,��C�W���3j�w^{���r6(|-ϢE��_~Rd?�
�<�ݳ謑�n}�8]�W���C)W�I�N�j��ݲ=mʡ�����&)��[� X��/̆���џ��� $|-��Ds�jyW9RAw��u^z�)��7�TK{�CRm��r����K@A H�y��������8s��u�]��SO1�-��`_;art�UB��{P SL��J�xT��L�`F�XL�yT�:�p���ʪd]������Yh�" �*�'Й���� �:��}`��yz^��?b_��O�}�_f�)ۥ� ���:%}�Ct<�`_����g��X`��1�񹉐tT�}0�T ���wd����:�	��G8{���Yk[ V�>������8��[�]��s���ןuu��@jԎ���z�#�s��HK#�K/f��籑�P�b!I��~:'�F���{C�O�- �k�����A�	�]��WL����wlw�LC�e���.i�w�Z�sT/0�=�����U�P���	qIrL� %�qp����<�. �Rv
�E�B�/2�>�w���.X������I�SQ~����öy[5��]68��6 ��M7G12���X�����a�ᚫ��y�����\�k��*	+��|u9����@���ί�g\_�-���X�E�T�;*���iUn��u-�r3�����d:[_��n  �F���̫�|��8xmMۖ12k_��&�S�[{x?C��37��!�V��e1��>,-����b��g��=m�G��`e�2��Oז����=w�V��B��#HG��a�`Te�3F5&J����`vdf�I3��u��,�V�i��ͼF�|F���߱˻@�c^[���5�^�mG�/h�C�JSOdg!K���y��s��ǉ�9X��8x��k�8����d#�	G���hM(�ސlc���EC�a	t��K?���^��Z7�޵�f��Tk���*+�X#��F�_����_V9��;��7w���<�h {zU�h\�H�#�A��!YĢ�Eu��A�d)v(A����m���^:&ܻ&<��]�)q�E�fE5k:x8t�`u� \	i��d�Xw���&�O0k�A�g)�#A�<���3��2�Er����e�o�e]�;"�ى��I��E���g%�	�Ǣx#��fCE�!$��� #�o�4b��i�_C��E�Y"@&�L _�՚5�a���.9*zL���|��CǗʗ�(^Ә�7F�3�X�h����3I$K3ې���5��p?���<��	>�g�Kf{�?H�٘�>�:ݼqA)��8;��3px���i<�g]�a�����'d����9{Gi��}�򫮱/����c��M6���A^�gt�?�1@��h�/!7D�N\Sa[���]�r�/l���?e��͔ÕB�B��bWP��J��NGo�5!���5����T�� �������N[���->�^��T�EC�up� ��PN��5�!$ �~�bm'�@�
�G���J��9�^�B�v�>^��qg�=<cS�U�� JN�T1�Ca���EGZ�7vM�ƒ���_��,z���k0Rϯ.��Jf��- D��1o��*[�$�;9�8������H�$�����;F�CS'�|��ҡD�'���A�X�`: �{Z�@}��B�� )��I	������/R�7Tf@ (+V��K��`%�~b{51H��?���3{�=�f-Ic�xv�Y��d~���n�Tz���B:�Tb3�ŭ�Ͻ�lլ�>cQ�� J R9 ������/)��t��+0��������X����xd�{+�|u?�
 p2\ )`ͥ�*/͵���sX����|tTtt&�+�"��V2�;�q^����!��0�#�e-̜Zn��:���}��=o:�-o���?VF�0+����>k�şw��5����6&!�dehL�(�^>@�%�������F�E�}�_�ht7��J�����"4:��Dy6��e���*	�� ��d�X~�,�-^��<�%���}��S�d"[�)8�ggڞ�� c�VJe�w���(�D����� F��ꦆ�)bI�I�m݆=>>^S[��7Fp�;e�m�y����I$�F��_Y��8�J+{e�)���ML4�y�C>�QM�Y+�����Gƭ=$k9��|X�qʹ��H�V���!FY�}��?�ů��%@vVw����h��s�&Y���G�0�+ E��Y�Q4a��I��ڣ���*;��� eS���nc �W^y����w���f"C����A|�G������"Ɯ���K��^�a}��ښ��d���6u�4wl����3Zܱ��hL�D�be���X�q�1�#�Z2�������P���Q\�Yp�d��P�����LG�Dhhi��~�6�CK2�^ؾ������0�������ӟ��w%�ʨ��ÔF`TI1A��J�1@�"�8Dwa@%�$ď1dBüN�@�"(kQ�%\�|��( ����*��mPP�.4�B�������.��>�q�\?��N%6S�Mqa�Z��&z�<4��;W���������h�����فdI	e�}V5c:�4CiM��6��R�3e��ұ��0������q�㷷T9��Q7cz�-b�o
����x���LGc� =��PL�U׵��~�;��E�RN����6K+DC�# ��0ݔ��w��r���̯���y��kZr����8���G?
ʌ)�k������_��>�x^"*�(Ix��ĺ��~)W�Z���g����t]i����8o�1��?4/ I�|?BY���x��x�]��B�	��hnWA�� � %t��	��r@*�H���A�b����g��5ir�(ݏ�a���j�n�h�X���3@&�1���A�H���8Ȇ"��+z�$��U,�@�؟�S���g��NSsPžd�i���ُާ��������|u���o���i�᥍����^��t�)�q1sA�]�Li���}�Ao)��)j}��@bZ[���vuvs\e|��P��:�4橛u&V S��׾����;]C�� �m��j�<���RǪ��:�3�k��x�?�
��
��p�Kk�,o�uRW~����~wU�Vđ�*	*�N��A�J��͌�.p�?���&��N^gLՒČ8��j�9tZ2�(�3����y3�o��ďٷ�7^w��ݶQ3vA �Qio��r�Eܷ	{��'Q[�T1=]=�����=<s "�i����k�u��6���;����~�0{�C��D��봮�By�ۗ0l5/l���R����½�9$�f̚g=�_�X���ks�h���=��:ر$�t_v��)�������c6'�~�3A��4A��ܒ�(���m{{
/�<�6!S\ @� µ�-
��JwhS���B+���e���p�/��n;�k�>�#�:9g%uQ�n�-�R����3:0v�p��![O����X�Z���u/�p_�at~h^�}bFe�|���h�:Tc�*C��>b�d#��8lfF�O�4�ţ�_�~���.w��~~� p+I��B�t�0b6���3wp ������Ǆ��)��s�)�L�]uM���{��8�9cw0⢕�ص	}>ȗ̊-�,-�GY`<�z�N���U3A��?���D���7YR?��	��X�I�h����j�JL����hL��Z���<��fZ�̅d,�	 �P���X<*�d�����jRP�G�I3^-�dۃ��v�~y	�����ŢC�
]�����K�6ye�� �ttj1,$�����B�ya;��[���a]K��s��?��Z^��� ��2��n���0fEq%��9,Y�O�L�1��$oD�C��H�L,���-�������ٸ�V=��
�d�5��3m����g����=�R�,���4��}.�T��K�;��C���Ǫ���`Za7��Q���Yte�[##7�3��u\�L�"�[n1�LGU
`������%��Ɇ�"����5�^���9��Yg��:t��ut��{"����#�_�ʃ�ygd^g9CX�t�������Ϙ9�[鐤�&&�f�z$��Y�\�3E�x��^r� �e�01!�3
� 	p��O��F�B��H ز�^IA4����C��8�#���>�~Xe&��d�cP
�$@b���F^_���O�� �!iIc`�[���(H .CV�!g�$Rv�sk�ڸ+J?H�|�����4b	@)Q���yV	�Me?ϫ����"]�\��N/ѳ��Gk�0僤1;�^|��`��)��"a�bϋ�ΤS1�� �fL�L ����b9�4$Z� $���%�.P1�Jb���h.�?)��i ����� W�N���$\g�cP����(fh����s��4 �(=�:�e��ε	l
�BL!�&��d�_�1�0���;�i��6�7S�D���c�z{Z���!�~�2ε1�ha��J�f�� �:�З))�a�$ ��3%�xn!>�F��ݹ�m��̰-������J|�9�T�ݗ-�j��*G����Bt]*�j���T{0;=��W�c��e$�s� �h�/l�j[�uQ{�4qz^c]���#P�GQ)c�z�	c6����L|$��	��a3�À�C��Фt�O
���X)�/E��k���8�jC9�}�y�`���:�W��5Po]~���i` �LF��1Mf��uHc"I~���O!�xI&_��1�Q^�.k�3��-�ZJ�-t�ǡ�N"�nx�D)�<�,M�4�܏N���'�3���������F�4<̢9�2�`w2ߙRj!����]6���}���*ثAH�!bHN�aY�����Q_�JL�i����Ȱ��{�U�zF�q�%�^C3� �gb��s�s�c�s[}�HQnV_Frb?V�/��)��u��_Ą�'��6�'P^�+��q
G�]v�i��ڷ�`?g�`�(�h�l��1?9�g)�Z�i�	���hȉtQ����R+s�v<�ͱdw�.0 � #�g����{k�k�o�#sb�$��@hچ�<.!�NZ|��{�>2#� �v���,��n�6�"e���ѓ��%��J��<�C�7�4>Gّ��&���`"y�cuF��a�2���0�h@gG�ed�a�Fb`Ӳ���.�9��������h)�f�}�:���s��f^٩Ϣ��W���3�<�F��ol9l�O�s'w:�3��𹖞:�~�??(ؾ[����o��þ	9�z�-�U��A(b�����ZIDsgUY�C��D���F/V2����&ԣ98D�&V�Z��2 M)SJ�7��0
�Viz�8��8��|�T9�$��x�Kxl��wH�P��`t��d�)@�k�D��^��r0/*N��x���ke�������p�����䥥�&�`�g���e�bO� �b���&&D���&?�
��}t'�bs���E'��
��}܃^��3�b�� ���+�g�q�aS�1�]ұR`�� �(R�܈u"B��>��@�	 2��>ى�q ��� ]�� %^�^��}�KeP�a�G90?��Z�̫ʵ�0წ���b4&��9p7��l'����N���*O��Z���S�e�X,��a@Rd|�Q��ƥ�~������<�8���Ut��ټ��mϑ:L ��%��<��b�"B~_2}
�� Te���o�CZ4n�f.��ih��tn�n ײ���̘J軒nў�ėdD�Ě�)�&�W1���)s�Y@��	!�ܜ��m#������N)Т:���(�J9SHp�GY�Oa�:15!��K�rF�����F%	�B�֕5�g�i ��_�0��yx$�
�c㕰n����(Dc�J �I~��&��h����6�03�)���|���k���(���do�����Q�m���tN�`����Ρ�{���ib��{�qd�����Q���:����?CN��!D��t�-;y93'���iJ�\�_br��h3����u��ڇ?�1��SI0���1yH����1�6�kf��$<�E���6���.;�o¶n�	2���tΣ�c�\�Y����AW,�ȂYS��.�5o�-9u%c���ِ�`Ŕ�読�؏��u�k�c���B���y46S~���&�p�8�OǛk���6o��S�s~F��p�e����u���9<a������D�+1e�'�G�� @CEWk-c���.�Y3fzC�IKN���}�l���nI9T���a����ѽ=� �K��Cv9*}���8�/��|�S	��٦t���c{�G������@�nKKOO�DRvʏo�w������9fg�XaW^s�=��Z\�� I'SםL�"�;�!�r����a-m��B�KFf�	,�(���63�>���d�}Q<d1Tr��%��h�c$�2����t��M8l����l�ڢ1��*���~�m\_k;���f�$˜F���ut!e�Ӄ�B��|�M-�a�5�[4t_g���{i@�7gY)����v�4�1��(n��� 椢b��4Y4s|�T�%76�̫����:�ZYl�������f��û���V����'��I�Z�XP���Й2��M��aHS*����_��?�-��ӏ�e�N�C����17���_��	�Yu�M��� ZkO>�*g�e�l�qz��@#Grhw���������v���0[g?����8!�2��dӡ�Z�Z����Q~j罇�E2�?l�hU1Y�4�:��ގ'^G�}}x3oM���7h�K�/1?�S�Ke׀���1�`��^g"����v�.�ޯ+�o��g�%L�.�r�����x�`�iP�@�K� �����ff#���P%�x-O0�1�� f��#6>F�9=���Q
<�D�F`AdF<�����!HG1�1#���mae�akG���Fņ�˽���B̭�C�}�v$�׵�"����Q�#�I����V�;x21j��]i�����O����m�SmǾ�>�r���z�kݿ��5��?u�b��׼`�^�.�̯b$L;eh�8���5-֊�݆T�)�Q����WoeD�ɰrH`�v�J�є�pπian+vS�-��C���3�0A�ɡ��$@��/ز����F �c�yK���8��3�(�iy���'��5/�Xҙ�[��V5M2ب�F���t�S�o�� p���^۸u��=��zW�c�g'GM��&�����{n����;J�< 4������z�O!�
 k��ߧ�w���>�mb�����o�=�P���x�e+���E��K�q?k ���e��f:A�QW1m�+�%!�ý]$�>�����?�N�}m4lu�qaI!�6P�1a���׷س�k����VQ5��Z��d8=F��e�_l�sN���?�u�7Zy�lb�6[~���>I2y�=���v��ﱝ[v�oŞ"!��1	���ڧ�Y�[�A�����
�t#�  t6i
�Fu�~��otM4���m'"U�r�� ��n�G=g̱���Gu�w�͞|�)�m�s����6����S�t]Ո�W�;��Fz"��(�ƺa�W4�G
כ��Q"3�O�^f�h؎�p�w�hb�b��w�����і�}�'���0~o;��l<�!�E�� �p3�L��:��x.�ﳚkl��E�:	�8H|������@gL�C#@:�a�IO���U=����%3��*?ˊH�N>�t|:7Fk��/.�Hg��a�v襧�wg�16��*z��l������{{���v�{�E5���@�K�l@
���GS:�PVz�~tN*�D��Q�\�e���	��"��j����Sٸ��R�٩��N�NF!,^�zv�-�5m�5��,.�y��ڰi��8�yJ��5dW#��ު]�0��D���"�؊��ڪ�@:�Y0a��M��gA�kG��X�A�O\&s#� P�1z��������v��D��� 5P*��#N&���� ��t�t%�)���̾�1 ��X��t��q�v����2й5��]j;�v�I���Ճ(\Y;����˯~�K����?:A~	������ڃ���V�Z���:/���fR��%�! �����7�n�4$���u�9l{��H�4�t�\;��-��+.���:����]��ņ�œ�r�8�K�#}��P�Z��	�7�����Waa0vܼ��+4�j���:�28�ɀ�/�����:'��k�����w�}��)a�fDeO�{�D��i�0M�t���(mM��n`+�g{
`�ϾRv��8�q���#�RY4�C:��*�oB�[�ُ1���Cr薐�rJ<?!M~~ڗC��ty��L����@/���(#h�l�+?��/��;n�,:�����W�A�{�k����r|���8��j
�f��h��#>#�kmo�M���2m>��[����J+���n���������z�~�A��R�m���V���U�B���'?FךH�������n��RP>$����f�<�)MI���3#كp�G��߿��LE�_�5��/��54SU��Xk#��◿�1�R�.:5�~�[hð�!�]�u�mY�mS%�( �wcj� %C�����
J�4��i�'I,��V��aX|x��5����c-������a��1��!���<�D�CO~z 5���Mv���;=׉Ƶ��Z1&��w���n��m��9v筿C�^M2N��uh���sܔTɨ��}~5��Ҁ�N��J�b���|�#�����ec�z�-�7��\s2R]��Tw�G�M�@3��0���*���������R$����;/}������V�M?৏��LF����{��]��j�PR��N�r��9�9x͕SM�f�l�4��6�����:�k�jH��ܷ��)%��K�$5j�(��7�U��"�O6�l�9��S8Kc�䬁1�yZww��C�McL.z�)4��ڪ����Gm8�"�}Ҁ�t�J�����28+�؛�/)af%���Y�'��}[7��0TNd6�c�� ��U�H�a��IS(Kg��������a�*�D�޵c|ժU	W^{]eNa�Nna���&����0%�d%#W_|����R���l ���E%-�����L GW`�4ԥB �I� ��ZVc14\��l��c��9���	c� k<H���Xsi�x���f�/�N[��Tk�0����@8�k~v���� �"A��}�A� M�Ժ(s�cD�J���+̥�e���-�P�P&�#	<��6� %�n��d ~/�=����rI�De|�جCd��I"ДDk 7O�Z}���a���.����Q��B;e����|�c�7�a[����Lڑ��[�j.F'Q��K�9p*��=�i�f&�7��g�i��q�m}/6�p�KuV�C�rLLF����O0�����m;��d$��d�t���~B-�=d̙�hv�ҍ�4GhͿ��S�鷵�.tE�4[���(k��&G��f���^o��/ݛa 8�sb�%��O�ɬ^�5'����n�Wm2 �\N�ӯ�O�N]�|�d.�ʧL�nn2���.�~�d�#.�a�N&�J�^U��k4���H�%Cu�!�+��vS{�5;AR4
3+��x_HM�lS�Eq0,jXgm�cdI�.�D�� �54H�[åeC�C������T��|2H����OG�ܹ#9��������&�`�`)ץ�U�P*�.��}�>�����"V����(SB��Ĭ�����:a�F�Fa��y��k7~J�1w3`m�c-���x嗱,0�v���E�flټ&���=�\9�O+�A)��.���Y��ztD�H84[�����YK8�Ҁt��)_&�I�Se���F�P��\>�{�Q���OO'b��{��-,z�i�Ј8br$����A-4��;!��7y����rJջ��X�ʕ�tO&3�[�fq�9�'��^�o݈����R��uqY�Mtv��-��b�,Ύ	�ܿ��}�?�ȳ�h5���,��_��0���.����՞��ɛW��[�D����L���ї]v�uv
ՁX5`H�Fɺ��0��S�����ى7]������4|*�3~j��d=�*.:F��~����OSnw۠t�M�LdiB�XG���D]����H �&�H��+��	�M�f��sU>i��tP��%!�n����[�����.QG�d3j IN��M�2B'if:�,B��П��=�pΕ��\��L�������rh����.�V�eL�L�J�rC�����N�k���Y���9�;�����g�%���wn;��E�w���f�	�6��!!�А�4Ɛ*٬�F>w�&^�����}[���-i��S7H�� L��3�&��w����y+��_`�l��m�.;-z+���5]s�BB.�:H
���/o���sg΀^�C#[v֙��X�m�r�΢;��2t石�f���ۏ�l������j��)+�x;�w��c�2y��Ç��5��0AM�E˱G30�e��A����T2�Ҫx�`֨�M��*?u�uc�q��~XEDR��A�]i�>l�%�Ⴍ�)��,��]�繩AA��`��N����Ρcu��77?`���k^P	����P��6g!Yc���wc0+S������8�t���g�O0��,�"X���m�/�������7��EN�(��]�a�����}��5�0^5-<�K/��֬z؞Ƿ���[�v��_|�=�v��~�=�A��_��fΨ�UOm���X: ґ�����Ҟ
����>�h�:�T>��SH��r�؟^���k�X���]��^Ĕʝb¤%����ǲ��2G'Qn@�;3@ W�LFc�T�����ÐES~̊��H��HyXFa�*��("s�>�,j���{��F�I��J��e���@��d�Ǝ�b����J�^����#օ7R]�}\�<�0���Ac�� �8Y�!�s���Hj&�F���ٟX��X�Q	��s���Re
qD~R�)>b���>$�I[6��tt?�򯟂����Y��z�ۉM��_��~�����t��xb��=oCR!�rd:���_��/�)!&hD��ey����:�Q�	��_�H#�eK����>o�ad����$G��
c�Y��挄	����4�(�$�j)�FR���@�!V�"5v�[2!� ��!M �*�����w�zW��%�e�O���DQr��HɗX.y&&HdA"�����6t�;Hx���Q92�x߄'؏�[ۉW���SR®F���>��!����+����њ�3�}H/`h���3Vش�27n]�d).������
��˖.�lVs��WX�d&����X�a�;��3X���7��4�<��sv�=baQ�F�}Ľ8ؿ��r�,:;��bL�u�{}��,|�2��ϧ�o2)������	 ���$*@�j�6E�qҏɂ��8*mV�b��*`�I�v�Y�L*�]U��`�yF�'�ٵsmh��� �!*I~��ƫ���zI�Հ��}�J������f���t{~�N~0_���K��kf�q��.Mt]�\�%�~X�xb�J����9��$�	����²��Sx64���l���2���#0�o毿�uv���Q^�q�Nȓ���:{�C]]�=��[��^�O$�q+#g�፣�`�z���v2��?��J(:�}��1�A>g�,��w���L��`�����K��O��Cdwz��MH�`F�?��Y�c8HS�n�c�f<�2�U�����QZ��)���#$�ҡ�����ʨ�6�ʟ툂Sb��XՁ��FMc��A�	IP�=�{#znN�ã�#�P�ݍcv�� �2�8�Z66�����;(�P����e��c[v<��7�Γ82��;�ч1zl��K�L� �����BQ	F"�b��������W[�8�a�W��oh
n����Wi�f�l&]35t����DS�e_���tB�cjy�ۯ���z!:��d[d�t]y�%02�e�^Ɣ�<�0e�9v��1�m^#��3ݓ [{��J�tW_s��V6n&#�N�z�Jv����?f�^�^��z���\J|�������U�S�3�!�+}�7I�u�eb��Aف��$�`M9�0k~(��2+��`"�/jv{3�a�$�2���R��A�>N)Y�!�Mx@��JG�$��lH�W�P����k�"%?�[ObCbI:��Yw�L��d�D�کw犁�u2r3ث}������?Jv>�����JuP��Ի%S-of��GiE��|�(�^�_��c���E�>$V�?��V�⥳�_��0��'or�y00ٔ���'?�A���~Di�;��Ϣ�m���3v��v&(�r�@_�:�8k�a��L*qF�`1�`� ��f�P���P	68��i�bF���]�-�}�����mh�".�F�b1����mE&�㘙ӂXϯQ����*	�������<�dn��$�I�'1M�ƉĥQb�����x#��ζ&�ʿ��[#">�xkMx��3/������m�ê��P��B?,PM��uD�g�D̈́��H@�7�T:z+a^$E��{��a����3k�V�QQ�����P����>��4s ���p�3�=�2�|*��CG3h�M�����/t�� ��eQ^�6[:�#�8}�T���QiQR�B%������ܹ��a6V7�ޮ�Y������.݋�,thX����(��
��}�f�J�ǽ��%��q�:nqH�V�(�Hz��-\O���H�M+�0�Oo&;�3�Lj�8�k����G�ƗOf+ N�Ir./�#G�:h�Ym�8OԐ �a�IVOɼFWg���	���+a㢑��ݟ�V\���� �Nh�u���t�ge�VN�Lثk�Ml��B��@�PQaa\� ���IZ쎇���2|3Z'�l�(�w�-&����A�<mL�Kڣ���\�`��y���Sk?Z���v�C�=�Ρ�l7�ٸ	<���p7U# H�C�1�1�/e
��A2�'������[�o�3<����EZ�ǔ�S��]QjK�β�õ�� ��zb��	��4D����/��`�KFу�I:A�
AG��j?f���Q������Ѝ_K���S�SƠ0��>J����y����Q�`t��b5��x�)�BkG!�?k*���p|4�E�K��I:����4w�V\���.���jM�IH!�Ŵ5��KVW%f���)���F}�=[�q�Z2?��7\�����Y�#H�d�5DYRe�6\�{(����7��O>����.2��Q��@W?e�^f�%@�'p0�l���'0ao$�x�5�n��p��:O|�W�p��&��^��@ߟ��=����^�O}�?����t�����Z�a�H9I�1���O58 (��#6AV,���5�*��H'�v� �VI�bf�25]�����0z�V���Rݻ�_�B�ѩN�Nb���>lk�!a�%�:8����`��T��0��2؊�A�6�̣�~����Y��<����v�`ZT���@M��K��5!yʓ*1%��H��a!��=�q�Z����F $��v��?��o�G?�6�Y��c�4q+׭��?�Nk�n�9s�8x�v|�6�N���tP��L�i��Uk�{BoVaW}��^ι�?������{^'����_ �Y���3��3qwW��Ӣš^*P��J�
-�X(���N�@�=�L�ɸ���[��7y9���r{����7t:�9���k�g=k�w��t��40�M�#p��1��[�p-u��ˮ��m�+/�c�w0�9~�h�4���TI	���~W�HMd$,���Tfu]��
V�3 v@�f@Q�{U�TZ�<?A{:g��j��M��O�0���r2&H�����x:��B�i)��ɱ�E� 8��ŗ]H���9��3~5�3�����*�d��\˸�B\\��@�iS��(hn��L��'O�eE4.����L�m8�-t~+�X)$��ei�b`舱��X;��Y6e�і�-��h����s������t�����M$�
�h˫0��T�%�\��.nP�݂*I60fW���P���M�G�?9��IS���7�v���4���]�@�4����	-3�:* ���k���&��e(��1GAiu;�}'�{�	��|"R�f!�t,'��J��N�c%�i��J�c���k��m�O=�l�B���)P�ԚH��#0^��h]�I5�c��S�>rs\h���	,)\������*b"D֒�;������	�f�g�G��A�?��Ö́�$776u�?��+aq=uv��	6ax�k��H~�⣬���('
S��T��x�
vK�8a��N:�J{��D�@IΥ�&�c�=m?����EW�ߟz�Z;�i4Mi��p��!(߆`�������:iC���#6V�ƹa��A��xڙ6�N��[�ڦU+�j��Ҡl��o��־r�5V'm
��s��.L��e��_��ք��j�O���s�0p�7�ZIi�]L.#Z5��U��R��a�E��N�[s+�u�V��:�V�Xc�}��=�	�ۙ�d���*#MZ��n�?�._ҕ��w_s~+j�}���m8�|i,��6����[��N	���	[VɊ+��t{�:������z����5'�э���Z��� �V^Ͽ���[x$���qK^�Ϋ��~�;�h&�`�����ec�H���_��,j�T��x�L�Łbk|�����;$����T����U�ꟽ�`%N��WY4?H�w�}������h��8_��,o�CV��5Q.lE7N	+���x���ђ	b@��q�Y�+��e�kv�ULF):���"�A)F�d��e�Ay���2X�at�N��t�+�t��g�ރf��,��Re.2�(��.�6&�B&�����D�|>���%"552�ws/F������}#�Y��ڰ�Q�t7mb��+#V8�rJ[mѰF	���� ����:�����^%Gr=!��a�Z̠�Ѐy��󺅎�_�v��r�|�[�/�6аg�]���:�����]��+l
 m׎M4�q��s�s�����=��?aA�k���l̸t[���U]j�|��t[c;�b2M��V��yUE���ǳ�Ŏb��a�R���X��X��#&�*�>��'m�f��F�9%��!���″nQ7� �X0����ʦv1�.��4;��	�z�`���9F�����Jpq,���.v>�yb�u&��|F$�W�i�þ�NT�b�3�)�A��Λ�1=b:M-0R�Ϫ4��qJ������]�8�{������"��3��Q�y�����UKd��FY�w7R����|�a.⮑���w����9�x[�f�.���}��J�ih$R�pO՚�c`��4^�$���K��X#i� D���r�i�a�-&*�����P�WF�jj�nPV3��i��SU�2n��e�T�6rU�:!`H�hU��KO�Z	�XVP� ;9�*��CN�`Q������e�N1l4�*Y�.&O�c���\�2��R)�� �6):.����2-�\+�U��hR��\�<����*��bCT$2!i+��zgi4��.����?���A�L��S�"��g=���y��sc*�SSj��<�і�h��������n[+�;��UL]m�RE��~@V�BܑϠw��}�i|+M���Y������S\�x��f�=®���-�Q�ge�� Xz���ѥ�sCf�V}��h��	kV0�W�f�=��:�(+�Y����A�ª�Y+].�,n�f�������[�?�@��=;b���c3��0:��h��d��N�6.�6nj���/]j����G��Q-F�Z|�g���ľv��h�e�<�w4�L j�=��&�~ʠ=��ul�܎)����oTfzڎ+)�M� N݈S����F3�"l7�>|i�8l�h�m�:�>��3l��C�Ǌ��l>C��'��Pz)-+�H7�� V��͝5õ��%�8���4�+������K+W�6���k��d;���y��t'�+%��^�I`� ��L������w���_z��o��B��h�O�u�Jx\ i`�m�yH`B��E�e��HI�����hJq�V�s�CS��s���� R�e������ X���oM��ƶ2IDXz�P8�*�qU�4�Ƣ��Ǐn�Ѿ��s�7"u�n^r*e����#�e�}��3(�O��6�	+���b���WR��{��;P6kd"Q�\�k�K����(�ZB��X!IJ��\��H��j�$�{9�2OjeMާ���mF^�8��U��itZ�7�	�������E�yXPu� �z��	�^���׮��*{���e�횫����z�ig6���3~�H�a�^|�)���}嫟�[֡����;�r��cɱ�\����|>f��I4�6[|������驔�:(��9�9cZ�]~�.LC�x!��._r91=�}�v�����Y �AQB�<�`���Dr�r~��f	IW��\i����SO�k?�=�ċ���d�v[=����`�О�?[��S���)T8�m��2��+�*�_q�͞��~y���hdl�s%���v4Ev���N���Fl]�ZGsU�&�O���K.�d�o���v 8�0v*j�\���Q'�h�<���(��t���^,m>dC�3����H�tL*S(L�Ȕ�`���5�w�P���g��(�z����
�*����md~
��B��4m۱�4)s�G���q�ճ��_|��Z`�<�$̜�&��/,|TZ�NȮ-�����0b(�Z�ǂHװ�%�8h���$��������qg�N��+>	 Y�a2צ*O*�sU��,�ET�i#b�:ky^,ms�L�eGI�X'�U]u �*�k�cy1���c��<V��@x���*s�_��� I�B��"�0T@�)A�����j۹ �锌<� �4�I+Ҁ�/���q��O:m1����i)߸a����;�,n�4c�O���z��m�열Z*%������f�1ɾw�Ya��G�k�t\q�	�cD�i5I�$��r��r�ױ�nA����e�� �4�J�(BZ۸��1^T�Z7�+�*����E�}>�ݖ�{0O}�&�Ӱe@�D�]T|;e��S�Xd;֭�����4v�]~�U6c��ލ7Xف=N���3v-�&��|ֱg���q'���B{�Ϗ���A�&B�W��V&��ؾf�Z�:��'�愂<�`�/1�(�D�	h�4���7��,;Qޙ�J�����fg�{��g����R��▛`��,�������(�fX����z{��5��;�е4�2N:Ύ=�x�����o��� U�[27�D5�K��H�M�
������{o���*3����޿����yd=�R��He�bbq�*�錈銃��%W|i���w�E>��-�O	�;��b).:ɞ��,����m��5�:�t���ˎ�]�؈>	�(�-ی�B���{���������v�����l3ٯ1F��~B���~f�^C҉~�3G[Ѷ�n�S�ZB
f��x��OU�	�S#�X�)҅�!
?�^V�ҟE1!�L3�$��؀���L�0����@�McITD*�����YV�����1$��r�֗ �_m_��7켳N�3p9�|�2&�[o�P�����:�����ڷ��m�2l��r��X�ܜd+ۿ���(�]ƞ-kW�9�,���(����7ݓ؟n�#�r�l:�V��N��|	'X;��y��Gٓ?I�ڙޖ|�>�B�#��|��⹯����L+c��b[Õd�X:�+�Xt�b����Z?��|D�\C��)�k�;��a��X6D��ш)���[Y4�u����tX�SN9��I5א�aX44b	�:e�)���T1��-`.��lO�q�e�f�r�㝿�aCGY>٤9D	m��C;�X6�8�qx!>��s.�W�&�+W+4�v��i% �qS��6XԮn��;I$�Z�x�k���i���c!ݶ��$�pM��ո2���R*)h$~^�vLL�����YtrFs9��Q��0,����R���wґ4�^|�{���w�]{c ���#���p��L5�֩�� DG"�d\G:��$@|�+��.� s}2�M�k�r:$��3d�k]ݚ8�SjFK�9� .���a,�"��(/"Gr@�oB��&�NA������Ϳ���԰p��`?eH���OM��>�|�E)e�NR��#c{�� �}j&`�1� ?�2��
y�e��/a(Z[f��z*F�i���J*�^�}+.+w��e����7��C�<n�8�N<�DVtUВ�.�#�����ղ��I�򲭺��N�|��)D�#�3�7r1�⼬�o��6�t�	�E����k�����@�7 ]��mQ��p�:ȟ%k��93v�4�����_���n��Me�˛n�9S�bUF�/%��]�
K����1:e���{D:(#��(�\�a�v��l�;����8w�V+���{
��w^�_"����c�:�n��OaXM!�d�)��br�ߜv���B&���6J���RL�%M��f��g�m�V��U�Le%����U���B:�N8f�- P|�ttoųz����)=0�Z����O��Vw_��WѴ��|�Du-�~�5��}�L��厬@b�f��������Õ�@�����/m� -}��/�p�a/Գ��n�^�Q
�ċ	����O`��eН<-gq)�,Ę�h`B"L�{���]5N�zQn�t��'O/)3�X-'#�Ϥ�R����ڙ�mk7��_�����aL&L�e���I:߮��5v�-w�y���c/Φ��N
�v#Z�\J��)�,�(�ʏPe���L�Ȥ��L�E RY�bw�\88�D�m��R����MW���� �TLH�`2�z�MJ�y����[=����P<�z�Ȏ8�D�����~�s[�KT#��'�M?��*4�o~y����6a�4�<��w�u���?���<{w�ܳE�	g�:�^x�m�+ �mۍn.�E�P<��L�g����kw���7ʚ��˸�k1$�&����ш�;� {���P-��m���e���K���-����֪��[:�S�D���aB�3bqjQ�04%Pˋ��DG= �O��	;�B�ڗ?�X8��r5 ~��=�����m(����5!�N�|*3�¢�0�u�p�L[0g������#���ׄ�(�%Ax���a�#YR���dۅ�=�N?�LJ�C��_d�����|���]r��r4�{);�`��z��h|7o��<�dܭR: ��!��=�vn$���v܈1V�=�(*N��!��NTԴ�!x1]�T����.IqR��2`U�հ�5 @��B$���/�\���K.���`����F����ٳk;��\�(b�6�K������ս�T�>ޣ�kSu��;9Gm\��n���Q<X,�M��+m`��1���΢&E	d����K�欦��� �T�F�@�n�<v�r%R�UW�R/Tzw�H�fQ#�Dg���ꘟ�N����`SK{$���9�&9Z�1��C�$ ��1��V��{�p�l2�/1�0�X: �x�A\�h�����H�VU�x�����iN$�������N�rV�}����M����??H"Ox�LZ���Ow������Өa�T������.�E4�!�z�kY���*�
�&1p"7þ�+�4,}��{�7�����)S'�r�:�p" _��6ir�]t�o�6�7�q�t���JƥX�Zr���=y��W@�F��E��h�������f
+�f�V��H̴�q��YX�X���}���Oa%Zb���W7���\V\�ͬ��Y��K8�،E+�2ࢬ"�Bf�rd�*.0����r�ȷ��)��F x��K�"�C��
�!1=\8�r"l��>�`U:ijІ͙?�a,�w5N�m��5���-���f���� m�t�SܸbH���l�3ֿ��5�b������gj�� �e��������V�.��Q���q�I��Ctbd�[:�>�z�(���,��+-�fK���"4z:>}��(H눛���q��|%�!���d�j[6��}8���X�;c�fJ0�D��ϵ�;wؗ��<)v�ݷ�q�m���hOU���9
#��)V�}�qL�j6P�HR�4Ib��6�"%h�9�F�yY7��2u�X�"?�Oa��!�&�OXv�ԓ��"��٩臒lf�˗}`���4lV.{��_v�]y͗��N���DǓn�>�89���K_�Ʈ���l������� �Û��������W}��8���~{56O2V%ڹܫ�3�6n>����0F��׿�`��s)2�wV���bb�pD߳��Yg�=��3�'Xku��&>��cVTD04r�������@�o$��2U&�>=[+�q�
��$V���p�I�I=�^Y���duɕ��/���8�/dN�NN�.��~z��z��M6����Mw���J�@ KC%�G�*/�n�`vV�t,�$����,��Ek�)*˝^�X�>4������Z`�����ݸ�*K]c��=Uj�S�	��DA�iQ��e�H}�s��~�6�Q��=CY9������<�	ˆe��q�m���f]?bZ�����չY-&U-��t�]�b��'���ͮ�	*�c]V���ȟ����;;����Cخq^Mp�.���
��Ts��Ù�e�/�(�7j~�.� [�Sx�:\�i���8�m`�+��u�
4�=���s��I�[]�;]���~4}�8keq��i�i2X�����
R2�a:D�*O���Ӕ�&�W$$��9-���SS2GV�i�D��1�����@WR�ڟ�sOA�BM��MM�h�BGUXTl��P��j̜��LS&�y�N��3��=�$J���jγ-F�Z~ԓ���+�ӥ��Ao7j�C��Ȝ���K���p�8a(;�5�ݔ?T��)�⣎�s0MZ������i�4MM��Y�qh��!�v�j�y��N�s�bK�����d+����̂n��E{KKq3QB�0ʚ�E�K��V��q��I��}��*�"Յ3��L��A"z��"qA�b3��'��U8�BVY����
m�X��BW�3����t�M���.��x�� ��B��(V=�m+�X���Up;��V�Xʰ
���i,R%lET;��s���Ī�@�bGu��{�1V�c7+���0n��yЎ;j�=��k�P��Lfql���#Y�%21ESVp�����w���G|���'1a����l��k�4pk�u�jʑ��×���w?q+�q���T�#�h�`�Tb�Pvj$���&m����o�;�f��`�̓{9e���:��uh�Q	+̗���ݸ��6��I�"漖	a4���Ӿ���L޳�+/ò��LD�Z)x<�ݰ�2`5jY�h���&�1J�!�
�=�<�j@=m�Hc�R�D�)I�{�@Q��rX)B2I��N(C9߳h�>��2��T�-XZ(��ŧZ1]ݫ>Zng�~�]x�y����{o�r��m��f���
���/O=�(�\�=��3����j�I��|J�����ŝq����fϛE��>{���05����V���·4d�y�[m��H�Y��捳�n��6o�C�P>��/�gλc�I�	�v̱K�Om�?��n���HC����پ��Wv\�a#��~���/�+;�nP�5PiP�; ��If�����t�3�0�U����B�ba���WIwl��M��#�(��@t�Ӓ&q���&�zc}�d�O�Ɋù>�>�ۋB5`�,Q�l���7�<�.���ztI	 �[G�4�rZю��c�n¡�����px/A+G)���%X�CחGV��D�_0b�����2���E?7��9� M�ٔ�Z�K�Ё���Ƴ[~��-���1��v�3��}�D���1��< &ГH)�+_����,�+�o{ ;��k��o�:?�.�b�<�L�����)�kjƬ�5����f*�?U	Ђ��R��Rf�9@ۢ�I�U;Zb��I&�Rr$�6tt�G�,�V)��6���ʈ��8 �8� W,Z~:�SѥX(��ڳ�2T��z��ٔ�#�w����r�9�s�PV	_l��T��'2�/3#�>�����_��q�\�H���	5C�0�9��0T'n"@��$�p�H����Ys .���@U�\�B� �:n������b�\z7o�]s��8)O��.<�&���p�e�ܨ�&]`{�gS���<u��jL�g@�O�O��NV,�N�C�p����.�� L[9ځ�Hn���lth��[D$�v.���$KɉwNک��y%�x5tه��`v<��G�N�c)��U��z|cCk?��ˎ�q>ZA��6� �c	ƪ�5��0;`q ��J̾���#�h8s��F�5Ʋ�[YmP��V%M�&��(V:���b�eD�X��;F�+��q�h��2F��zn�&��fD���IX�K</�f���i"X�V�JѿQ����������]d�u�(I����o� �I9w��2��o~�e���0��qݫ�#��J`U�qG��]������OڍOb�����=C�0�V�y�0T��D0�z@�C>׆+O��0�Be�C�]�A�b;��9�ȝ�Z٪����TL�b1�M��\sG��-|��rWW܆Vq/�B��;'����;��ϵ�ϣi�R��oH��9k��6�����^y�w�-�ӯ����s�t��.O̷!�v�v��������$�U�ڤ�
�[��?� �pd
�4%4���C�Wm9�5��W\z�=��C�k���ׯ�k����a������i��~�����`��J�]�=�|�~���2�,�H1��j�{{7���,���\m�9N�xr�M �U��o�Q9a���Xhi�m~�}�B��ԍ��q�X�,sv }mN��cN`��T��ڃ�@[uV��r�q��s�0&)E�*��st\��3П��^%dOdZ��^q����;n�ܻ���~���pxF�f�7�U����\�x`���7�Ɗ��r{���0���w`�p/N���|�M"�F�1��O:�]�����r�T�˖� caB�]�!��Ә���i�hCK�f%{v�����q�4@T���O��(QL�d�^Et��X>e�Qh	��o �w�uc6��z�*$4#T��F��h���<�3l��X*,�:L�7�V�9��<�Y?RN���"T���Ȧ4�X/��Y����y�ɽ�j;�62<����,x�Y�
��0���Ju�N�0���rn����K�"�n]%�(fL��X
�𸍅���h�f]ۚ+��k�*C_�DL�,����(������K&�p�ufr��PV��d�'c�8��>CY�.։:1֙��ґ*�/k���l����)ˎDț!���<(�,'�w�k��15=��1t`��L ٤a��TU�<���Q�} C�����x�5�{:����gK$iT�T�D�s�FO����o���(�q)���"G7�ǝ��q��2'�R��K���]�;.���� L����&E&D���� ӂ�wkuP�G���ڦ�fŔ]�����.�Qc�0`'[��T�xbYQ��1
��1��"P�"��a�5v�K`T��7L�K�p1�_:�$[�j �'w��ŔЈi�}Id5\� ���.���}�nYQd��$�3��"�������4[��}��<�հ�=��Y�|���,Z�wl]K��ط��ޭj���s3��p��q6�Db�r-���g`���m%��ӵ�֠�N��ۋ���x7A#��ЉBK��9�z�E*=���Λ+P)�e'���'��pMJ�JE0j��8���s�����_i���q��c,��B���ȺE��z�*ꨒșNX����C�3­&k�vt&��De(���>o���))>`|�	��}=�)'"ҟ�9-f��I���i��=a}0`���j�C����zɹs��f%s��-��^�<K]�b����]���]�w?�n������ �қ��Ŋ���kL}ٴ���;JqC���K����,��Ƶ���f(2*Ӷ�*�7�o�ϝr&"o�?ݽ��i�H¿��>��T�i�o׫��{0f>��7�(��o��k��^yӟ���������_���n$�b(F�5��w=�UH<�N�N�r�9F������އ�&�g�l<�m2zS'���{�u�ɐ�`�>ƑhEz�L%��x��a��(�E���$`=$#�L{�÷�¢��牀�h�7}�v�9縼�x&�ND睰�G/���g ��8"��*+~�nl8e�{���h�&���o�i!ٮ�i��Kγ�n���e�����u;���U,���3�Me]�N���[��;p���ΰ�_sڲ��+)iuGۃ?���~|O�c��ޞz�Y���I�V���^�ϸ%�y�e8 ���̟��K�g��N'�n:55�u�@�l�G�x�D�!������o���t�'`�6���&�j�$�T46e0�H��f�+k��M@�Y��kF���ߙ��~1����1�����Zi# ��w�]x��'��r�[�㋐�$R6C�e߹�z� �@�j��.�����Tb2 
~���pP	��O�_=� ��U$���Xz��w�U�g�������7����k�b��������ӗ$��E6h�/sZW�g�!k����'��f�%��+*1��1U3�ZtĂ���4�(��w<���<�Z��خnۥy8��r+��vr�9Q_��$�ok�%�E����fq��9F�.jhQ^l �`�)�#v���F�'�2���}#�`����MZ3��%$�h�u	�U�Խ���OYW'����!C��kjh����rd;:�j�Ń������G�vl���k�G�[DU&7]\�E���� �"���g��. ���.�M�� .x11}ا0Aь��Y�А���P�d"�X�p�B��q|���ڑ��V*�lli�#TÂ�� _��)6���'*=*�?VY�T"��ȷVB-��ܽÎ��f�7�)cDp���;v����kP�Y�s�"X5�ٵ��͞�s���껶�-�\�s��;v��X2@�_�*��TZ�	��,Pˠ���\,�P ���� ��9 ���$kB̟-#n��à�s�t�s�6֗Xod/ba܈9�#ȻJb�P�."���p��z`��Y)eБ�
�Q�s7y">Di���m+��p�h7Z��V0P�����p��^h?��:{��-v��g9S�֞[�r��C|�w~�W{��U.�XV����5\�j���nI������;os�p&�륋Ւ�!�0V)Da��F�E������p��RU
�f��˙[r#�8�������J3�I{2G�v��?����S����=�;J�m�o�����϶̄.��0�����=��{3ha�(\���u|)%%"鄸B�_�����ۏ��NѲE��Y��d���` �_a�>�9�����OP�p���Jǥ�u�ʾn{��S�����P`]׎>C�B����a_9�����PV��Z�`�N���F�Xu��tGF�s��/��[:3��]�"U��E /����, d�f��	Be�L<�f}�m!�篏a�B�iWT����׊�h���� _B5�TQ6ه�|\��툴��L�W��>X-&�h�ZC��"�DǖJ�ᘒΞ9�n��{�{���逋���_`#�؝w>���(���y��ƅmo�N�/)�5LV�Ĝ���Um?��Om<�j,�^h`i����?1�6`�<Ѿ��/��100�5T�0^��lE�pO�^������"��o��0���V,�5�1/��>`��Mqa��=팳��E���?�ݮ��v����]w>́6Ke!s�$
Ȩz�u�&�ʳ ژ�@r��&۹q+`�2غ�lʬ����CL~�]J�*�&bG1�f��L�b��+Z02`L�`%mtǋ1����ekW��M�R���Ob�F��vԒ��n���^ʡ��̬�;�[|��>����ACs��(��s$�p���_�}6��Io�vĢ���yͱv꠷�ԩc�ǫ쓾  �Hc��*�(C�ƃ_��,H֨4 )���@y2 � ��l�����su[2:pr0c�^�-w�KO���A�������L��()��U�S�.����+]��� m������z\��_��!��#�>iH뵰l�3Wu�#��8Ъ
�@����s�q�JNJW{�q��X,�'�)���g1H/YxlbdWgg8��TN�����.2���Ҭ
��Y_CFF�'� �H�f~wԕ��"x]8R�?�G�QJ�nko��������М������OLU,eֈT0�SS"�S� ��b���r�jİ6�\V]W�.Y��mE 4�����S�0:[D��7�7F&ЁȘ�@#o�(2A��1�G�[���w�M�=}G���W�J}���%�W��:WjL=���x�I����R�+p����n�h���ߵH�$�T�E�L�771:���6����Km�c=��Ī��
��j8]@��@����E�o\q;�	��������h[�AhU�E�_+�NL�r�F� ������� �%Z~^�eª����w�I�K뭄2iyC9�}�=�saN���>��o٫O�hw?�������:�h_���0��Ȑ6���h_�S��6~�X4.�6����x���XMk���i�	��Q�I<�T��f���3&Oum�Ut��SQ�]	z�/ԣ�)�Cs��ǣ�A[�V'���浛��� �s�Me9��ٮL#=�駜L�ĩ��a��*����y��A�fc1������-t�IkǷ2C���}�8b�k������;8�Fwû%����.����4@듎�'�wG\�h�~ת���u��\��>������H�ue�.��8�� ����f7,l$!��4�4��B�N�=Za+n�㋖���B&��rᯫuF˓�Xe勿Q���g��Gީ��}�����a�ԩ�C����P�DR�ˈU�W2���3U�a �=)��ީT�/e
0*��x��F�FhN�8�xX�{�g�b��h��Z�C�8�rlM�^̍�6 �E����3�ui�y��G�a��ԙOG���ß��� �z����v҈t�]w�<���?�1��xJ�]�:i��<�!�ʻGX���2e�x؛:����Ǟ{ڎ;�T�.`U(�-<r��"{�mӈ�H���3 ��b�����w��n������?�m��Q�䲳�7>py��&��=���׮�::�f��t��dC�x:W}�<��fۢ9����>yǽ�O�3Tkbܡ�{���h�M�8���~4�_��[���]0}��ҙ*�"4?�0U�0�q�U���Y3'w�a+��i��XXb-R��{��$�֌�S�dݢ.R�n�p�"wΡG���ł~[�[ �A�=@��r#׶�9�`p�"M����G190���u�L�փ��h�R7c���[ 9\�l�6A�@�b�N�1��9z~�wM��
�v��?�H��s�%)v ����Cq�2C���U�ա�+�E�QeV�Ee]�2���|������}hu�?k;����O�
�ʓ.-c Ø�1������<���pʑ��p�U>�23�;$p�	���.�}�6)iԌe�)���0�1�1�O������ t�u�� � ����$����������H�-FT��toz���d��h��2|ر4�P���8t�y�P2�� ,�A())��.��xVi2�+��=fe+B�F�2�^O��l1�&��)g����:�/	�g�J(��%��b�D�F%Q=r^�L=~Ū� �|��O
���^	�7�;����0LC���	�Du�U���� xf�1�v�Y)���1\���Hʓ�G F�R��a��+��ʹ쪃+� J^N�-\,�IЀ�a�A>��tX9�n��JX񎷜I�(3���k('� ��D��LdX3l���˯�9ZLY��aV��\(�5ke�������͟�^.�\��t�d�_B�����+	�V��p�s�p���iD(��Zl_�+�Wzb�[��n�(ʥ	�ОXZ��)������$�G�Lc-��S0IL����,�Cm.�:���q�������G;��9�ؓO.>I��]�L�T5������^56��� Dli�q����$��/ׂ��}$��Z!��$T��y��D��M�qǝnr8�]X��iT�t;g}��ݳ)����l���_]��r,VFlR �Xu��S��dbܳ{,Bx��}�0�\+���\�=c�.��[Vn��/�a[��c��٢�\�YE��ˤK�^���Iz ��&/�U$_�~i���rh��h��r����_�u�_K�[$�\W�*�X�ˎc@�1Ls>�f�Xl��±=�ȊR;�. o�
V����윳/�����6|�p[�|�}��?��{;����=��R(e��-Ӣn7��"g�~���7l�}��v����XhV���ȌD�/�myC,��怵�>&Ҍ�*MY��&�e|���f8�0k*���ڍ?�����2g�i�����b[�+��G�#�i?��w-�h����&�nG�U�	P�k����6}�ilk�
��U��E��fQ7c�lΰ�,��^B���kV��O�e7r,���Y$R��#Vi�TК��/$�`VK�Ņ��Y�s ��㜓�xk�"��N'F5�DK$��	_ K��� XAl���B��>Qf�A �F� ��tCi��:����_T�1�!�.� �
����.+Y:xc�b:��}y�gB�>ķ��nv��捵�r\�F;̗����|_o�)b9#[�]�D}�쐔e���0���~��,F]�+eF���à�_��{T��>===��b�o1~RJ	�Ն�x{�ٺ���ͷ���� ��7ޱt	~�}Ţ)Rсimc�F	�3�i;��T����m�7F֑h�Ұ�Ħ�/+3g��r �ڒU,��קa� �����c�j��(�|��Huꗟ}�Z b907�h���EO+�'1�Pn�JwI�:�#�|�٧^N������6r�����{V��,;�H<���nD��X���Ѫ�s�с"}
��� &QJ��Dq50g#������v%Af9.��,��铀�����U���+�>�R� >H��08	��!ٻ��ba�)��âu���K=:�}��H��Km����ܘ��t.E�X����z91�V��B�E�DL�� `�* W�٬�G��T�~$�6�v�9]01���Q&���CB�J3�7j��!�ĀD���<&3���T`��5x�'M�`���J7L�_��̎?n�-9�H{�ɧ�]�$Ͼ�
k;m��D���{�t��_��.>�ȬxUlW�m��G�@���c��r7�[�I?�V|Z�qC�u;80v4������9l� ��`E��-�_��t�h����La4�:��w�B��	���;��!C���𳥁R��� �,zd���=ݍM�D��@L�츔2|m�~4����qDw�-$�tTeq�㺎�AtV;cM]Uq0^�
xf��` �b�p���}�sTvQ�����xSل����q��x��]s��o&��w���¤y�ģ��+aBT���8Z�u�8|�[�%� ���8���S�$"�������>�θ�[t$it�i�:���1t�Ȋ������\��yo�������;����&�]d�E�MXt���{��6g�箿z�f�﯏�����{X��ٝ�����/��IS)��]C�0u�|J����{���Ү�Ʒ�3{�r`�~r���)�)>gq��o_���v�u_�[n���/����/E��d�1,�Slgy��-��p���k�*��g���YlB�����r����w���H`s��/H��=��}����
ۏV��c\�'Y#���K�R�)i&��y�G�3�������tmzl�+�sm���@���������&��p ̛\���~��`G,�&~�)�9�o=�1=�d���z�i t�Vy��1[n]�0@Y�u�V����`�T����}@����[`u����*����	�D�YA@汌*�c[��2���f9��"�Tbt�h�Q4�XKo�57{9��[6B~}��Y�=���yyy�O���c�J�n���Gj���z���ށc+�A篋�w ��U�������Z�T�{}y�.�y���d�#C��=#�`H>�o����?����Jy��@�� <����J�!`kdAƝ��4��G@ ���g�_]O����9  @'���l��{�a���Ķ�؃��L�v&B��8H���H�j��Q&�]j�CK�jH����H7���T@�����`l��30O*������J 3�ۄ8��M/"�(��-̻]���s���j����*��I�k�Y�vB7�U�XE�g+������������葔�j(ä���a��Y�����.Nu�l۶�!���U�F\�w:�d��D!W�Ň��+���UF.��dʚB��j"��^�LK� �*4!�fN����y��U��x�q�K�Yw7�. ۏV~dϿ���xU���X���ܼf:�DC�+��k�پJ�դ<9�bb�I�k��KX�F��OpAup`�� ��W(�M+�ï�=����	��ܑ�NLp��
1`�J�=F���̹V��z�-n��� �JF�
�`!	cQ6{��@�\�x�z�c�c��" 
]O?sS_=�N7lG��6�ί�t֣s��5)ֹ���,��l�;=������@{�s�^�q��K��I@_�l�V���9j�ׄ�F�X�L�O�M�"��o%����1t1H[�p"�N8�z��)M�� ��}W�Hڀ�9��Xl��'�8$��Y����.`�r�%�!~�����P���V3F��9k�k�׿��uԑ����g�����#�llc՟@7�^���{):��^@`�+�F�#���6בʱ��4��a�Y���'w��y{����(��a�=p�{U��pS�K.��Y=�V��w��};�����k��?�vʹ�Hgr����(� �0~�o�Nd�Dʱ�`4S�e�� ����2pc}�W_z0w=�w���V���n����6y�͜2�NZ0��9���(�~����mȂ��W �.ݷ����e�nSi�QW���q�W�K�O��M����>0)��7�2�i=���N���볼{�c_<���u�����X���--�v� ��y�������(M�:����ˏ����m���o�Ǽ�Qn;���у�.X�죘9l\``r� ���"=@����{���I�:���y��X?C�c�m[�q�c�P��	aA�R@�{/�\i;�|��(0��k�1��]G�CS�]Kj�P����pk;�'_�N!1}����G���nc�5��%�>5�������p�p��괋����ɦ;'	Z��'Қ�a\��2nLV� �J���CQ��J8>_������ܵR�c#�,Pt�uW�ф�Q8�w��ŊH��t��b�sr8]�a����ˠM��/��� �e���B�Q���Ǆ1���X�-�|�2]C2]0b5�h���4�����FeXl�6��zڹS{i�d��#�>�	)�r_:���|��;�`��������ih�*��t�`J�J8N��nh��3��Vck���t����`��Uy뵗m��M������
P7�X�IǱ������B�[�:�"�LKm%S�j9?Y
F�ʅ��E�p���s>���v����Eǟ��kc�L��i%�aʘA�B�l���Z��}��٢#��|%2H��M���	����ɔj�'}�Y�`";�~�'���#Ю5J��*G��`�`F,�B����bG��������SL�7��A��ba���wq��: �X��sJ�q��^�k"�#hea��h��ع��GC�e��m'7�EQ���#=Hx?"�����_!ɧϣ���+���&���Xu��r�y�8�﨑iܿtWQ��hU::��#�wWf��R��Q�a��w�� r�f��J���~��O�l�����'
؉,hn���05EhBGۨ�6y�" ����:7f�}�S1f}��Ka R(��w�3fγ;��R�zđ������w�#��Q<�ƣ����GjADЎZ�]AI
M�`|Ȁ쏷�~t���d�F��%���,���b���N���jW��5���`r:�:����� W���}���§�������΂��fM�����u����u��U$�Y��'o�6�%���	�Ƭ5��wW�mo,{	+��ujfq�@��Ƶ� �;�l(V=�&Z�l<QL}�9E����Y-�W�6�R'�f��&�:��T)Rh�J�LFN�D�_��a-=�&E�����G����
h�1DH�8�A��p�����(���H���1�^�NO���ʚ�����C�x A�]��?d݂���h���	 �o���n6�66����"X0��Ҹ ����ޫ1W D���:7P�u������z��mPǰ�	M0�����i�P���)��b=�m��{���k
4
љ��/P�c�A�Q��3o�n՝��r���A�x�dC���՝��z�tɵ'p���>x`Q�� ?5����`����F��G^��� �1�?*t>Ч�l	����@�N��El���2��.h�4��0�b
���%/.-ױ3�6�(��R��sqc䑿�����l���P��B9�c��Ϝn]L�1�-�����| �nt7x�e���RcydQ��r��p�ެ�� c� 44"��0����qI��8t*ˢoJ�#���>�D�)�[�)w�&�n�m����M�a3����F��š�h��=�7�mg�#���.G��a����������|.������`�LN馓���Qc`��C{��d�g��Exu؆��--��R2�he��ŧ��Ym�b��؞D�:�|���r��f�ǉ���9��n�;���cN;���co��lQ� �|�S�;KmĘ�hlle�#�>֎�1{��W��w߳�����O~h?��A,6�r����D�$�@)��M-�Z��:��,�E,	�i �`� tJH"5���Î��O�T����I"��<�ݯ��vV0Ͽ�.�[��aKU�매����y$��d&�N��Z:[��72ߎ\0�vm�;�'B3��.+���Y B�L�F�S��(�u�|!�bRl"��y<ZZ���
�Ӡ��G�ƢD5к2��G�)i=u��t�Bb���]WL⚑
膾�sg��z��}ϟi."�z�B��������H#��?wy�sl��24Y��=g�ڑv�=�GX� ����I���U��̳ϵ����؏���o�������v�%W��ž}�������1�Pl�S���*��V]�����%�RQ@��q�`,l#��
��a';��v�p)>������Fdo��e�t�����y����³�VÃF���ѳf��EX����'ڃ�h|�/�i���N۸��� �LjR�L�8#=ߢ�GP�u�n(�]Gg�۴�Բۓm�K9)�,ΐQ���q�z)Ŏ�73��ls�͚5�r��݁��n�Z���X��Ag7&��Ĭ�0Tc�o���[&�k?Ȋ9�աo���˛������9ː:�A����6n,��Y����u�����;�k����� ��� ��
�O�C��<?�y�"�+ ���i����y�<��;Q<#1?�
]�y���{ [�V��{o.�@���Sگ`��;��}�.	��\{��WI[�f�]?h���ب�h�a�£�cU&T'��s��S�0\ZZ"j���`���(��RYTI� 	��"0U<�<fA�}�z���V����<Q,%�5�V�b��_���˚�I%���#Po�e�5s��7_+���{a��C9��V����5��xA��I�k 2�W�5���x!��[��q�O��zj�"����7m^cy��j|b�=��K�sG�c]D�щ�J�T�|���̡�32��lk'�ך �<:0w�CS"��D�q�:�1:<n�����j�3l��m[i)aW�(�4�� �et2�������z���b��5�4{�=��*�+�N]�u����F.�:�TW�j����2B�u5s���_G�DƍD=�-���tط\4rU�r��c+�_�'�e_8�Uk#���l����Ȓ%'u�?��[�րO[z~��T�I#]g��}���G̓�w�mC}��U�|����t��v��>S���{���o0a�J.8���~x+��y��`o:��>��50w�}�v{�~���7/���9	V�Y��`���Ю�1TE@�i,�$p���M|�glٳ�ۢisl:��)'K��W:�6h5p��Xϵ�@x�3��m��ve�]�A����bt��3�d̘� J H�Y�d�N+ZF�Q��1����C4\��^(,�c����c%��}�uv�UW�Iu�����,,��1k��K�h,�����:��}:��锸^X�mߵ���̜5ӾI�نu[�o�ne��P��͔ 3 m��������κ�>V�4٨����M'%��gV˂R��ɱ���I���\�7ű�s\:����'i1�Nnf�yN�G�!�x"f1QD��kal+� ������@v ���oA^�<dƨ�`û�f&��괧	��Tf��f<전؄V.��@���u۴n�	XF�W
��bL泦͙����^x���(�u4��$������)�X�gϚŘKg��0t�ɃJ���E�X�	Ӹ�}�I�������:���Ϟ9z%OO��:�n�PH������~�Q����v^0���]�x
�<&�����\��_��� e�a������{}�?�
lJ��֗��
tn��
����&o<�^�3�T��?=�L���]�T�{��p�~��7x�x�������y���<
�y��Dm�^�ڃ��ߤ:��9����A�v� Ku+�#|U��n�nL5��C��� ��NVs��3 b�o�d�5�-�{�s�ʭ��M�ۚ<C�,M�6ծ���Z��Y3�W_�]��h%��@�A����08x��h�AwR-����]���D�E�s���_��A4��?��j���F�^;Ds��I9�l)m���ǁx�d�ӯ�黸(��i �t��aDjd9� �A�i9V�'m�#��a"`u�L�J���6i���؂)�D�G)s-�m�A��a��G1㢣;{���6�Uc�N2�(�V2�_=
?������o����� @�Q���FAi+O89�`�O�,�sbЋ0h7��DA�~�����~r���Ä2�r�X|������FsL1�D�SqĜ�����N$��t1ťXڮ�d,cW'�-��v�5}��ݸ�V/_X��+eh��έ�h��09���%G��I���u�l:=_���p����e����$�����������_t��t�'�(�`�C�{z��^�!��K.E��lU!� �-�M��ۘ �Q�	�q��[�Jt�є&m#ˈ�g5� �B�-��Ȥ�&����Le4�C]���.@|.����
{���l5���
lZ�q}�9}�~� �x�	���c/.��\�u�(lٸ�u�����o�<�]�9v��K7q-&����0�~x�m��u���u�SO����~�E��ysm+v/5,2��ޑq��'/�ـ��e+�EG��Ǣ��`f�Ak�x�q0z��T���f��ي�[QI�2�H��|VWW8Q?È��zM����^���SMEB�ьIS��jRT��������M��XGÎI����|�G�`ţ�������}-`=b8�C:���m����ԓ�"���S�B��ΙC�&��}k��`����#c�8��]w۸Lp�����c��U�^.���.�Ă���I��ca�%iw����:�t>���!敦�I�#$�Á�>��( W�
��P�Jsݖb��v`DBo��yL�,]4~�@�'^L�?��V �|L����mu&����<������S��Ib�1g�<���7����}f`<2��O�g Hz\㵎�zY��nP=?B��:����=P����=o�?h��γ6?�W�-	2�_��Q��������^�${ׂ;��y���8V �m��Y����8p�S�A��Js�a8�!�dGu�����嗮�:��a��pnD87t`�%� B��ĕ�c��wC���P�Ç���v�������֭P�|v+Z�(��v�ǽ�!����=
c�o�	�M"BG��>�'�ZXL�5�P��V-"Vo�JZ#mǪ]���=0fU�hc0�꫌xi$��#+/���ܬat��Y��!t�kB#�Π�́����O��M�D��tm��0z;i�G�.�3������++,a<���9tlʛ���?��X"�\�r���֤�ɰ�%o�^��� �"�F��^.����A���V.��D�W:�ZZ�1R�h>3�|u�p��"TQ2��m��ιY,� ӊ+�hZig�Q�u�[�mweS�L�|��#J,$�+4C ̆�����%�b�6<�v��ɠd�d��Y.��9���X�ܖ,^
HK�S����$��PG�����Ob�����;��gL�?���=��l˿�Yz�W����[���0b�±^�ar�4^�Z�Va����3A��&�9l��	�BX��狰�h�񝫬F��
Jve�v���(Z%M�6m�9e��X�(�j>�+}x����b��\�V@���J>�SV2�r�6�+�iӦ0��X���#RƝ��P,"4;�y�%r�*��{߹�N:�ƚm.��SO�7�Yi+W���XU�w����?�.9�f��}�6{��w���Yt��~��r�D'�qe�����E�;-/k��~�bJ���{�w�aLl��  ��2WY8
#��x$�J���
��#��neLE�
@9��n�%WSC!`TM�-��4��ݔ���k`��	K�謩n`���eD&I5��@5���Z�3#ȀM�C��}m6f Q�ʜ��/�� ��+ِ\�w��B:KG�22�����6�܄y�(�P�1����
��UF/&�r�.l��bl!c��m��k�J�í �ls��a�LD LpD���CwA�����`��i�4",��H��w������H��a$�8 �?ԥ�@��+}s�c�䰍3����6)9���:4�j`r[荑������~`�= v�����\�X��\����$𖾟.��`CU�?X�|��
l|`�=dA��S�}�3��r�_��Lt �m�O{��Ι�@�� j��b���{y��;��QH����(�q�3���|�k��o���s�̀�^�@M�n��BWI,,���\e��(�[9��(J���0b�Q���  �3KyTI��;:2�+�{���_�4D�uեx{��t���Hd�2C;f$B�z��� *tQ8c�04S��{nl.����whmW;@P2�L�Q}k��ڴ�':0:�"&�Xy�W��W� �e��������A�+N���O[�����<E�X�MKy��%U�>���U���K[;�=G⳵rY�e1�a� u0e%8F��]���e�:Pd�QV�XM��|�6���� ܩRCA�.�:J"]�"ɓ%Va�JZ]��Xѥ�wR��k%*��~   IDATv�V�<?	�P�nV�1�9�[&g{��'D.�n#��6���ߍo%�*;PRA���+y_d�5�����OY�c ��4�CU0"φ̞΄>�
Ї��x�Ύ�g��v�i[m<����a�b8V�W��VQ���t�����خ��:�>x7�'=����7ze�5C��$V Ӥ!5A'�t���ZD�Y��l�'M��K�����%"���`�����rԸ\&�&۱�5�0�6gy��-�������tR҄��S܆�p�}����;�"SV�h_v�P&6O� H�߰��P�}|(q@���h��B����W~��c�N?�$��R������/����� ���V @���;���,J�/��=��$e������t+)�DS� z�6;���m;:&���Ib?v��ηaxJ�h�>���wٍ?���~�zd0u}�>�%�t�7���=I�����o��q�=�B�=:��~��M��h��/^�m����9��a��6c�Zo�Աx,�9@ݡ�}�:S�׮u!�7��Vb+�Zd���o}&<�֮�n���n�+¾D�������3Ҏ[���`���C�oƬ�����,2zz�#Y�؅������[ɀ+F�O������/�Ϟ6�D�A K1�
��Ẉ$�}��cYPf���*ư�q��D���	A��a�'a�1Pw�@�0�8�ۼ�	�	���,�cR|7������t�yα�/Ǧ0��+s�/�(���0��X����恃?�!b޼}������3�3�\��<vȉ��:X������������D�m�O�/��r����I���������;��U=��!P�l�=�4�y~���=���m�u��� ~9����v�[Q1�����0YFKB���OZE7� �jzk)U%���hA�h����J���	x �q���.q�A*-� �UO"�`��]��[os%�`L�5�`lH[4*��k���C��߁#wB`��@��	��`F�jh�ޱ��ߵD�^aD'u >��gG��OV�p�rL�g$ʇj���#��&b;�ɗ�p����*�����UƉ�C�2������vCeoɶB-��FKK�����8?o�||��ʯI�0ζ4�GX]/�4�;��S�fY&�=<?˾t�g9F�l]���}]]}��)����gŸk'���sB��Y�F�ҫ�W���1��)�-9�H�h pH
���F;����D#�I�C�sN�r���l��qCn�]{�	oΠ��=,��M��{0d���E����rw���yLjQ�b���##p�Yg� 0����N;Y	������7���
��O�b�Y��(z�4W����J&N%�[8`(b ��k'�S�1*e�Ya����Ri&�ໂ�h<�'��8Q�>����3g`��I���l^�6�nj| 5�3A��w�U\g*Iƪ�Y�9���z��Q��$dN�ѤNJ�0E�М�au���f�{�˚URG/�z�rXP]p�ٔ�Vٶ3�9��m���V$cB:�N<�B[r�4���>��d3���RB��p��ee��e�^���?G#��{|��&�0�.����g{�������K���^t�O��p�0��3NV��ڸ���aѱ��b�@����3 �\~u�kf����bѐ�1�bL ��7�F3S����{\6�w������_�ܳ.�o�[6�ݼf]�m��e����a!�c/���늖VU���X�R������٘��bŊu�曻l��	���p�'�񲁮�ᣇ�P��x���yJ�8K"I����&��b#F���~p�A-�E� �>+�2'�^2G�`�z�d�ҩ����y��(yI��`�>'P�$��N�U��8���W�<x��f zyB���9�{]r���{�\��=܈彧cZ���+�y�)||)���C��~��>i��E��y�tL�SY~l{��~���7�(� ��X'�!�߃ , �d3���1�=���}</�V%`ǯ��`��?�wh���:TRU>0�k�����������)�x3Gp�6�[L���D��ڹ����.&�u�:�ղ:�����2Xw�����y�Ť��$��ɊA��$�;�fb,���-\#�Y��<�-{$Pe2�9�r��Xi�@�k�F�V/�D��UԄ�;v|��5o�e�:���	+'�Jvm�hF�Л�bz��HJ���l2z�j�pw�B4i#
h��r����c��l�� ��n�t�Uv&F�]��*+X&G�RW]�r�t��8�ƒP'����q�����ڎ?g�}�ګ�݆��p[�C
�^ʏ\4� ��*ϛ(.�N��0W��o�7�xӅkK�! ����`-t�ESQ�.%eպ�=�b�x*���s�u��@o���(4��/R���gO�`s)_F0�*;�����8�q.���e�UFDu�n�X|��2�<�*����MGl����5I�[X��7����&#O5#��:G�l=�����	��O�O��?ۣO���@��k��2Ol"d���E�p���Nr�- ���<�$W_���a4�R l�*�g`��eW��By1ۗ�����#B���<`C�qIO���V�k?����i�$'���U�p���\]zl�&�:� Y������&uW`�i�z;�����q�d:M�6m$�k7�����,�t4f1h�r�s w0�</�4�1Ó�a#�b����h�x<��H+޳��7�N�5Ҫ�x�݁;~۾}�V:$�ڕW\
s�lK�]J�s�ˉ���b/���͝;�>����'>��O�����~��ݔ;�7܈5�\��#*��n	�s�9��b���'$��YY!F΋��S/g��e8���L�k�b�3w��\f��A��m����L��ŦO[8���a�}�K�bAw ��#Q)VI�E|i%qt�>���s��,LI1��52��T���;����K�{��V�^���x��?d����;�k�~w�[�X���J��7�	]Bz�09�s>G�4{�(t�������[��`�5�z%*�߃%�`���%��%�_�����sL�o��퓌F?>q�����E=�/Ʌ��cE��2��<?�w�q�Lg�<f1��ʞ@sP#�և~�R�׮܇P��_����1�}h��1j��G����=�pz�����c�-8����{�*����U��A���{�AؠX�S3a�j�H�{�1by���3�x	�K2�NF������TI�e-������&�m�$.S�1�ڻo�:{¹���e�#�MQ�.�;�Ne!�O��|���m϶x�"��%���$�N�VOu��eC��v���[n��v�	'ؑ'c?��������ڈ,�j �jr�*�#�CS��%n�6����h+R����3���n/���5����#m_y5%:���K�Zx1;n8:�۶���6~��3q��)���Z�!�=����j����"`�Fɲ�h~cUn�&&@'��vt`h>͊�&��$�}@O#�!��dE-�\YS4��̎`�P�Ef�ֳO=b+׮ &��^gH�C	����.V�2�����7q%�(��v���N��]q����mQ>�"E �]�K����Odf���
btQ �X@]�g�Z�.I���.F�uEj�)Ek{���[���gmX�C��4� �&l��u�.S>M��� �2�$uk��"ƭ�����T�� .��w�<�0\�@;4��tz����Z�n�|H`xf`�π+x�9
���d ��Q���[��:Ri������)%����I�+���"A�2f�5�X ާO ��7�|9v1�i�+'s-�0�<wsm4��im���G��_��r{���a�����.sM.a0Y���κ ���Nk0��A#%���Q; F{�0��x;X��ڥ!��'?!�?-4�]�m8"�1��߱u%{�WLꥤwh�O�[kh;bqhV��c���~r���[XE4�-������)������N~d/�tI��8�ҳF�;�+���`=#�Y_�ʗ���N����6��qWm�d<zR ���K�������ü���z������?،��7?�kӎ\�=�n����|�F����z��q�gm��#��2��������?1T�*U�%�:�ӧ���T ��-����eq��`�!4u|bTNfխv�Q#� U鶭h�M�X����:�[~�#KGo�¸�Yl��kE*p��~N��L�mu�>�Y����t�+�6�.�p�x)?&�X�^@<�ˌ]��t	����'�6���4R�Ɲ1u�!!#Q�$��'yF��q���{�'�ܓ��]U�{�[�����W��L�@L��{�6��{W�د�إ�x�^Ёy���C#���z������Vp�8Ȋ��
=6n8�8{!�W&��X:�@�D@���g����*���F�S�-����?yO-
��V
���A���:���Ίc��;�tvj���{p^Ў�H��,�n}���8=�-xf81<��?'�w�0TVLd,}�J�����P�.��α��4�1GԸE $t��I̐Q�p���YVV�Jk4q>^c��ݳ��d��8ڤSaW� ]�A�|�uY⋸��$hg�����`WJY똓O"�>��Vc�����^>v�e��{1?7%��,�cSrR�d��!t���M�J��,{���[��2wl܁s�&�̙gZBx.����V�R��M���T��F�Y؃���x�+5���#���*A��DD�DrЛJ��i�?�:��=��&�[�0v��|�9:p��Ԋ���A+�iJ���1��9�Y�V�țHi
��*�"����==�]z�X�'�-wX6��!tX�ǎ���N��aD����9�$��6��kk0�����A���I&����4�#�Q��d�ĒoE�SFz:�A@^L�2��%��#Y���;Rb�r��Q��7�{MO_�J�nr�]Ҍi�w����uW��;���dL�W��:��f��}R�BJ���h4ĺ�E�E��-�QΗG��h��\��(%��J�'����*��8�A�
�Rn������� !�$-��$< �D�i�Pܖ|�D�wɍ%����l�)bx��Q�C?!��k��F���k��Oz%Gq>�P/�*2F+u$t���2�c����O �h��r�\6i���Ds��駎�(Wj�'e"
�]c�t�R������J��)�k?����@�E7��*��w���@�Dn�@�:sQ��B��C }ݽ���QTeJB`���:KzYЈ)���|��n�a�0+Ϋ�뿗c�� 3/=���c1F�bd,d%l�"m�/��v�:s2��G�$W�c#�d۝��������捰}{�b,��.tR�1m8엣}�`Q6�.��K�b���W���hB���_m˺�VR_n���<�x���A��H{�͕h�vڔ�m^��p��׸�2����n�?7�~�G�rbTMC��ؑGN�������KD=���w��F��m�>��5��5����1Ym���� �(����y����1�n�+t7��~����3�J�q���p��XL�㸦���f��y�e2^�'4R�^�1�R�v���a�N�Z�w!�n�`�µ?<�ع��??dm�7�'����	�Öo��$�;���2�Gƒ���MG<��4J����hUR���Hp(M��T�R�����.��	�G���*8�dӂr`�rd�Ϻ��|�����u��<��4�&���BI��4��Ba�G\SA �h���Զ;�)L!ܢ9<�\$��U�I���e��<R�J���C:�}��k�����</ �T�OS'��Vc�^�}��"�������<e-h���f��>C��t��'m{�3U2���tۮ�=g��p�#�� �8�l�k���!�#@C��8� |��8��X�c� ����@t�Xмչ���������{j[]0�����b�@�|����0���.��5AR9�x�k�8���Xhb�����FRCo��%t��S6����ʡ8���%�g�9�x���왗^��6@��c�v�8��1�m����?}4m�%�s<���$vv���϶��[����u���/�v�d��g?��H��fOk�Z`	�۪*�`��d:�p`:��)]�Xxh2^f۬��	�}���NFT�@�X>��xe9�%'%��؅�?]X�DS�Ѷ]��V�6�5&���)��r`ڱ��d?�ȣ���~-�FN~��'L7~�zw�TV6l����0��[$2)r�hV���81>�@�=݌��ȔN�s&����/�EA5 ���V0|�(����q�S��nm��������Y7��[Ç�J�p��pNC;�y[o���$���*�C�EB&*6"ItFɬ6��ń���n�d��"�9�	=�4p��E܍p[��� n1��s,��O�}��*=�)����8�rM���Ha��hӀ�.Nn`���a�@9<�(�A�/+ƥ��4��gj�~�ɻK���FG�� X���< �c��N��ñ��} ��b'���7 N����?��HlB�P��V���ƿ�����F4�:(�'��-������lO�/e���@�~��N]��:�!���XM	2��Ȏ�O�>_]`�^�y�	Rz��#5`b4�$���9��V��]/�'���2�u�wk5w�@����d�:�k��R����ƒ
̃	���I_�l�<=V�Ǘ~Wy=�EO��8�by+aS*:��� oV>|=�
ׂ#0�E����3_�#��7ޠ�9��~�~�+(j{ྻ�,%p�E��.�؎Z<��|�چ�v���V�b=��ť�؋�o�~CK�ѱd'ͱ��o����E�~��V�~��7'��E��C�U������4�ּ� �;������/ķ-���׶t黸˧r���sϽkg�y:�2X8�����]z�%v�}K�W^v
�0�#G$�o~��=OAα�ݷ�/cl���X��؇-���e���t���\3	��=F	#[Y�۶�C�oIt:6��c�)�_h;��8�+ ��0���BE	y0[���l7�IY�g�%q�~XF��^~�e6&T��S�/_iv��e����AՁ.I
M�YMrm��q"vM�j�PyPL�T���\����M��_���;�\�g���}����2�!P��4_l�(��Bб����g�v!�i�S���]�q��c%� �s !���Z�i���7��{�X�9A��W����΃�F'[	0v�d�$�I|O���@)��8<��m�!]�����=;�]�8��k�8tFB%�m2��X��h��-o�pR���1���wup�a�]Y���S�#�W��`�Qj��ܣ�l�E����.��kD#n��Ɣ��bCT��`�h h�0�k:����Z�[S�����_{#����8��F��i-fզ��ؒ�&q:�j���@(܌V��x�5
G9��-�ǵ.�m?�X�U��K�S� e V�M�d]�`��0[d2�GXuBb:~B�-&[H�#��vW�e��J�NBxyZ50��7,:d���+-�$��bp��a܌�6���&D�m�Ҕ;��Q�#33�����_jG.�k��08�h݆u�m����fn �/�GL��L:���Z�[Ic�D+��.'b�O/��B�5�ϐ��t)�bQȥL�1[�z3��/1�N�4lL\c'M���E\Lv�*7&��T��Үᣖ� 7��t��Ȥ<%p�ɗ�3���q��W�ީ�O -p ��6$�};�t��I�&�+�q�'�c��P I��"�OO��Dbu�����,��]�Ǳ���c�4�#D��E	8�h�G�F+O�n�	dFG%�����&Qlse%7��m�}��Rte�#�)�m�ô�C�J׆�:0n�ܗEÂ _���T4x����/N�Q� )�
,����̊4��zT���<����1���i��,Z����S|N��>�,#u��y^�rေ�{��[A'[���y_A��:lSZ9C��x�_ݹ��+Uj�e���I��D(�d`v�>6+ =�p����>5���������Ic��
i4��몙{���3�29ձ�o��o�M�/1	�S (��ae!�V�1wI����/��pE��޽�q�ˎ�[�*Q_��(����klweݞ1v��ؔ��O���.��L��g�k��k�v��t�g�CmWQ����;��(3"c��/+������QX��b�0���� q͆M�JpyA&�$l�=w��M����y�v�����9�N��tÆ����>�]�3��X_i�gN��Ů���㏷E�����o��W܇,(�;;���p�E;l��aVVQ����8�4!
�/�#�%� �\6 h��h~����ي>��9-���WS���b���%ty�l�q���x_��c�A� IE3�L,z�Y�'٬�Gؤ�#����ïQY���k�E%6g�d��:��B[����1ᆭOmC3,�&6���胺o~�&��=`i��~P��,�E�n���?���^���� L���}���ĖK���B?��n�{�:��=0��<0��!�q����k��}ܒ" n�o������8���0���'���`�D�A����=.�m����c��z}h��x���#��}j�f	d!�!$̵�R�A�Z�G�lAi.%A���5ӫh��w2V����e�_�'��3M����iW�2��&�-�Q�e	|� {=���.J�Ř4��Z���^@T��0�>P��Ǖ7H��s��Ԋ�~��& �#<~�(���ͽٱy}t� a������N?s&9fv`?�|>>3�1m�}�7�ij'Yl����(�mٺq�0��I����t��g*�>vb�Z��]q��0kB�,[	�ҙѾ��G���.�)H��چ�Ѻ�k���W�j��x�-@Kg���tp�a�J�?�L!����UʳҐ����T��d�u�m)�^`��q�V������x�m:�:�0����5+��ɱS�H�u��ɱ��Z&�0 eZZ&,��B��\��(!�^�*���:,�A,R�FԊ�*��kBY��T����P�]g��V�O{��JL�j\WZ��
0��
��ނ`��ק���Հ;�q��Y��db�B��H�V�)\D^�͞���������$�G8��ڄIs�� RM`=���G �#�,͖��g��S%@�j̀ag � �4�0� �pcu���O��v�%.��D��Π�������Y� g>�0"_�hJ�1��du��9��Ⱥ�N�%&Mh����qX��)���$(�X3A�-0pM茺��'�_�Ţ���y7��ć��8��6��pBz�Z�M9)��,#`�5�&�΅� ���:���bo�����X�����9� K U�:Sv��KM^e��G����S�K�ar���r禍k����@�.�Jta�hR�b�`��*i��g? ����ف�0ƙ(�y2�l��2�Y��cZ�K)�5!�,�rt��x�yB<�������#?s����� ����7|��h<���6�3�8Ͷn߈m�G4��۵_������w��㏲�G�`+W�#Q�]����D��_a\t�]q��O=��ۥ矁���1L��+���vl�ᘱ����z�]~���=d�׬��	f��W���[�W_��̛M��6c<�.�F��#?wPG�9ĭ���d�m���y6MY՘ss�i�RyL�g���ZH!c��l�G����#���?��}�F�@��#��۽�49��b��65�h��O�~��1��:IƼ�N�~`�����,�߻*t���"-,��;�k�����v� �����j0@ژ�\�mr�������z��C[��'�q #�, ���?����J����`��{��^��x�z�yׇ�8����;՟>�(�.�����&pa"'d�����>��5��o�E}*AKAZ���*JL��j���(A.��,�2�
�\����M�Y,�&	��k\���fѯ2	����f͟c���ݾ�	�@�3����~��\�bʝ�a��a2�~�&���ۖ��[�t���
�ePǰ�'+{8;
k��PT� ݒ��>@av�G�2ԉ�;q�OF/Q�S��nѢ�\	/�|���P�8&�d�'�w��-6q�d�0u*�A��>V�0n���N �iԐlˤ��K��Y&���fN!F	[����(y���ig��Wg��oe�!#KM@�,b��-�UB��z�0�5!|��
w�4t �R �Pb�Ā�j��A<	��T�0��N&�n�����nFƒPE z��-��U@�� �8�a�6�h%؎J,641�㼟.o)���������QO��������-	���6����68��L^;�a�@��mJ����y�SYQ &) � �L����+�A��$|�:f{\��Sן+ǱE,
��D�.!�N8��P�ӭҵP�y`���2�T�]�uiKt��<�*�.�\�d
���@��fɀ!I�];���J��)���=�{ ��U�\�4&�K��u9 `����5��}N$�iX�@�ǌ+�Kk���vU�e+���D����ڿ�d�f`��M#Y���$)��F�5��*�2"�B���{
8J�#qu8b]]=��&J{������1��T1\� S����D��3R~Q*��5���
1���b�[Ak" �o�&<� ��N��YQQ�vȝ�y���lZ�����mg�|�B��߽���=��)#s�<C#�4W'�L�a,����VQ���л�ڈK���� �Q�ۍ���Uq��돒6�eA.�@�b{�m��	x��;��tX?|Ɏ�_���Ⰽ�i���cl|����ⅈ>�s���=��������E��\U2���~$�4�v�	G���L��6�E��<�F�Θ]w�b����f���e�@K�c1�
��U��FP?{�����Ǟ�Uk�Cbr�`�4N�ӈ�A>���u+^�X�¢()9�sU���X�x��d��k<�}�Ø��_�Bs��m6o��kF��=���Ϯ��Ag��=��K���{]����r}��M��J(k�����+�z �_"�?���4�����<͛h���{N( �Pv�M��~ �tTAf��y~��}�`���`y�z�>�؂6G���_��3����'��CA�w,��;P���1a�Ị������HIA�7L$Q=є9q`b�&BB=��#���p��,�|}`�Fj#q���&|{�F{��q�g`��"GTw��f �+ȲSN;ʽ�閒Ym�1A�1�v11�tRb#~��|#CZA����D�#���>�2�J�o���e5:�7*o�����f��>}�l1r)�Z�wnن�"��/���j^8���Q3IubF��$���?�~�!����@�瘱��}'�� ~T�]|,Ḱ{��Х�ľf��(��xe0�w6KȐĽ�50���@7R
D��]����x$�n��E f�4����3��])Jz�0&Fr��l�����S�����&��2�3fN� ��n���竸'0 s?%��>JʰHрu|�����8$���]�v�N�N�p�g'�ֳ��U����6�ro%��'� �В���t�o�+����>D�Z��VGb^�q���C��8�P�0�U�7� Ez4il�B*� @��es��8\���@�X��4��Y�uj?�^�������KF�':��<ia��V��شd<��/p�r��]L�z�Įґi���ѵVO�L $��AN��j�d�,Y��hWۡ�F�cb�%us����q�D�]��:	%�ҵ���6��{Heu�M�i�I�ԯ}�S9�6s���܍&��iL�G�8j��WO����u=�Z�%�[f6F��8J>}:n</&�R��euO�z�Z�Ɍ���%T[���a`�Pgp�J�LXh�R �.PR��@�X2�z��K�qC�$�0kz\�5N�#а~�:K��b`��ep�dB�m&�%v�&�B��bc��{m�7>��r�x�5֕�����X&#7�����c<DP����%��T�]?%�K�˕ԑFIT��[ќ��{�x-�j�΁"4X��eh�kG��0��,Vu�$�{��l�Ĥ/�p�4�0X��Q��?��}�l'F���{�q/���{+���;w��A[,��rL_��J���~l��=����[s�]z�lh.@���4�k6�kX̯��ﭦ9�1Ll7������&��I��5cb8�welYz�u���T�_���č�<�1N���Ǥx���Dx�c(�=�����@��P@�=�?��'i��W����/��`� �R�y@�I�L��X����$���p�Bu( }��8�s��?o߼c6�5pp���w�������P�Y��H�T�^��&|�r��F��Rn��>��$�|�9��1�¥Ux@+�n�(6nNǌK���4!�"���dJ$�����*5�?�('����֊JJ�ζ/� 	�2�Z�F���M�;��h=�L�rFN���9�*�8��o�d�pž���'?��M�_`�}�B{�����{�v�O�oS'�� ��:;�J�)!�T�g{a]R���^�FҦL�ni��Jz�*����\�{l��2��p�}񋗹���}/���V�fuC8v�>bɱ.ܻ�<���:^,���^�`= ���D��UЬI��V`VԉJ	 .�kD%�p����� ��u��v4K�$������ ��IB��V�BTJ͡sI+v��T.�^I%��S�� �)�s+M�W��Z�r-Gc��:uE�R�cz�D�e0~M�?21A*`�I2��'&��Uv�����&��#*F`�c&"J�n���g)!�~���U)!�e��]V�IW��f%^W�J"]}��(H]̒��bұ2�=m�sx@E�bY�mݍY���16v�(��bm�8��%�ps/f��\��4�.��������#�k�N[�n��&`����& �Ғr{���}��9t�N�4�F�ěJ��b����]d7n�~(��m�η�cGZ�g����r�|�v=�k"c̴)Sƺ�~u���{���x�v��cK(k���D)�oU�mٖܺ.���>;r�B<��"��5��m4�<��{������;�	|��PЋf���4�&)=�ED�J��Q���/�\��$b�S�U����6���<Di�}cL��m�
#x1_����P��
�:t�c�T���c7T��c��s!�X��r��܋�ֿ�S�p��^����ˀM�?��0��޼�L�%���������,n�6ľ��a���O~�U@��Ӧ�7�{o��ka�:PT�65��T��E, ����I�����b f����s[�u�Ԁ1�d�^�� ��r^i	6,V����m� ��ȳTWQ�ֳJ��eܶ���L�[Qdu�o�+��k�v��D�ҩ"���[6��������{�K.$��ő� @�,�O#������m�M�8,.��o�7���F�O�X�xh	��l´�8�ϰ��S;�mkKF�-n��\3����P������Σ-j�Q�ǚ�'J?K㟄H���y��&�j<��~޿�L�<��I�Z��?��W��p�5��� ���L�ဘ������_��@�8��e0��/{��@Nh�8��Z؇;��c�eڮ�ƍ�k�[�0d�Ȃ���0���g�M}�xQm�@V4~^��C\�[gg������ڷ�S�y��>ڦ�-w�p~ֺ�EG,p�>C�~q�ol��Ev�%��[o�jo��~�Y6c:��
���?2Ε/�N����0�(�'�k��k�o��w�a�M4��V��V�Mɲ��E���$�s�\V��7SS�1��_�|ˎ�q�M9��`��G�l�R;�8yqɝ��N�)��b��U�"v0�d�����Ӳ��ȼ��r{����ekV~�ׇa+ۂ��V��¨$�W��饉җLVGci����"�8>¶�5h	��TU�Z�4!C�)]�Q��b}䯣ɖ!]qO=q� �mb� �v^bL�.�3�7�bH�ñ���ꔩn5[��5&�rD+~8'?�2i�8�La��$��>��4 _?v�g!��>����R�s�DĤZym%��%���n�T�T7^N��t�5aKK��J��U|:��U��Q������Z���D���2��(�*Q�I�tԖ�0��o�����R!�W�z�]����~��y�}�{�ٌ���40���Y��on����>��\{���)�*b	&�A'�[X�܉ȺV��k�J	{f`���-�s��︋���6l�h��_ؤ��$L���}��۝w��$[n��v�C#�K� ��[��랶?���hw:ힻoG�=�]7�|V#ݎ�쮻���G�>��*@p�ɱʦ*[x�|�{��gx�V>��\c6���(�85��5kֱ��afZnC'-����Z��k���LOCE���XT��0���5�EF�_�CU���o�<X_+M�b�D�H�"C�TyB��1Q.h�M����犱��K�A�k��rz/	��a�0]UǬ����zz��.]7-?��*�/�ćV�X�[Wo��z��V��ݝ�z%�:ՀW�D��g�?>�}��gۍ��ǥ[��$�.�}7�7����w�ƾH��,>��75A��?%GV�fo������;h� Gr��Z������r^��qƫ�=�'+�g?�!V7���o�`7�z�=�ǀ>�R������~�.�M���.��5y�<�	��W�&��(�3���~��oe%�v饗�	'L��tR��0�� j({V�M��Ϫ�M��������J!8�8���p��_��-�D�r�Ģ�H�sY��"�˯A�[i��r｟�Ն�d�4����`g��)�s��W�v̩:���	��c��Z(X	e�< ������?������柸��*$�uC.��_@�+�����zeH?c���L��G׿�.�U��O]�~ Z��>��V����q�,�`�X����r�R����5y��*����/�� ��F��V�;�#4x�x��ͭ�P~��B�#��^��nO�'Z۱a��r��+R���Q��nZĚe�0���v+��c2����nh�����,�y �[ �_/	�Sq�3|��۲��p�4�Ʉ�I�|5;� ?���ϱbV�>��Ӵ,{��&�0�-93V�K8oǱ�Y�{�:S	3����@����C$LP=���x_y��>sV�C���v.���l��}�`/���;q�m��<�LJ2�w����{��R1�M�*c�5��T��Jb�8:ߒ`I�;u���Q�Fkq�Q�(	ag �)�j�ז�@� >i �&�FF�#&C�{)��\��k4�a�L`E{
�
���vX�&[�&�iPwY�ʃ�v[(�$3���H�J-���I��D0�EұX�H9#� �嫝G[hd$�+�-����y�6b,z8� ��)�u�$�W�T�����= �Q����8��K�����{p���#�{�ę֓ZiŬ���'��ش �zb��dۛz(��IO�p2,U+���H�l�%� �5-K7��.¥�3�c5�Prn$	j������p��\6J�|S|MvV*�݅)g��G���i]E=���!Nㅔ�2�JI͵�â�.)�`���Н�ñ�KY3�e�	�Y�~z�	�`ɣ�Wp͖��8�
̑4�����B�y��N�R�p���a[a�[yn
���㣦�X CBJ�|4�`*�[#�)�<^3A7/6*C�!�OJ��ˏ��T�W�r�d��^q�K�rO54SB�Y���3���֮��q��5�¹&��Z����ǂ��W��D�����QJ䎮�,��j��뎺�3�$���e��Q�u��]�b���R�Z�]��F�C���<�4��SU��^�A�F\?%/��G욾�������n11�vy�U!��4a�)_t�*�!�K����An�9@�ԛ�`����؞�����k���g�=��>z3W_~�}�ҕ�==i+6ͱ�^x�����a6:3��l�&�+K�\�l8Bא�
0�1 V��Ҽ��xo%OH���G�.l�lN�a�*��d#���JΫ:��؇V�$��L�V%�&��tlTy�_V�4��ǵ�{Y�&�1w �� 6:��Hts˂�F9�f��:�s _-��Ӹ� �M��C�� _Z�V&�Ǯ�p��Wٌ	�l,�ڂY���_�W�]��b1�.e�Y^;����;�R�]jz� >̝O�p��+c`�zŌ{ �H���{0��*�5¿�����`0F�_����>k0�
���8��?�*���_�=�q������`�,�y�_��ퟝ���P�q0V���������`��c�� �^�18�1 ��9�=0�ק.G�Ji C%C�_�a���*1(-o���SϟN4��	���G3���5�hO>��FN�mEhԹw$TuDVc�9v�H[�v��n9��&�D�
�`��L]w��<�^|�dR�$����������"���V�eu�����c�i�q�XTVRr�c \��R;�ؓ0d�n�G�Ph�����3O�s�>Ӣ�B��#��6��Ȥ��Ŀ�&�75{1������3*ˌ��bB�󭶤�m�c�	ά3��DÄ�0�́QɆ5��jD�J6��F��H� u��_���iRP}=����� a��SN'R�%!���xʬ+�Fi^�$�u4��`7�B&��8㥫���M"�~JD�t��N%&�XސQ��01M�@�8]u"��E(s�@le�aJ8��K,f�L,��a��U�I�/�:��������U[��T��&V��0M�EYw��JL+ �EQvQ��|��u�qQ�.G!��LHa�.��8�%�5.f��������D��k�~�V�wY�Ȼ���T��?���t�&�sݩ���=b@n�ӕ%���H���F��S41�^UD�N@��֌X&r�T�e�e���Zm't���&YZ�hk���~G�M�8�ǘ�j)9շ�ߺ;a�aC"�J�q&eWS=��.�>���WQ�g�Ȧ�е�>PJN�k�t�Y	���6�-�7��&ei�:9�ݚ�)w�dC�U�\ā��'���h�Zد�!� ��r5�y�N���p[���
K���)f��LX�n&�z�+Ջ�����Z���А����XS��i�P	��'�Z2��6,	�;(�%�� L� rMʙ�َ��@��C���&m�@�7�
��4����$���H����v���8Z�K�R�T"��6";/ߕ��N�e�<��`��՗]�tO�%0����fW\p�=��ۈ�Wv=��YI>eg�W�ɩ��}u�Ӂ%3N�("Z�&��L�h'ITĀE�������D�`�Es��W�ǒ!h���) �T��Ή0˃J�(u�I��\�H���@*3P�
�r?�ڛ�1�%}@^��N`�k�;���t�ȩJI>��Q�4�,`:s��=v�`U¢/���n2nU�V�����Y���`�$�H�d��9��=P����ݥ]���Qk�x��d΅�X;��〳U F��_���A��/�+C�J�J��{O,�$�x̓|���P6N��p��S(�� �`��-����Bپ��?H���/K���?L�̙�����s���;�?��[W�<ؕ�1�;\S���y���� 5���44(�ǣ��A�K4a�rFS�`����	KPx��M�)3�[6:�~D��hE�ϫ�l�d�����hiF0���$�Ὁ����b\�j���n7��JOm��խv�QKl3z)�Idڂ5ś/���e_��
�Y�i�w��׮�%��$Ii�����a�fPnQ'&�np^C�hVf.X���~�[��cW]v�3�Ǌv��/Z5,�pߟ9�J)�VCi���Qj�6�p�3�j�D�d��{Cڸ ��r������V�aZ��@�x#��]��F;�c�[q�OL�) �(r�¢7@�g�> �eYݭ��;�$$�%�DMDhu�,+�%P�~V�LT�i��b桹�v,
?m�N�qc'���v�B#~�G�b!���L�����z[ X.P*��<�����O��ܠ@5�RE¼��n���t�GںM��U[lLW���l�_z��0 �aR�p����2@��2&ӳ���D���Q*�Kb"mRǦLW٦@���5�����W4ٻt�Q�j��(�<�&ؙ�{���ٹ���]��
w?��SL���EV��D����t�+ht3��#��W�l�8��b:v�R�/�ieB��,���k:�*v�c����M�J�W�hl���^b-a����V�n�b�bw"%�*���l ��*�0|��X�<���xZq�Bel)�����0��7 ����z�VV��h�"��0?8�9߯5;�l̆b۾� ��@ ���E�@�M;�]�y��!rG��� �2��+�_DL��S�"�޺�g����EA5�6���sS���t?),� \�N�N��$-3	c�N%6Yz/o�_�J����K�N�+�aG���,(��Iسk^e锓aYawd0e�|�T
Q�u��s����NG9<�6o�k��O����cX� ���G�I)�X�4���ڽs����u���½W
��I���kY������0��nW��=P���t��r�o�����'��so�1Q�,:�4U*��Z}�b�e�5�F焮P�]e�t���Λ�ʸ�ad���� dS`���<u'�s=W��;)c��4�r��y������������ZQ�^�c�)3��r{.v�v��W'�L���	��IN ����x#�@�0��u��l��x&�L �5��NV���P0�+	9�㕠B'�>�����/�b�n����&p��&k�1�y��/�z��1 ���~��C��e�C��(z�p8
"���ݟI�1�^��{��8�������q�1X��S�����gZ�������uh����i]´�e��k����-���c�eQh���͍VW��ܸ\����v�o��fWd�`�t�åNȿ��Ov�Q' 2^`�LtIi�Q�x��ev��s��j��S��)�8���˗~���k�9����߭���2K����3��۽ö�7Z#�e�����L��3�:�ȑR>~"LL��Ty
�����,K���`5~�L���A��lM�}��?�)ƪ7���e�"m̨���GI�rY#��n�/��;����*��o��' �bV�=G,d��a@��
qn��Y3'�}�ȑ�D�e�A*���ܝO�{d�j}tH�{�:�%Z��_����xdR���`Pl�lЯ�4� t�X��ᙶ���)l��#9�b��,ݢ:��5Gs�+��(*c���3��{b��{,�r��!� �D���(f�ey���g$�)u�U�����腱
V����p�>`���~�#���7̑s[oe�%��Lٰ�	����d�/�#V�wi�� a�6�/u8���� �}v�_��m��qE�u���Y�kPy�5�jՇhT�%3�~�X���5��o�0q�D�Qj��g���ed�D �f/���6�u��,'tl�)q��"�?Et���V�@b��.bX�V1���86�	�ח	w����ڍ�'�UI
IçZ��ڛ+��+78E~X�VՄ���J�%h�����\+��p�@�<O�M$�p>T����u�+A�ج8@��bI?`�s� �c�ڻ�c������������~
m���6k�h�2`����\�A�@+�Q汝�~:9>�hUΎ��|�}�Ѫ@�:s Y�����8��K�U���`�1�ė����p�}�x��Yey���q�'ql
�ͽ2�]1)�ʢ���γ�SF:����W��
#9�lF��1��� ���Y::�"�VGM��b�<D�c�z � �>�=ݓ	��3O:Y��;����O)� ����7ʰJ]��a�!���$�"��:��]+=�F���l��0.�;�Nt��(�^%MpQjuQf�pܒa�d�҆�u?�>`�ٴ�k�~�[(�-��(0� s���\7&L���9���f��lWf,:�&UZ4�o5���?���C�O@}æMV\ZJ�zC�RIP�`o�il�CC�ɾhR�y��ݯZ�🚭n��ã,�Ư�D�M�~��M��@A�P�	���������'��,�D>�c�1uz��m�L��ͼ���i~6)��j����I $Ѕ�o�k;?�����3�9=�6z����:���3�0���w�$�>���5翦���Ԑ}����2a��$���j@����~&��i"�S�`�]+9L#c��� p�b��
 ����QD�A�?ŭ���
��m���\"�VR�BH/+���d����.Fg��q0T�j@�ʠ)�����w^}��s&L���@h���aO?��n��gΣH��8��DV�g���p�=���L:�/!��a��.�P��Z6��]ۗS��6Z� �m�lD	a4��]����k��D�gp��ѓX�Z*h�߽c�ͦ���D W�aO�tB1��B��c�� ;4u�(G�oڼ�B2�<�s]�ۿp�	��F;�N.1��+�#L�n �he_%��.w~JG�J̆��P:z�RV�)�J�t��R�;���<���;��-�I��n$V"�����n���OX��tס鐳;���;�*ǕPb�3��u5*�'�v��l������㑕�k1LV���R�?+��d����ǡ��C��D����I�L���Z1���F��HM��YB�K ����u�ɾ��\L���Rl8�"�E@wG#n�����2��L*�_���wO'��p$O/�9K_J&�rld�J�, �T��X|�y�j�F�Ѫ�dG��� S�����AeѡrmbJ�R��ڽn��"��>�#�0�0`��،���G~j@,!��k�_6�	�V2I�RyIݫ\�r��\5�:�ᷗ��klL��]��ň	�[���0�T1�1) ��L̑�Y4ts~[䳆.�������|V�h��y��˗��S*Q"_x�ɖ#^�XOF�\��@M��W�Ka�*�)Ҭ+3N������E��sp�W⃄�z�b�4�Ӏ'������Ĝ���%�g$�����sTU'�>��ńɠU@-���륟�d1������'/�$��������|����/�&zԾ����:�i�ȥ3�{�����<{�u|>�.w��d�Υ�[���֥�	n���}����຀!n��L��:,���r����茯Y�$%�%�J)��ǵ##\e+� ���.U�lU^U��"�t�j�˂��~mmL�"=0����gE��)+ku��N���-��W��0���1����U�3��׭�?�{ݝEήc v��#��r?��[h�r�g,�#fY	*�~���*�[�C�S��i�"�<�3O`
rBY��_�d�ʹ�ľx%+?8�:?��&���P��s���~��M�^y��^�_�~����=�g j0���������X�1? ���WB��;�
�B�͟b�B]���;������^��!�B����	Ӱ,�L��a��us�3�UT�AbdZ*:��|�}ܘZrwc�����E'b6f�IVΪ�����U�(�g_x�9�K��1���a�Dph_v��VDd
���s���Y�`f���&,�x��T�u%�46"捦,�wj�'�`㪕䥍���`+;('����[������<�ZY�5�3�@ܔt+?��B|:LG&��
`�R�]������Yq��W'�X:�����r&�ݔ�d��lY	4V��%3*�csm�c�� ���Q2T҄�����Ȕ�.�@'`��h��=z��?�E���a���*<}�&�0B����Q����E�3��ilr����4�BR�`Ҏ��<��A+!\���c��9�eO\��^E�4����
���E��3iK��+��)���@�����W	8���\��;xYi�&���?1���K�o����C�������Q�g�4N���l�f[<�Ur��K����NT��[���&�M2)Q	CZ2�س%����])�0����q��q�n }]��l�.���|�%�
��q�n��@X�~V�b�4�����ہ��k��It as�+�`�v��`�JȰ܌׎���ޏ�O]Ě�z.19C��8������a�"
���V	���E��;�Ʋ{��O	�����ʌ�d�p�0���c��Y��]	��)�0N�0�"E@[�h�L�1C)o�0\��c�`� �:kc8M5VBsHe�,:6#)���07�S
#h��{�<����?kSǏw��a �G��t�L��bc5n�D9V��p��1��U��T�=1�2�q~e�G�20=���Ps����8K@�&�d4�b�5��(,g����2�ǲ��
�CR�a%qI۰�ȥ�gڜ�����#�/\i������;��� IqXvT�3/�e��p�Kvx��Wa�16�E���a1a�q��(�����E]�\x��QFM:�0�a�����#Uhj���1���KP�] �>��q�%����JF��N{e:�Xy2w��c`�@~缍�{O�vCc��'ԥ�LIV�Q��$�`����M��8�v�rkMQ	�Ի�1;���
�
Y�Ds-��
@-Y<�1���r���L� &0���8�J�N�V%��Ռg!!�I
����|�	[�w�gib�dF(�>�'�cߗ��3U���M̃� ���Il�ǰz����i�B��,���?�J����@��~�mB@hi�c��3�.��^���e8�q���p�E���K���0��򳀞�L�q�o���2�~ zH2�m����cW���x����[��8��h��A�ք�j�'#()!#"s?��C��=W�z�=2��T躊C�����m�-Zgy���{���<��x!|�Cg�k_��l۹u�����ZI�>j2Z-%5��Jc1���}95?��<���6�,��%0������^y�9ص-h"(� B���s`�a�R�b��J@U0z�s��[��悜²��gOX��}��1�C�i+��ifUG7f?�J*�|�2� ZdF2������6,[f�W]�ae�kW��I$gN!�v�ccCX�f��d�D��߰
2'[�ZϤ��nF��10MW����5u&�M�i�N �*w1�����C:F��`�����5顔?(�(5���n!P_��i)�9���te4
H�(����X((
1��]���®�N�u�!���K�>F��	�7	8�k�p��0DL���T�I�R���c�v땕�J-�n�T�F��2	�_*s�s�t��sRl���َ�ed�]~�����߳ES'Z)�鷾2�n�e��ُ��Ne;xV�L�bE�kGGY�VL�b0 �>Jw�L\���a�(#Ic�<�8���λɀmWɤ_
���$a��CQ�XBՕ�(0ߥ�Z��������a<�� =h��8�e�$����#��mΣ���"��	���M|m��"֏g����BC�����u\�c��	�Yߢ�4�(�Hj}�Â �Z�ql����`E���
ߩx�:"���p4C*s��Z��VP4���Lj�&�n����������W3�7�M?�.��^{=�W����@"���2�TSJ+M4s&O�����'�z\����)�	,�]�J|�yk��2V�7�T&�v%�룟j8��0[��)�D�+�!324́�N�&�W8��_4n�����"�7��k��ٲj���_l��|�����G��g����,�����~j�-����6+ގ�3=%E0Z�t����X��lk�&�VY�+�K��{)���S$� ZTt'��|@�|9ǰ�a�6���r:Y��$��t8u�84^�6aX&��qx	\&&ѠBY4����	9�Y��,���TX:��0t�MX� c}�4D�x���~�GV��>�e8ǡf����H5��&�{h΀��l�SS�Db��M#S�k]���5`�Z��E�͜�����틆��z�:<���ѩQ5ȅ�eU�=�b�?Y�(�M��.�����4%��~`��{�7	�5U�<+�N�B_�����ͳW��|���f`?��7x`K?=o��ޞ��`6�%3��x�#������H(�}����1�﫟���<y����}�����{��b��g���B��x�n�Ot�(EDqE�W�Y��G` <|�/�������:��l_٘�PD-�u�7��?tI~j�P�C�oDJJZ�|d&���3'�1�&��/��xԹ�7�Y�6�D��5��dJ������6�����hs�g	������ә�~��5IȱϺ��{�}۰j���֛v���>Kfr��`��%�0�u ����t�톺ǽ+�f��S�2���Rn"P��B��[�r��4���\�x��|ƹv筫��G_�3N8���mf����VX�aW��S��Jw$�v��K�u���%bb��.��zс}�gb�Z�@`y�.Jz�,V�*�v3ah�O"�ϝ�\�K `P���Z�����w����Iڦ�,ʨ���g���_������h�:��=���~����8��i�K>"���Ϻ�R�`&^]u�隙��쁭�DC� ;�L����"�@3����m{�
�y�V)���{KUR��hI�2�x�A�K,��]��r!5���30��Z�z��+�f�:��ɡ�c����e��0^M���M�����cǝz,�1.`[^k*��qA�� ��0��# fUU{m|]qt��}�	�yW��>��R�3� �z��Š�d(��*�?��݄��e���|�3I�X;���6R���T�8lE'6&q�I�>��aрe#`���	kl��a;���$[��PTL�<�$^��X��&�N���ab��+ʊ`jaJn}��~�x�� @�Y�D��(���Q�{~4��� {(6Sjj�I�Ă��c�1e��S��X+�+6�`6�i�z���6�";<��g�|��U����X�=��뾃P;ϱy�@�v����*�Ny$Tv�ܯ�'Ȥ����P�~�|�������H0�,Pjs���s)�+�\l�|�jj���hd�*��co�_��p%o�X�E,�	�.�X0����羕'��咫.C5ζ��mC�?܅�߾]��6F=�ׇ}֥�w�\�bm���-ܰq�
��g�=���#W1���.������1���ko-�3&�E��
����c�1�!�t5��?¾�ڍ7ހ;'(������T��'�5�^hO���ƣ�=���c����j���r$�mݚ���U6k��3��ǟG"҈A�	6z�D����l��4H$P�����	3m԰QN�8b�0�gY��2$h��hG?Z��m����g����l<�v�	s���y�~ >�HX�lư�����s�Q-�e-�CH\X����� ��#����Z�	�Ϙ��O����z�.��BK`����M���lb-�n�������%�g�
?�eC�m���?�����������y�
x�����7�{9�Ol���j���w���?���\y���U(��x=���7�q��1�f���#x@<�]��7���}����Ǻ!��o��:~�X!g'QF`E�Ϳ�V���C2a��-�hw?�e����+|�@�E�D�h�������>`�&��K�;ו*�Z��K�_��f"ؼnP/�Y+^*[�F���K��[1ìi,VeХX�δ3��~�&vح��Ҧ��Nƞq��VV������Ͼ�;��o�S?`5�b�e��6|���Ͼ�/R�-���+e��� W�`讕�@,E8������9���?�Mge3y���o�g2J�`$���	�W^�cN;���I����` ۃ��{~���6{�$2/'�2��b�m�8�Gbp&�q �(�F(g5����N����`0 U��t�E�Ti�9@�)&=ɞ|�U{�7e��1���`��4jt$�j���;�Ri坞(�F�f�f�
��FD3eZ�Ms]���r=��9U7�Q�\ H%�`�����uK�\��g��Ne$��hkG{UcPu���(��8�
�f$�W��W��%&����sK�����Y~��+�1&7d,%�X��t��X�A_��bLw��βz��/�,p���=P^���:��-ء�"��3�1'X��m�h��D=-#�V���0�g���ؒ��%����T2�(�Rb
`���Q�[�j��-&��ڰc����~,.��w��.�)M������r1���k���6�,æ5p,"�m��舉i�|�\�ʪR���ﰿ���J �� �+�t�k~v��ix��1o������	{>Ҟ�5۽��N?}�M�1��� 1L�a�}�p���Ɵٚ�+\fk�_��{OLb�d�A�>�kJ�Cl�4^�n�	`��1��X�\�qi���K�=�}h�[��N�X��`�_{�O�\�j<`�$�Y*�E�G���2$�����~���NJ���9�2I�c[�j]�l��Rt�80q�O���f���Qx�Yg2>а�����8���ﲋ���Ƣt���q�_l��;�� Ý#p� �YW����3�>���0�Ϯm;�߾� �� �E���O����f���`�cl��R;��Km��Y��K���Ǝ�d!����50��f$2�E��˂/j���������`'�Y��j+֮���xԎ�H��i��<�L�>y��v��%%��{���1��e�E:�S��촺��-��/��u��YW�}�7�.@��8{Y���l�Æ�e{���v4|��)Ƒ����҄�KuUk���e�%,�>��ԣ��N��$�M� �ψx��=B�K~p�I��*�4��A��y��z��1�a2tNզy��Ie�P�
�����/~�
�B�����s�<6��"3ş�������>	p����󥙧�� _����Et4B7���3���Q)������f�h��Ϳ��9�X4[��	��?'tC�@�J	 ��B���b3�@E����`9��Z��񶮰7�,�Nݎ�gδBD��5�y�6��v��NC��(�,���Q�m�X��)��L��f�u@��K��m�pYݙ��,�=��Kt5�_<��p��k�z�q�cc�N����ho���M!BF"se6�q���L,�_��_ULF�Z��e�+�w����Ⱦe�x��j����Q*�����M�-8��sge�~���tw3��ݝҠ"�"b�q�㱏zl���-" !� �����_����|��������0������u�k]k��ۑ�u��\��7�_-�_4[.��I?���#^���{�4��_�nr��3�ʋ/�$g�쇣�y���6�u��x�1�j&��:0u�mb���y��M�a*��J>��f:ɼ�b-���ѷ;�ҪQSx	��#�K���^L0�&��m_$�:�4�F���je�T�C��i�Di�0]��A�����A�\ugڞG"�zK~�a���%ЭF���A���/�}�R�]�ث��ʾ��_@d+��˔�_�զ݃�� ��͑�}"�</�͙%�?r�����eƓ��vt4��񀙶�����S/53p;Fo�x��d�(U�c��>{Q�V��2�����O@�r	��#e��҈�j��]ce ��D>�=p̔�*+��P�<�+�R�߬`�)U���O<(+0a+C�/^j�L_&j-oj&��� ��43hpsEa&FŚ�-n���a���� .�	Y@Lm ����o���}�G�%�v��r��2hP��������"�<��ص��<��B:��aS1+�)��![wb"�� t�&�T���U�������~_Zz�O�������, `���ȅ�Ġ^Wj(R�z ��m��84�Z��ph��r��+���Ҹ"��ԥ]K�ǉ�z���x�X�!W���*J������˱��a3�h�jx�;E��T�`$ �ɚ�̈́�I�+�v���4^~X�Dbj@�y߁<֧��$�;��ȝ�:hhW�pm4\��F�Ȣ�֑hA3Ǚ�](��ǈ1����t��7n�0�;�K?��x{ ^j�=@�qc$&�f������3�D��a���g_�ՙ�]@�A"�"�>�Ǐf#	#�,����-\�ƊB	rKb|h�~�8�^NEAc�bc�B�,dp�Db�:!�h2�q4��Q&-AZ���p�[��ðiC��G�MnN	������+����]nFO��;l) S��zR]��.Q[�PG�5q�'g��s��y;f�gX�?Γ�����p{̷���3������c�q0<��h���\8�C;@��m'&�k�l�c�t����������C�o�����"h�\g`v���y��־0h�	a>��/�_a�AFF�4?z��~!� ����,��W��녈�Sd��a2�o�|����LJ��#����t^~�"{��T'����KWSZ�E��I��~:`�@��i�4�������ɪ������a$`G;�����Ȱ����zn�<��M{6Vh�Kg�O���+D�0S�w�B9�єcG$�MW�y���������* f$hb��6��k�ǤN�_$-��������TNnq�eh���x�M�c�~��SN(5�`X�@�R�}��I�d�&�s$E�N�,o~����@y�;�J�e�~�K,�rEV���v�:�����F�~�2�ܳ���.�܉f�Y.�1	��� >�O���l�z8e���j�i�hQ-:a�\j���(�����@���f ��S!��������?-�. f7V��ǘM�Uck�"x=%?�0�Y
���^k��4^�h�$��<��)���Z�4���ɮ(�j[Jk*d�́�W�e3��_�ڞ}�T#G��yRX.��b�]�����FJ�ڽ����1&���R�1�r|O�\2w�$v�!^���|����Ų3��c00q�Y�~��8VU��S���l��o���� g��pՕ�ʕ���T`�;[V{k���lS�\���۵h�\����q�)a��J�X�d�	�D�V�O��\W��؎.e��LE��ղ���̓'�W�"�HI��M������PzB9�+�s���p��,�O��=�ʤ	�d/!�G�~{��[%�N�k���(�2~,y��h+_�O?h����L��=Qn��R��R�'�cݥkw�Lq�����MWt )��MX7�;�d��R�Cm(T�e�V�E���S�q�Z�ӼC�k��vT7��5x��Z9տ�ig!�U��Ԯ@�m�tm�F�5�H�H��>�ˈZ��r�w���[R+� ��{b��ҭG &���5i�w'��3�����RvϾ}��%�p�������e�X�)������Tq<�.�}ʭ-tㆄj� f @���x�ÈcҲ4�Y3��CF��%k�Y:w�#q4���r\j���؂���1_b��R_���bsAC	��0{��8P��p�Kfm7�e�O�w��b%0VX�@#Q9`
��=a#irqeSS�&];�@µ8�RFY��B���3�f�ej����/�0����K��VXE��k%�������W��2�ޔ<����p� LA�y�v��-+<�Vz�,���mM|�l� t���'T���^֤�ܥ�`@��κ�S��� ��t[V��3x���d��y!kE���|n쿷3S� �ڏS1�sbaΠξ���]'f�.��:��T���~�8;:F��9��#fզU��[T`a�f5�5�ٍ�����i)BsG�J�@|}��W�%�/�tޔBaB�d*�3Ѷ�9�n�d���}�a�j�������ò���d~n2q�9��0������Ҏ��7t��{h�qdtWbWJ)a08�& ����S� �a��y���ԉN�j�k��q4�K�6���X���� �;�~���_�e��(~^d�|ˍ�l��|��$��c���cWQ��8�[LD޾�M`q\\<�q�({�D�X��w)o���wH���>[d�C2'�*��+w�A"��IH����"6��L�v6�}-���	7�L�3�8]�t�y2�K9.��O�`�#yU4�H�v6� m��4�@c	nv��`Z@�1��!E���P���k��F����R(�}8����6����C #pG/����2̑CC�������Z�������26}[�{](oz��k�I�����ɑ�S��ǟ�
��FsS.G�^��	��m�*b��jT{��V�~�� d�����Ar�w�J%�$��޲��!��a�`�j�΂�&S�TP�eG�[z���̱��x���
z��&W�=K^}�y)JK��cF��B'K�C�M3�,_��@�+`TL�/&%��yx�x�����&����C���o��t�~��
���h�Ǵ�`�|���r��Ζ1C�qm��;=伙C����4��x�,[�[�,�.O�z',��;T��;A���Dʘt�}�v�� 8�W�S��7]%=aw�]2�X�$���O>��'y�G���"S�:S~�xT<�8�.&v)��`��Ѓ�]\���|k8f��Р�X⃎�����l�d�3�%&/@�� F�K�Lz,(�`8=���E��e���Q�"a\]��r�a������+���ܫj�`�yƔ���W��ʕib��Sa��؛�D/� J�$r"���N%�"GF�#c��'K6���%�|��6 ��K^z�5�.�5��]êq�a��T�\��&��(�:J��]H�BDlo�9L=^at:Fu �wW�P���7��`QII�M�t������d��Q3d��H(�~N"�՝��F�S~%,6�At��~���}�%���@@ߌ�@㺚��u�M�P�9�-���Ox�/	�X)# ��� 5!V��xܹc�ӟ�0+��V/��q�S�T,���n�F݂(h�lG�����0 \c�T�� �&�4f��];���do	������^
�&x�y�0�A�}��o�;�B�S��,���ul��ֶ�2(�,؏���9���0;`��A���� ��؁�3 <��3`��s����]��s���ά�}�ґ�q�}�o��S��6�{�����ЪN;���0%JK�=~X����������),Q�*7�WW]9���Y>��W�	qr��i�3�V��2VP��͈_	�e�<�{gي�;�s7C���2e�dy�W��H7�����2"AJ��(�N7:�LK���|a(Yx����;'�C��?e�2ʃ�YG	�f�{_Jh��u��3!l?��5�%����<�1���,ƈPW��R��z�N��N~��hR`���S��Si+p�:n��Fqd�9V�-�U�09�Ig�]Tt�5T���[��$���Mh360aU�r�7f��H&�E2O����iL��%�my���%�6��3H���>�AF�5����be�L��z΅�:(�B^K�	H�
x�D��2n�8��'m�ԙv������4_�����XZ'�:
=�;�,�L�.@��i%3��hs>���yDx�TX��:D��eD��SE��d�`�WX�9�1�
��A_�-O�s��8��s�{*��s�P(���PFJ�������U8�Y�8�7W������%��f�#U<�N��Ң�?���S������-о�v���ƒZ����i7��
��(�WS�:s���F50,K���(sg�+��"kݪUt!��Z&
�������4��ǟ��5$���IcxF����V��URӹ�x���K����a�$	����a�2e@gٴr��?f���wK�� k����ze��U�ۼT��������W;���٣dצ-��;�Rƭ��.;�R�vt`t��yr��R�sPb`�Z�8�`��6@�.2b���K<VD<���0H�b����%��*��ʠ������姃�;��z��7L�v�Zp�eY5�х�d�j�`�H����g�����j�W|����}�7��j#��@z����4�;��j�7T\^��5.�v4t�J�������k�QfF�	�Vӱ�G�\�
%�NO����} �n��c��O��_|Q�Kb�o��녿ˡ�R�%9���� ��С�X��� ���q��X����J9����ZEX�kp��|��!��v)*��� I��?����B�,��z�EF���IZ�����Rɮ ����6��W��ڤld��WRhR���L�*7m������w@Z�j�8>�>��|�m[g�s"3�9�z�z�	����R;uV���)�WӵL�Ud-�x��h:�?�t��4�Q+>G���pi8��@��v�c�u8�״��쬓�=v����rfu,F���Ϸ��-�f�iV����H�,��۲�-y}�L�$;�t;v@a\��A�u�����1�vpc�b;:F{'fG����r�3��߫�DG��um�����c������9�-�j�lV�1�_j�t�gDXp��������]`��ê��*��U��*=�{��D?5(,Pvm�JcX��Y�$��E	,R�8ۚ$4�+6�ҟ������S�S�.��!��F^|�=9�.(�ҋo~+��]���ڍg�d�2p7Ԕ!T�l�J���.
��"V]�Y؆��1s��pu� �DQ֌����3Ϡ���<�M�aӖJ��e��=�S���ڳp>O�[*���k�EW��h�b	T�D�oڈ���]���_.;w��Z�X�#ɒWR!~��I8D��b	,��=��H���ђ�������[o<%e�/��[Sd��Qh�B��u��߸针^ǻ�8�/�s�JYF�@OO,+ F�(y���.%U�AÃv��2aW�A'M-0$�O)��&��b ���A
���S'](oi&xE6��6��)Gsp�6hxdh�T�RX70�Nxf 9q7��`���Ș?�h�vZ�J����͇�m8p��j7i��	��U�eg�J�tW�X�k�%���w0E��B0�݊ I�"�=���tb�i<�lӎTͰ��a��I��pJ:絑�!�^7���+%).\���+;��Vü�9�$�ǧ禡����H4��D�Y?v������_d��Q*��<� ��L\M�G�Rb9��0�rS�OO*gI� �%8ߣo�(�᪕呇o���˖lY�l���0Jn�Ŀr�9p`�\t���yθ�y�q�ޱC�#To�l3V<_UD<i��0�H9��']z�IC��OÊݡz6ʪJ�h Z(@ci�L���h�K��Ug|�+��!sDAҀ�V-k���>Y*�����[�p�¤#U]����C݁a!5�GmE4:��f�����a������?������8Q��O���\��,�?e��a�����Q�%��M�L�b:�:l1�m�B�ٝR\9��8�9% 7M��v� �j��8,M�#���Y�a0�$���5H��#�~r�c�ݠ¢��5L~X�F�����Zy��_�~ �����sJ4ľ4���cG����aýe��4��\v��G��r9�,��ܻ�x���#���?\,�4��)m�x cX\��2l�0�/����U~��"m_	�՛JF��M<'�ǐЫ�<���<��a.r�5�K���2�9 �v!�t�F;U�b����Ş��.�m��97���#���h�hWg���1��\S��Ck�a��X�Y�N�'q��3kd�$�v���- p
�mA���%�ӱR'����v�c/�c� �s��X���A�T��__g?���\G�;�^��Y��3mvPdg�����`/3;�[ֿ;����Y*ǿ��':�0ݦsI�:G��������#.}\]�w�|<iZi�w�$�K�E�񫮸\~�u7� L0���B#E��:T7����U`I7&�aj�n�

1�ܳ��d�?ԻOZ���f�G�m��4��:��D�.��d5��@ժ����h�\��kKū��XQhk5� !����A�d��=Г�8���*��Lzt���u4���$#+W�O�D�Z����hc@�l�ZJ+9���� vR�kHF���@��S3�H�j��y�嚫.��.�+�z$7��,�|Y��|��.˚V"w�#X�b��{=(k�a�PƄ^��+?��;m��8�����$��E�ʗ��ħ�`�HI��;V~���9��<��oV&̹`�S�z%+���$�.�_9Q����mD:�"G3���8���.�3�c�1%C�,�/	�;�c�P��Og�	�s�P�8��﵏ʖ�R񦣰��,����PC�+ۡ%<~��	�j�c��ن�vV�� �l�R��rQ u�Mnh۪5LM� %
�tR6]�ڕ	�fz0���7&�ґc����NL^�]��~ePڴ��LP�P`�B/5�UD�@̔!@�&k	�G���'�����zR��~ص� �J���X�+�P�^H[�s_VVp{�����}��N�it�� X"����Z~�%g ���Y%�d�o���o�_c:Վqou%Z���R&��L9�]/I�0|���/�\s�,^�N>��s&;��wM�~���� �4�؄x:�����_�rt\F���, �ԏ q��FI&����{Y8 �`Kx��Z��CON4�� ���2k�b���ED9c��3L�~6 ė<�Lؔ�4� V�����	`�WǤ�%aWBn,V��qg���I�%���jnQ���u�>h���o����"w�D��O�*�u�t�f���$�9�gNC�u1�R�Y;%:Mi��۸�"�f��+�X�UWxa��	�R*�}Ǡ�:��-�<\�}M�8�w�̚>N�͛s�(�<�/9�� <f�9_u��8}�8~���--*@7���E����;~m

��`�S���xr�3�~�ȝw�M��)��n�����DC���o:��0"�?��`3��D�ryH*l���(�캹��Eq���S��oxr�\r�8l� ��e�/Kѽ�2	&��5<���4]�q�m &͟��0]�bA���<#ޔ<9ϩd�j���?�Iw��6L~C���e��"8�R�J=��� �����,}�g��l_M�:�:�u������X���:bb�>Y������̬Y �$�);H�3xv �C�~�Qy�d�����gg�:����3貿��{����m?�� �y�.�m���X��~� k�������}���d�<��8����fhi��ҥ���]9R�4��?�{ ي�P�qt$��WޥYBv��0�u�@#�eͶ��C)@�% ��/��}T�����JVT���J���w��&���'_*6�て�yյ�x�
Y�f��0ڿ��Y5	��ET��Ɠ={��N����0��Z:�ԙ;��z	��[C����Ȫ� ���!6�>��9a��U�2q��xJ�m�����Yҧ{w	#ʤ�	��UNUI�exv)�C���t]�`*֘U����U���TF����bY�	jg�Y���� w�;=)�� �4�I%�	}��LI�+ư2D>��W	#O2(�/�At���d��GӁ�o�|0�7V��$��_X��T�IS� u��V�ҝ��
�z���ȭ��O7a7�M�#�h��%Q�m��/�/���c��<MG��A�4s��~��C���_Hj��Dv�+9u8Ϋ����b�\5E�L�H-�T�eG\�)�a��o�珿M�IEڪ��Ҡ����_�;��z���&����[����9�9��)���h@�~9>��T�ƶ�]b��S�It�_�ӗ�?��n�i_=��i��rΘ� _�ʈ0���׃�$�CC�
=M�\{��Ϧ�{1��A7�sLn1�ٛ �#{��\ʛ�h��$��|�5I0�@��K���Y^�$� �EFnc���?R�i|��;J6l�+k���[�IR����=^�=j����'���˽w]%��:@�r]�b�g�!��G��ӏ�ӓJ��1�A���~��I������~c�TUp�B.)K4ʦ��R+�v���>_���
e�q��]�vI����FCd�ĉ���kW�o�V�H#i�QoD�jV� ���ʂ���F��
�Q� �H$|1<��	�CY�L�`�Ǎǹ����!m��>��ȱb|ȁ���+0>6�>�U���
���0Ś�E����C]�s��k���8�C�&6��(w�|�/|?��{���.�K)x���k����5y %d>��k�~{�x�yt5ʨ�2`F��󏣡b;���WʤqI0�BW�����O?D3�~l&��
`���`3��$��b�[��8c��W]�9�?E�1������`A�I�X��a��-O�<��H0���Y��U�I%��tX�!(U}*l^lT�)!F�$�g�|�p	řZc���RCs����E\Mg�v��5�d^��+[�. ���"�,��:���dl������\tb.�&q��gm���1C� �6j�Ag`bcJN|��ڙ=k{��M��vT޳���v����K�fo��鶩�f�]��<�L�>�[��۲�թ����1�n?gΥE�Z�m?�&
��y�� ;zͩ@�3�ھ9�iN��KMX}u�wqa�Kxdtè��-<8���v��E.a�xQޘu�(5���Y��$����T,#l���]@���t3�НW�xt.yEe��H߅���3����� M�LT�z�����U�k*Z�����mA �P-�TVԛ��q�d�O� �\4*b��]4ύRK 傊Bt*t-F�Q��+/1�AC���?J'؇/���*R��Rn���L9d��
���A���:�6�8�H����	A�����9�4
݉��X�J�^q����z4^���w��D�1"_��S�dؗV�#Z$�I1����]5��hJ\�/y0�RDa�Z/���{��d�����\�=�Z(�h�qq{\�y���!�;�Ȍ3�˹�_�l=�8@��֜}r�ġ2?�6��� ²5�כcY�Hà[(�P�+�ĕr��<1@F�7GǠ����O�l���
��(͕S!��~L�PY+������
��Q�yk�1��ѽk�~m�l� L������Gi���v?��o=4f��j����V�WȮgb:��-�G�b-0Fv�=(�⡕G�U��޳�8��P���i�x���_����/�<���]'�g�Y�-�R��r�UdZ��Ͽl3�)�W7��Q<�b	�oeq�C9|�j��ۓ�$�(	���I�'Y�a�d�v�A/1�]��-�E<�ʰj�#�(ƚϾ��̙}�����_~�����y�h���G�s����(���'1"Vf^�7ٲ?��C0ah}¼M|Y-�`D�'V"x���Q�_Agf#~{�F�q'�(��(�ee�8������0���>\�;�<��@��`�KN���6Q��ԞFn�`�;��z�y�o�ƨ�g�@J��xW��՝�mb~�����(��;*4*�PFL���ח-f�J�{�rڧ�ǒt�mG}ƭ;e�o���Ǿ���4��x��(@m�X�[@��ܘ1g \<8�g8c�"]�tP�g���,Y��R�����E��:GZ������pL����*1T�BGu�Aqr,�n\J�Q�.һ�����߫��/׷�{�&�7 � ŀ���]%LMyI6�"y��c����&���"X�H�l�%�ٴ)��΄�Ì�tCRJ�b��S����b5�.��'w&>���܅���{�+4���Ә������6��d9�kj�S�5�W����p�x���������;*�'y;�r����.ķؠ��,;@r.�l��33�~g�;#��Q���d�p�A�T�f�������:�>Y S��N�N��v ���9�η�����d��d��d �:�J�:Y �b��c��0�Z#.�~��KnF?9sdo���ץ�V��˄�d��ć�T\�g��B9>��It3d��ѹW���'z�8�؁�_�8Jھ\U�*��v�>�	 ؋�j��t����bJOJJ�� ͭ*�֖rt/�d�^ ��e3��cH45���BV�ah�0��x.�m� 'Q��D�4��bmL�ZF�X-"�E?��ߪs�e驓���T��VP��Od�aq��D�ƍHݧg?4>���$��HF���ч�Co�Db����=�> � F�WO��4��� ��� Vo�e��3�A���K����XGa��Z���E���l�bqS7q�{������,Ȕ��] ��!0|-�J�OV�ay���ē�cecmqW��
��˱�X�c��/��/���'9��nS>PC���L�V� :*���E#cwZ�X��w��	�Fצ%3�1�?�Q�kз��la���R�������!g��tl\���6�Ov}���1d6�k2a�p-E�J��s��]fv�t���m�5�ī�Pn��N�����`�p����S&N69���]�m�U5b�  Z�E����Ŀ�����-}��,N�M4To��l�HW�N�9�0/w=��_���dЊx*��w�R8�>�k)�m�a�*Ä�T��|���0�ه�8Y��,Y�0��!���M�i������������}�3��.���3��W?��!U�3�(���׳x��UE��;,X ���t/���kr�dJ�m��YD�����n���!�c���\�&�"��)U�f�0��|p\Հ��G��7�D�q���9m�����-��\!�警���F}V�>��ԉ�i�n�}%���f.���SRRh��#��~�{����w�xH,�Q�w��v�Nq˭7�'�?�Z����ڥ��d�GY�5 �W��B#��7Ưj�@y8��q�t�и(�7��س���`.�`���Wq�k)m{�Ì�K$] ���m=�q����+0�ހ�y��4�՚�2�2��e,�~��,���caP��0�x�yTI
	�����0�t��3��ȹ�2G���*�.T�쵌2x ����Z�v�kg:��4�̅*�6��dq=��v?�W�"q���b0j�xEzS2UIG��=d�c$��n}6*�#h�0���Q��(k3��(�di�l�����:Y�Dk"��-�#�x��`�T �1�8��
��Y3��\��}R f1u�y������,������Tl���ʎ�3�(:�����q������:���t��?>����F�#���v�c�o��A��Ϋ�۶m1a����rd[s�[TddKM�ζ~�^J��K��h|�Jd��30g�K��K��2���hX�W�`��A]H5�{S�R����J��*�F?��Nɽ� 78is��3XǏm&ί>�Z����� E����ώvOU�2S;,�������A�Iǔ[�fLt33@��T�4���Ȩ�CK� f�)=�z�ل]<	�t���a|j`<`��(V |^�p`�S� b�I�J&�6
�V���\�=b,-��l2)��# L_-O�\�]�Յ�r�H�ҫ�-Қhi������ͣ�#��L����.�Rh�P���j&g++��5�Es*˰��νfm�7e6^ό�|�|�{)ѿ��S�	���)1Dc� H�: �F���s�aĿ�O����&!6.e z���k�6eY��Uen|�jU�V�_�|�Q��_:��x<N�X�u��U�����i�4��2�na�� ���zu�������[3
ۈ^QPe�;u����u
��N˔��۷{⁴��Y� `�����%�o ĵr.6�2mt@�|+�h
F��(� F� ��`�Z 
�0wC)�7b����� �o<�,��V:�)�|��rY@V~A!�V#��/a&b�`þV�(��,*���C��3��В�i�aX�H��mL-��lM�z�fJF�U5��w�Т��ĳgɔI�\���\�� ���v݇z������#c�aq�����+@��By,=-M1C���ߙ7�L�w<�u�.�]��@�r�پ=t4�դ����Ŕ�=Y�ԀDtQ��Q.��
��`2�����qxWj)��=M��'ڤ*΅+�٫�""��*4��h�Ԗ��v*��z�<������U���.]�X�hb�୛\8k��U���c�����BG�E�*�0�U�����:��i3�2��b�K���i���eIL>\�V0c-�ܴG���O��YE2@#~^��T��` bR��#����5����(wg!��l�[��8I����i�b���]"��Ⴠ�2��u��j��2J�Mh�#�1bSC��.R"����#��"��7�v��2��Wl:����.��`�T��u�cM��2a�5'#W�Z@sP�E0ej�[@3�A�t~t�3F7k�a�Y�i�N����Լ�fF��1�ζ������:�
��Z݊�:g�J�\��;xp����3�d�;в���og��@���������,ٷ�}3�ۺ?��ʩ��t忓�4��Y�J�V��ߜ+��4�]�''d.�q�����΄��@XCMeE�q�]s�S
�b0C� +���lݰn7�� &eP�Ͱ-�nL\~.�7�1-ѝp{�n�H�T�?w��&wc��qi��Ώ����Y��c;�&~�l$�J8��"J%h"��?���5b�� �O��v1F`�ZRS��w��:��gfɥsǙ�EDX��!V�i,����%:����b���[8R])�)#֋����U�:�y�fU`�4�l(�Z&��#F�
����R�
Ahܹ{/�������m��ؼ%B���Q��P�z�;����WM��VVkc�i�@��/��'�V9n߬��&L�+̓1��
�b;�g=t�c�j�t�/W�<O��c�|�x%��]�>��q�ٓ� ���AJe���&�gQB`�
�qjt�P>"���0=�Ɂ�L~ЈMP�n�~���(�5\�a����t�S��ܚ�K�L�U�4#���>EGr��D�q���R����R����n��`�T�����tQ��_7��)-��ˎ}���GZ��� :����5)�c;1\���_})w̻H<����:a��Y~�n��ĶT���V�w@�v���$�1�Yla>a� �b QM#O���,8�cg�ƮC-��FhC?@�%<?o�wUz�m���S4h���T��LC��Zk	�)���g��}��w�L�Dgr?��%Fn��<��B��V��]{������&AD����r�_3M��W��(�ǝ?��:�&���� ��@(.@�QZ��)���h���1r�<���d�ɺj����[�����3�� Y�q��}A�������B��/2� Z��������ͩ�E ���*Ɵ:E�z�-s���f)����q�kן7�?��b�
c>�d>ςR�Z���'�c9�t�mmxp��3��.ؒdcEɑF�*:��Sf�I��EE~9�|������F�t��tQFw�B�9R�]A���a�{=Ѫ�r�)Qv#����G`��P���=�� y����³'Ȯ5����#�m����].�~�&e�2i��W�Ƚ[
�u�����8�L}6cv��}��{��*%n-Yw�W6A���� ��0��Tj�JR[ƙ���`I�3�grw��,�<s���l)��I.�Ru�ù�Vв2�:V�bHSNL��,����V	ʹ�g7�t�{pf���s��4�/e-�s쬊�-gm�}"�H(��s4)8�,@i�]�paׄ��,����/ ��|�>ۯ�~��[?�:w���x^m�οS��c��y�+�8����O3�8
'���&�N��t��Θ:����	���_.Gz�Ի���:�7�w����0H�=H�|�=y���d����8�Jf5:���J0��[�tʌGc��`�.���`ҩ,H#�-Դ��ge�u�^��N�� t��[n��bM�F˽vZ�`��k�7��>�V���*-Ṕ:���(� ��(K����$��b�50D9���C�*[�.w���D �p�}X���dSBX���~?]�|��� ����>n�Ei�K&��k��ߝ*�R���,����R��tz�VN�#�9�y�B��Wj���A�=3�1͔.TT�#��*�xSQ�rG�����1�Z(�p�e�/꼍?��V>ã�H�-�$��X���Jz�F��i�dT�D|�T�(gO�.CG&�&_31�?��{?&C��}L��3r�D�(�6�".B���V� ���b�T�e�+e���.e���������`��5x�M�u6��" ����ޔ$��W��L�7�3ݐ:x;έ��Qz�iiTs����y�2vؚСe�����9��z��nuR0���GM+��T�����|� ������g�֣�^ �#L�ar�9�������B&]�$��;�;�l9B�hڤ��¬2�5F�r���K
����_�߷�	8J���\�J����ߢ�*�{�O6�I����~�r&�V���޽��sG�]Z�W�NPM}�tO�'o�L2q�_��-S'��j���VH3�_��=��Gj���S�-K�|�������	���^ӧ��M��G^=�5���r�5��-?;��"���U�h@���Xn�3�CV�!_P뙄���"��NJ���GL��?-��T N	���� �,!��O#Ђ�옅�簼�R����T����s�sf��MNF�.�4���?`8��&B�c;E�X�Zr8o��>�r׶�g�m��Z�eˈa�d�����#C���/�]vn;��� �I��\+��9G�zw�����.����f4�,LJ�������f_:�]a�jj�a�x�9͊�`�sЄ��x3����o���=��n�2fD���3����S{ig��7݄ip��U�Ǫc[>|�������zA@��T;��Y�>~P%œ���P�ea�Ђyн�����N�]�!Q4	�����B2��]��nf/��0��ئ^�ތ��\i��.x�j7&��12�?:oN�gf�1�1q��8K�����;�pff�Y/k��ޯ���uv`h�L;x����si�>�:� �O���J�jɢƻ������'�����B{�8�����0Cq;����T���S��`�O����=
��ʨ}��Ƕ/����ǁ��E��U;����֜c?��=o>��/��٢���3���S����Z]JKҽ��j�5lD`=.���ގ�L�r�̳ě�G8���Nj�\�9v���7zQ^p�'1!A��\)OK����K�c�[Rwc����WƑ� �jz�~�2���LI���NP�8�3��Z8������j��#ƨ���,@a��R�j8yjG���2��L�J���)���x�<�tP�Sj�05J��8b���E��Ȧ]����j���/)��Nc+�����h�&�d�22������>t>=e���7���J."����̔�4d\)~@��aT���L��V��
`�d�ra��P�i!��|�	�в� T�;�M�ҥ�G:�(-Ǝ� ����0ܰ[��<V�ʶщ.���q	3��n �V�:!Nݗ��A���zS>n	�z��Bcw�C����ʹ��@M���7�~J;���P'�'�0ZO��n����׉�Ue9s� _��Q͗Qf�x��^@}��{ڵb�*�5�V*�W � M��G�
`����5�0�Y`rmcb6f�z�=`� r�����ad�5k&F����~����L�K�|�d��VK-��`1B`��)M�'��?Ĝ���*a"K)7�^�'%˕7݌�)NF���h�B��rӬ����7ޔ3/8Wn��,ٽ�7 ��,X�Ef�!��H�p���K��W�v�Y���wN�(���QT�#7�O��{���m�� ���Z�;��>�	�P���] %�`�����q�d�����o��4�y%�����';e/v2�5�	q.�x�K�q���B�̫����ݤ[e�����t���ut�E�U��LJ��Q����S.&n�{�aYE��ݴU6n_!�Χ�w��⑦c�+�K��d:Pÿ��"2
�CPM�س����N�u��ش���?ǳ�g�|��r�-W��X�ʔ�uT�J���˛��-��9�g�U���M����5&H�Q� ���N�L�y">�����M;�g�nr���r8��x$���E���6�x�9g���gʷ��H������Ӑ�ɧ�e���x@u#�\3��,T��VJѩhY�|������Cꃇ,[�U�Ѕ�c@��4����X%ūY@��W܊fՕ���Cu~s,T�0�n��Q:�F�ߠ���b|ѭe��;��:��	c��"2P���}��䘉�r�^�3���Zd',]�i�QS?��b�!��s���I7��aۭ��yG�u�l�3��J�'~�ٍW;Z��3v@w2��y�vPc}^G��~f}FG���hg����sb�u,g|���,�O_ߑ����r��3}��=���)�X<k;.�g���c9q-0�S�`ȱ����~�Q��h����2��2���[u<��S���{|��y�E��l��2�h�Ø�u�0ӏ����~�e�ȶ=}�����e�ƽ2g�:}z�b��8�Њ^A�ŗ�X1��Q�Dܘ �(�4�_
@��s��b�\���І4ג{Gi��4��)�hb�q0��oҖr��aX�Ĺj����jYe�b*����=��B`KY�_W��֓/_�>��jht5�����j�ڑc�t�e�Jv�yW���t��e���Řf��qS��/%�e���Drv� �$����2�__��ʋe���/9N���鏭�'>V�|�_+���ʥ�ϔ &�R�������+>ǅvh!��(�6-�}�`��"0��Ñ!��5ӓi�ꌴ�K0C�� ڵ��.;o�� L3`�eX7�_�����s�ҬF)0Va;���(� .!�^m��$
����7$;2��g�e�f&O�P�f�cP�ÊV�Q��2��*�77�,��hT�J�&l��8A��i�묀N��*��Q�(���´���eV0j?�57�1 ��cL���v����� S�<��T����Dci��U��lK5vh�nq�^dfoL�
�Q=ux&%&fo�0�/;�^.�)�� ]��`?�`93Js�#�n'�3Ь���zf�z� �h���ى��S�A��W��&g�9�LT[7o2���]�e
B�a.$k쐶�8r2/�\&�\X�P�׮x]���7��vV�V �a����Y�a��壏��/��gT��/�"H�/��~��Ŝy׾�RY�IFi_9g|Wy��'%����]�q�?��p���Do��_,��	���V�"������S��3��\8�$���0���8���=v@&�y �!�Fv���e�/��k?��Xf��\9o�̻q�I;@9��b2M5����NelgB`�T&�z�FJ}e,暙�gκ�EVB�|�#�5E��������{� @�*��r�o�d̨	r�X�)������2Ln�l��d�f�8�l4fz��Ө�e�VY�3�4ͬ�?\>%�%�7�p�3&��MR�Q,?�p�׮�*���.�#j/�㼁&Ol;�x�+yF۸4��Z�g��pŋ��g�����Y��;\,����yr��9 �/���ޕISF��wJce���އ�\QD���|7�I#��6|iP*�}pm ��-WW=����5�q\F'*�%�f����v�� <�玟U���e������)�7�;&�������9fLh�7 �U'f����V�p�����}��Bv�b�RS�t|��]i�:��?O��˙=��U����9��)8�(gPc\�g8�"$�j�-�d"�e�:j�^k?w}���t%Ԏ��b䜯˩��Ɏ��9
��\�	���S���N�9����h��E�����_��w�[�L�k&������kxl�k~z�|��"bL*e𰑲p�b	Eo����2Z�VLG5lW��{��� � .�@�QK'PO~(!�bJؚ�dU"Tv�7���Jt(��y�)"�T�d���'/���8N�q�	�ߥ��w��x�0��Ł��R�1E�� �*�-@�"O<�w�����«o�]��f2S3��C�J��\s�l��3R~�YDSA9 �� V�h@�����S>�����{e�91��$��@%�� &<w�r&�ܹ�_2�SzU����d)iq0(� ���.e���1����֫�Z 7<�(u��y L](�+�Bf0l̜ig�p|*i��#:$�T�R��2�n~�|)�|�h��ر}`/������:X؛����~2�`�Q8�kT��}��p�n�C3C%f�� M�j��a� !�$0#�wܪ�L9@W;(�q��ߗ��f��P�U~��� ���k��ӳa~�=���S6������\u��Z�@��� &}p5�ޝ�+ t庠nH���6K����S�E�N5HSYG�{S���2ʿ|�AX}�<(���������߻�&o��w����\�u,H�ӆ��h�:�1�y�^d�cՎay��?�N?M�pŢ��gKǚ&�`|��x�	����F7ު���2A��y�I���j�{�����Ha�;f���k�K�	���}����K>_yiң7Y��7��{��yse������^C|ݙ.�lk�dޜ�Rʤ�~'�����>ۻG����0���! 3��EU+�w��DHI���<}�嘃zr��������J^�1�R90!r�%�趄u�N�(W9J,Rk��r��d�Uҏ�P?�{�G|�z�3�~6-;��e��]t�r�ӏ�ɶ�(ߡ颼v��s|����2���X��޿s��c��ЋF�ĤH�P)�t�7�I�&JVf�Y��!�8϶`��kc�π�ñ�HĐ�1))�8B��D-^�Ҥ���G�-[nƌ7�D5��>h3��Y�6����ξ����	0Y@������F�F'�F���a�eI'����~�5s�ڶ�-w߁]P��0�x���/�W_y�U�$�����nY�p�L�?0o��8�R�W"�)��xu�Ze��ذ�X- x��X��FX'q g<���]�B�`�6�7$�|�2�!����`�(�O0Ȧ1�
N�Zu-�Ŀ5������R��l�X��}�SI���i�c/�Y݅�� {��T�}~����[�f��d��g@h���������OX��kg��w��ѹ��ͮ�sa�<v૟a��^�te�[eӎΉ�9lefk�־�g/	;��>���o}�i��
���;�(����1;v���S���E�	��vk����}��c��e�/kd+-��y�l=�} +7�+�,����i- �L�����U�	0 x���mbB�C��x>�RW +�8�W���5��R��F֠��d�+C�������=駾Q�j�h���e���5��b�c��
��b��0���q,�Y6����<�Ϊ5�` jd����/9�.�%���:����{��/%�U�fʍ���2z���XuS�I��'����LD�p�������d����ٛg��/~-��1�cf�K��e�cK�����Y��7>�_ec4�E/�;��>0'>�tR���PI񢰆���UX`\$�����'���#����R�h�wGW���������t�+���F�B�Y��dr����t��t>��\M�tօ@a��1p,BZ̕r`9��cvܻ���ǰ�&r��e�϶��A;UO��6���);k���jjð��SnˀX3E�D��������,9X.w��~n\k�<�t5ԬF�jT� �F����4��:j�(�$JԘ��)$R	ƥ�3��g$F��L�tj�^nn����kғ&�$J\9�za(�au��q']yx�Z�F6o�8��!0�x���屧ߐ/8K.�����{��k��� �>�xO, �lBS9t�TɕD��xh%�r� ��l*�.aF�9�+�v���_xϬ��(���6Q�����4��+玔��d�2~%ʂb���8���ҟ���P�
��6ʶM;��;������Y �~�9�{����o��*���	?u ���bp[(��E��y���*_)}�|�ŇaS
��d!� }�X^|���[`��d��fq��O���qQ$D�eLi +�{������w>B�g�,7��@钋/��&J�,p�[?�4�\|�>��+Y�z%��M����e�%��A�rZ�6Mp�6n> ���,&�/���W]M<�$�f�O�ُe��%[��J�<~"l��z�����R�|�_iF���k#@K�u���[}X����X�I��Y�Nv���������3�s/>#�9��n�v��?�����}%�F���f��	g˞u�'Y�0>�5m������`Q��#��dm41Nd}�ИĘ�s�v	��#�s��ť%�haʀ���z�������
�+$󵎱�W����VEt2���Z!�z�X�9�:� ��w��`��`�b"����>�;O��	��ݮ�:�:K�<�[@����>�'�����j_;�?;`�ZݲU�s֙ف�.�����y{��Z̙=FIg�s����]G@��>�g���lhG��t��(^���j��o����L�f
<ًOT�N������l�޽z{��㛖����8��A0[�?o������7�M�%�C�+]8�!L�]�{!V���;D�^]����ĪNKH���{x�@�Il�G��z|�lՖitѬT�C�Kg�N�u��*���@�Ӓ�j� J�F��5μ(�OM3��=����,��Njd%�@��ɸd5`��K�(4<�L�x��%�v�����}�+����W?����"A0K���k2~roL"�aN7�tr5���>C�9���3J��C�o~� �N�+s��_���⋠6�c�����<C"��gr��Q�,xFS���sϽ K]��B��/��l:��̝����%�
�ך���by��7еdHx�`âC4���i	CT����j��W#��y+�@�Ek� -4<4�w3`��� @�+�j�Ks�o�{v
����1�Qv�P)df�W3_���o�t)�=�nP��>D�����Qu)����Ź$3�{��z��),SK��#cb�L�W�L���:����^�$H����7p�0�䊖��;��F���e6 ����� ��n:I^��K�9肨���տ�f�0��6�}����f��*��Hy���r������d�����%��W?o�mG2�`!�<c��a!�ς�I�kV�w߮[�8;Mb`����Z��qRN�ѻo�AJn ,:L^y�i�T8�Q7y����C�up�|���2ih��
L����{��^"ǡ�p1�{!�?
��@�����}%�p|�(MƅN��<�,��y�JpeJ��{�LG6*�>Y��:!�y+��-#Gt��/�Hi+ER����^#���wٷw�<�ģ��x�Mʝ�^#�9[�,^$�=�O�h���d��!*��"�7��4���Ì�!G��P�<<���;{\�f�3�To�8V��:��0�U��̴<އ��� <r�P������Ir�=7�暮��ϻ�R����kϕ����X�	���m��� phM)��TQ��X�@	ϔS��ѯ��J���h�|g��5a�`y��oˮݻ)�F��F�4a�7c�u��/]�X�'#�����E����}���$�F W�����"������]�w�l:��F$O���ps�{�H��1T E�<]���a�v�jeV�j|���g�����)=*�]��EF҄Ʊ����6�h��Fu�,C�q��iI[Ӓ:��['u{W�5���?�|��r�_�����D��>��ZY��\&��׾[}�3��Ѷ�tr��I����sf�7;�Cg�hg��ߝl_�se?�99 :������&���Y�~��;:�����.r�����;����� 7�911N�$��Htz+rЪЉ�hX���N��J����T1��@�WQ���-�(��`mn� 2�$���@GF�����$��,���v)U!9��_P4��v_X$-������R���UDl�#�nei�p\�`uɆ"RO�*"%5�Q�D0�`jy���r�����k�f��7�t>e�j�ճ�$��mh��NH�)�?q��3�6��K�V��祘^��.� �:΅?��ūȥ��Ζ�0a�ƍ�|yIvf�a�h�?�Bp��L:hz�m`�|� |5��A�[=� [m�89JP[�$F�ɴ��9���O�����{RX�q&l��\�����[�Ls1�����x��W_���b�D'�!�m�^{S�>p��$5|pj����Y��6�]U�B�����r��B��� 0�#�ū��ff1G�_VT�~��j�����-�~����������!�ӡ���2����0��MU_fe���� p�
sq�{O�,T��k�f��8㺿jg�>R�u!P��G���J��yp�b.3�
��m�;V,���S�U�\m:��(!��8ঝf0���p4`݇�R�w��ۇ�~t~Ut�����'�P,]�?x�ж.� 1݇��K�ȏ���r��0v/ٞZ(�/�d<����`R����|����*�]���äKT �*E��^-#��Ax�}��/�`���7���'�9i��d1����˾��b}I���2����O>�Z#���7�r�h��>�)�8�4+D�̯��\b��+"ݢ��u�2�EM�>0�-.% >r]�!p�&���$ �����O�l��~�[bOY���؛���z\�C��G2��.��ͅl&�g$e���� ��2l�0�L����Xbxm��0¿����3�ă�ee��T�4U��`�Ș�e���ь�
,9��W�[?���fL3a�����\v���.bql�����ї��g���M���S!�Lu��x� ��+`�T'�KyӋ�����1ÓEA b9���=؇:�o��v6 �m4��\�n܇~��EJvN�̝y.��ٻc�4a��^+�Ƥ0�專.m	,��$��_�̜�� �[$��sQʂ,�.^��x���y���H�n}h����*��t1����__���3���``�W��_� c�,��+���VFT�f&5-�2�4�[I�>�;��0ݑ�ߚ��@M�w*a�}"�������pd7������;8�*����!������9�u<v���Z�k���6������q��-�\g�e��]{����̾]�z��˾o')w��S�1������%��(�5f�s��ۂHan�7�\L�/�r9��kF��ں��]{�z�VfMr��7�~�~ƴy�ŭ�|1L\��̝.500)R�ƥ�M�4�C)l۾c��	wM�=�J>Z�<J|�O�e��l�:V��D��0�y��B�O	���F�kh`E�ˀ^T�*U�z�H�!�+/7� ���N;uर�Mb���lG0�G�A'����v޹r��Ɏ-+�Ï�ԝ%�{�l�,���R� ��n��O��9gv��x�gk@oS'��I m-����c�>�\q�IL�T)�̓/�Z"G�������	6L�.�/z�Uu�+`s+��0��]�+UP � � ��[&�O�)���-�vl����ʻ_!�.,�N�=��)7N�1�.1w	'Im&��τ[��R =������ ��&V��>����xP���W�D��2�+Z"-/��O� �f�f��$��������c��o��@�����}������!r��U���	߆R+Bfw��j���g�ո�T�CQϗ�Zq7&,=w��WN��2�p��f�e���t�7V(�`���te�{Q ��0�X�뱩v��Ymq�p�"�8Z@s#�J&^M.�.R�Ǎ�s��r@ǒU�����,pU'��13�W;��E�	kr3$v�s�h�`b�>mڲ=�v"�)Y �$��	c�Zw��/�4��u��o|��5����2W����.��j@�2<�A�2�IrƘ$��7��]��{�[w����1I���j�ҟ�ic�K��ٳ����̹���bnN6פV��.�j
��ޗi�'��^JV>�|�2��j�4dGe*)8�<�d��E᳗~���S*]����Y��f��[h�IK?��q�<W|�ʼC;`@�y���\u)qܿ��X#;wm�����'F�ت ���ɍ��t�lۺEn��0j��0,��Y[C��`8��f:Qz/��3�s��n�fi��2���3d���<�n����ԀOW":��A��Xܸ��3H��+O>�����2eltj��e��^r����_y��X�2 O�a��(�ӝ��=U�?Z0��^0��t;��ua��� 7Wb,�%������[� �CW9�ʟ�>GXPn�W^(�{n�N��ı�e��4�����`�i~�gFwcǑ%>M�Dƍ����̺�Z�ox(j$��Z�2��a�ݹgՌY;u��P]H4��Yp{�A��%�,4* �m*�u�27� 6�Bׄј�覚a�AML�a�t}�clo�B�"�:�޹��KcM�΀�#ps�I��:bҜ��3{d��u�ov��PZ����u\�%B{g��HY�g��~���0-�v2�e��������ϴ�}*Pt��utn��#��6m�� ��{�h��̓�� ����2���p�N?���>:	RA�E:%�h�+Z��#�u�C(��O�n#Zw�տ
Y�11�����)S���$My��6MR)��BS�yeE��1�2yԗ�bH-���\���W��45��jd��I_cM:c�ZZ��PQ�x��Sb(n��I���d�te�s �4[�{���*�ƻ������Vw�}���:L�1T��1���e -�����,T��󚕰Y��|���!���k�E�H�a㥞��	�h�$}�巒Jya0ViYy��0�=T�`����<�p(�V�eJz�R���p�V�qy��R��M3\��9F��.u�X0�._��M������I�e�7+�������^ 1F�v�xRU�Q�$;w����϶L#n?w�Yt�M�<�����$�����d���&�p�)1z1� ژ�[�iƐT�r t�Aa�LQ��`(o���z��f��� ��s�烞D�"�H��E-�-<�1�*�ǉ�)�+h��J2����x���De�u� �6Q�P;lP*k�� ,(�l\��q�Ё��n�sK��tͳ@��9�F��0�U����] ��L�^m�ѫX�P�6�-y����2t�I
�����[X �Q���n��TV� �����r֡'�!�ї����B�s��̒�zQ���$�A����wK ]��gHva`'��G�H)�/���ƚ��j‪�^�<7���le̇�G>ݰ_��^�e��P������0n�Q�ڇop��S�|R���=g�\vɥ,4<�@L �I�{ɇ�.~4�<����>�]h���Y~�XSn�F/0"&�i�VF�}9e��Fә��z�>åqw
��d޵#�ju�j���,Y�V<V��W�|C��rSbKOI���� q���CV�8 �R4�`�� Ō���LK��É3��a�@�y��2bp< �@^n,#�s?7b��F�{��YB���a�B1c!Q#z����=�6C� lm\ ҙǳ��Br*��gɓ4�L�>C��|���a�F�!=�,V�a��>�Gg�3��/�D���A��$h���g��{\5��l�;��B����;�� ��CGe����h;�����ET����=4���{؀�Vƚ>4
r��qf�{�C`�;�#��mr��	���%�%�I[���e��z��fAmXT#i�e��H���U�j0�(#ֆ�O`�Fp��}0{0?�S��|]`�>_j�m���x�i
.��G��GM[+nXr�q��)�t���,�ŘX��d�K�:��#�NW�r�L팘3���Z?s�:Y`��{��bt� �#vNo	�����K�CK¢�m���޹�h�ۏ�jz���(u��sf��L�����������:'��[�E�m"�o�؏�h�Ϝ8k?��O�N����0�Y���UV�ZȲ1����0"`�|<['_4;0]��m{e$���i�'K�B����N�O+Q���:�ť�cL�H`����&����y52�)�h�	v��rA @(fg�����+���}蓠�xpU0^��wK��!@����R�w�=�-{��1h�/yi�a< L�{s(ב�G��WX����w��
�9�]J�s
��|YB|I*a������Z�"=a�!�M�S����@z/id�1j��!$����D�\
�5�_O�y�8	�	����Eu��ղx�@t��Q.�����Znۋ�d�'���f b��xZ�ך$�U䴉#T��D���w���9J	xɎT���r�mse��0-�Ə�}i�Ę0�>������P�"0�[Y'�\>[b��0�m��?/�\3�N�p9cT�u�(�_C���Os�I�z�ヵ}�V<�����c�Gb�,����ں��1�5V�F����c�0�d�&r�UYy���Mr�g�7*�~�I�'`z�XI���w��7�R�.$f�N L��L"�xT�$9��8���	KƈA~]��}����xR��%�%S�J��d�IˇŬ�L�1oH'��F��4>ᗡ�zJ-4\s�4P��u���n�E�Y��K�/�6�QD����W&�w��Q�2c�p��r�1�*�cы�(jbb+�ԤF����6ו�� W��Y@�ɒCϠC1�d�f+n��S�ļ�r] @����63|)s��Y35bp�iM`t�O�>X�-�������R�H���ΕM�����\ݤ��?�L��=S.:�|�Q&�eS�����r��g��<á_T<��kt�ˣ��)Ӧ]`����_�H�=d�Yӥ"�C��p�l?����2+����0 �I�x�my��y�h���q/�=z?^~����.iwæ��3�~�n>S[�ŋ~�����7r������d��+ijB_U���),o���<)�(̔GW���f�Au�[7I ��p"��in��ù��"�{�0"�PD�� �4����X~�����W ̌�\D�j6�.�]�e,�@2qQ�a�`|;wI 퀱�1l�`����⿲����b�CYӕ�
�q��x�e^F���	`!��j�Bv��3zS�����L��$A~��RJ=j��3�ƚ�(�VJ����p�9����?7*?� �y?�J�2m� X�F�>d�<�������STC����`�!�$�����
F�0���0bn*O�CЏp��;����N�F*o@X,����習;�E��3L�Ra�<5=n��V�lT=�@NV6�3#M���O�rX��_̙��)�&����ϲ�c�޴�R�v퓶Y��~����۷mgϜ�i/OZ�ľ=;���+��Y@�G���Y6��ف��J�� ��o�8��k��̝��03��v��c�����[�Z���cqx՜��_f��գgCb\����ɢ/~�q���y^ �Ȏیik!-��0~A�|�I�x���Ё=����r\�������ҌB7�`e<�*J�LD��U$���¤�� Y���
�����)it���dЋI5�{����ܸ1ѢD�jkA���>9y5ҒW"�
�TsC�Q�+�eMv+@a��u���_d֔ar"�b����ᒽ����!�N�v��N���%R�[�\z�U��%k�6!���`?�P���C���!F���>5�q��zg�uC3�7q=�7 L!�:�+(���1��a��MЌx2�4�����{zU�J,��[ �D����|�:4�l��)@7��[G'Z?&����0����:뜙rÕ���4��~N�����x�A7� �;c�q�Ğ�U�	#�M�I�L�'�FP6�&� ����b��&?��t6j��ˈ���
�Q��-� a��`T��ʱ�l�;$�اh��zX�@o��6$q�l�SLk>���ғ2ڥ�%��~��{(1))ҏ�� �G)Z�}��g��e�Ε1|n"~J`�&�~���L�ŒMr�źBc��k2�F��X�^{"�F\��;�D��/a0�C|�wt	�~�2�*��,���jd�@��R<����n��Y�!pь����'��@�RK��:�UR�9�] . ����r��t�`_�����O��U�x�FuhՎÍ�i+h��Rz�Qw�mm�-X˲�{�a)�@ ��CG��:&7��a6�;�[�γ��s����n�1���ݷ^�����&O�7_z��<x�m�`�Z,#��4�RBa��{����s����Wː���^\�Ϟx��5}��{�m��턭�c�J�6�'��e�}�����W�+���V-��O�$��_���Jo4M6�(��/W͛-/����x�l�$�6������=� e��q��Z��&?ӓc����sΞ#�]�e� :���Ի?���ˉ#�jﮝ0����Y�ٷ ^��8�M8{�<������o˙gM� �j?��фo_Ӎ�����K��9��,4ː�A��c]M�h�r�h��X��A��I�R{��V��No5hid(��:'��͗�`Wk=�ǅe�����·��X.��?O�n�<��u0_�r�Ug���>���ț4^$ �o���� RK�l*�_jȬ�yO�tk��ӛ�Q���.0���նJPT����&�8_��]U<�s��+��0��P�0��b۪�lPƪ�M��ٲ�g��y��d�j���wX��m��θt����;�f!Οk��nP���9�~:b�L�ݟ̀�cr@TXߛY�������'�_�8�m���~L��`������w2��ئC���Y�������osN:q�L�����s<�ky�Z����כ���%啾�SR�£릌��ӿKw!Vf����,�u�\�ߌe��h?4g,��>�\$�s���d`B�TI���AWU6��y9)r��!V�Q&����� ڍУ��T�� J>�����̣Bϙ3�J?\���e��l'].8�B����s�I1:�&�b>�ߴ���<�"�@�bLi�N�l�A/ ���zH<��I�zJ4 '��l��&� �b.,]�E�hu��WH4v
Ԏ=(g��H<L�l��͓����N�|��Dh�a�J*jd�ν�ڹ]����Y��-7Z�B��r���U>!�7���ѕ�$�q�14L��KWɐns��)�r���{��x�V�H�V��ɔ���
��"�3��� �3{e�@Y�b��j�C�vݶ=��G_�(1�����l(�64U����6��u�R�1�q�C<S��wY��j�@����dĀ�8���Æ�:x��߷�0 �u����k�I9�Ld�Q6�{`X����o6ˤ3ϒ��s�ĝ�EjR�j��C)�2�݃F�nݻ3M`�AH9�8�_2���Ѳg�ny�ەD�L0]��G�����:�S�� %���.��R��B5a10�u0$5�ӺF�#��J%���=.F��Eȝ��-�W��P�\<��~8�6S�r��ڨ�xjl��SWB��V�6D#�<��-�ˣ#�I�gL��;�0^���y31��S�n�ك�.5(�>DK=5�kUx��jyM�h��C2��:��s�+2��)R~X�"Q��rם�IvJ�<��kҿ[�
�V�I2��:D�4bl\�QΦy#
vҟ���+�ȇ�
�i�L�Pʻ�/�)_x�����@3�ڭ�TW,�^x�~=�V��s�y�2q�66<F��3YRrk�xf�<���e�B"�\����xX.�`^U�,܊��_��Z�:��L�a����s�M��[_�o�[x���ɷ,�A�XB��,7v$�DJĀ�6�ق_h@���}X��?�lI��b���k4?�A|% �g|�Ơ?)=)Q�ó�LYYLi Qx��p��Fn`�x��1��{�ٳ�}�ˌ��\w+^�m�����y���I5R�*
���hr�.Vip㢩�Q��]i8��0vtU�<�{����};��DȅR�	M��i>�֫�\p��r���M�M73/��Ԁ=f���̟��"?x)�z5Wv��^}%���q�>K�#aD=��I���Ri	�0����Jno�1m�j�LiѴ���F�6e>U���ӹBm���ڡ������"���5���E���쓵5w�٦�M��{,q�}���m��,0c�m/�9�N�m�k���n�n������ ������:@�r�u���Dg����Ιu=,V���3p�o�����}?��ig�K����|n�c�����N���H�ĭ�C}�,FV�7j;u��-�@�/�0���:�E|?������h�D���7n�
kR��8JgI3�q�x�`�ZІD�@JP��(���z1�'�ջ�0ږke��k]�Y���JOŝ>�.!�ѓ��]��*�+}$��NV�Ig�Zy������G�A�ul��Pr�F!V΍jTeR2,]��Ey�+xw&���Ќ��j��#�xÍsdl�hYC��7�~){���^��z��*��h��J����ߙ ܮ�)�P7h��N=.��a�a=�@��/P��%�X(���Ǟ��`�Su���
�N ��몗����ej�3��&�`eF��N'�#Z#\N�̔c �xJ�R�@sBm�L���*+[>|g�\p�,�J`q-�̳�E��/�f�b�,�S�dG��1�����d�����D�J�2�Up�Ҋ��
r8L�r��C�e�&���e�˻��� �Vn��%S'�F{�
����_�����* ���Tm�pc���z&�J����a�l>Z(������Ԥ�����?a��q��1�����_�a��Ph�{n�Z&��� U���t�sd�-��sO˙t�jg�;V���΢�áWT1�F�	�6
aGT�Y���Ѱ�E9���.��U��B���2��닦�Q�����B���{�epQ	���@S!<�"S-Նy����Q=���,
�]us%��}�t�`˪a��\d@�d�%��a�³�MsB3zGmv	�.��N!%�:������ń��FmtW�]�Y0��+WKe�/����������A=aV���g_��o�^>��}��{���S��A��N��z����ɻ��0b:�����0X��A@YP�����ƫ.��f�����,	g�����䫏ߔ����Er��/I\�A��[Yg��J�5�տ_�\���ﾻ�o����~�1<LW�PM��������}T��_&G2�JvF��\�Z��o���̑a�zɚ���U��0������ke؈���"$;�o��o�����%��Jd�Z���s�D�S9�:W�^�XĐ1G.�n��� �!��?�����X$Y���4�O�Y�<�H3ף��y�u�8V��O�3a�)��b-é�Y���>Z� X8z��iH�Q��`B�9O�=�0��Ŕ�[��+.�M
�=i����o���$}3%1f}�v�录�, �1|������QD�6��h�E�|�s��"̍JAb���5�Q��@�2��Swc�C2χQ��7�ǳ��VBr��O8U W`��J���|��g��f1��9�ne�SvL�zL�t;��0Wf��1���I��2�3�p��Ot쯳3Gv bW����x'۾�=hg��h�rl��:Y�e�*gF������΋��p�3qv0bV�LSG۶��#��~��ύL������YE��9�ݟ� �s:�����L9�OLן6h���,�7��_aD��"�GU���"�;q�p��B�w������j"I������ƨfB,�jY��I�ڥ6�LGvAtL��$�!m��Cw3�v����p毒�TӼ'������$�o2�J_)=�[�n[+YC�)	^�
�7I;vHz�x���Q��k�K�Ź_��t���ho\�t}u@	 �����odG��T�Կ	���%���\	�3-���d����_���dd���W���F���5�
����djB ������ �H�&7219P�)I����Z4PC���O��V6L]�M�!S�/z������h�f��������̆��=x��ݠf�0}��}hX��EG$Yyu�2f�ɣK51)A)!����F��IYX���[2P�<����06"F��m��,F�|9��i�	�MHG���Dq�e����D�$��L��v?E�2d ݁u���(�����H��ҷ��h�*�l��\��G�)�S�bi�xm�K�z�X�ė(���@�9�Hv���4�!s�|�� `b8��"ɫh�����=d�5�Ȍ)c�B��������O��IY�:��X��N6��T&?�aUe#�� 	�m�����r��L<c� �ϖ�u	2�-����d��
0�<�ä�@�د�D `C(i�ܵGr)o�A�K.j����jaA}���D��kZ�dM�#��ףQFQ��:�/^U� q(WL�&�U5z-\�z�dG��Ҧqb�yHHc�ц��.tjy��R�x�M��sW^q�$�u�Ԑ���]+)��T{ ȯ���9y�9Jm��"�����>v7�nCwU&�F���^��%?�xҨ�h��+7˹�ȡ-�$6���~V%X&��)e��]Ҟ�\�y�c��Sd̙�v8�j9�ҽ{���Gu�T���G���3����a�+�jOs�'I|�`���W���<��	�̟;N76,`�q���]���Hx��,�e-ٝ�h�r$m�6�4��&�}��8D(� ƟP�� �5����)�l?�lo@g$���q�keĐ�r�u��!�?�� 2��,��:%�Cix�[U�J�rU��`nVk�n�͂�r�/�Tj 9h/'�.��B7n��F7���E�9s�[�����I�^~�<�����C�4U�e��"c\��u��S��f��òƛ�"oL6m�"m����3�};�I�]%���@�T�#L�1a�1I�w���C;8��Ab!Z#i�i4�t�6�>]�k,�#��4�qcW�x�%5e��i⋴;Y�<;���XҚ?�Dg�����5ֿ����84��v��s��t �y�v�`�}�vA~GL��Gω�,&�����wf����g[��Y��~N- �?��?������#g���:_kO�+���~\�~��'�=�pu{���uO�������i��0a'̄OY����eV�����U~ˍ7G��A1�*��y�$��Gɞ��F���X�w�����7�~(v�a`���Z��`ܘ�|X1�2�T��)�E�WH_� 	R�@�@�K�^0�\1:oܾ���_XLl�;��1cz���u��58���F4���&�p+��C�ܦ���nʹ\c������>S�d�봼6�.�s�H~ ��Y�vIm������c?��׏��S�o�+/���s,,��ڊ��S���[ѣ�����]s"=}"$!��ND�G+%#O*��*f՛��I�FDs��b<l��R �^�7
}�g @�L@A ���ց�j$] ���O���F��X�ן���U�Y��;�cD#�5���t�zV��wT�~�R�b��1c�Q~�(�E\���8�wav��@�4�i뱃��k�O'_(,:=,.���q�����x��:���}�'�1/�XBar4�9��Ѵ&�:E�KOV��MXW�ĵ� ��K�W �X�2�0y�P.��E!XW�2&bU�j��k��/ ���9m�Ol-�,8z4�L�O��%Cp��`y���W_9}�ܵL,@����������-��͵�I_��T_L�)݂�d/��o
p���r�A�ɘ�2`�hx��D���),.8�x޿)6H��'5z�<~�Y���m���b{�]�c6����������^�P.�y5<]�����`�5]���26�	X� "GR�v�V�G�hr(d[Lx��0֝��z�E۩���$h�����r��	�VV˳�~^��.3/�#���U�������}��C��m��]eΜ��.@np�g����3�o5r�ݷˋ�>)�=�$l~y �l�U(J[���L^ZN��o� {s#8�³������8�H��䦜9A�@~���q]�^pO%��Y<�!�WMZ�+i тr�
�_�+e��A0X��2pd_I=�W�`{���R@��
d2�����օ�mIa!�����ٗޅ��&ᔺ}(��25�yDt���}D#e�f�n�'��I,/�c����Y�R�U�_��K��3o~��!.��]do�!4�^<sѦن�F@@];��U^��Xl1FiWc3��pF&�`d\���~�VU$�,�Q��l��t��$#%C.Y.qI$��$w�V3��)c��_������f���ʸ3��ZS���0;`���3A�n=,��٦y���d󜸸���7�#��XI}�T���KK�	`��Z.8�L�.���Ō?���߀5ާy��lˇ����<��C�ߤ�u� �eDL����ԉf=P;;�<�Z Śx퓵�g�5�ہ�����D��$��� �T:{���A�}?,0e?vcg�쬘�1{�eFg���̓�0g0������c�_����5�c�c�����X8{��?��lX�Z�a������2ss;г1&�8Ǐ�2sm�e�������e.�������'�^@�v��Y��wX�K�1:p�¢�_E'L�l����^n�J�N7Vzu,-��4[2݄?e/l#�K��B���1�}PT4<�ĥ�jt��tN]4i�t���n�F���/Ƀ������O��o�&�t,iWQ
+�B4"����" �t��j�6��M�>}d��q�a�Z9sP7��.���#_�χ�˱h��G+�Zz� �9�ǟ�Nj��, ����G\ ������aI��[�e�r��A8u��.����◜��\;�Ћ�f����>CK�'��}�,���Z�a�ԁ��]��y&9r���y���[a��Jf`ף��Ϊj:G~+�㯾���fҹv��&����u�&�r���u�>�:h�����/~�*�xiɫ�c1-�̙)M�*T�T��Ƶ�4߅('m�bp�Ɗ�їFDg�2(%J,������,Wd���20���9��(�t=�7� �XQ���`gI��3�-��j��o@|'�ƻv�,M�w2)�ˤ~���)�o�vB��� ʛ�d~��CB�7�v��=jI���RX�+pr�pK�[)��2!�0i� 0������+ƣh�" �S&N3%���cD�$I,�#{�<����Pm���Qא�^'}��صM�>�}�I�٩�p�C� �}�+�L�{V�@�wT�|�r�
X�a�ۭW��=e��帼��Dmټ�8��x�ߌߕ�-��({��e&<�I-o]r�e �Fپg��ھG��(�^Ù��V�$��R-�V8�¿_�q�Δo�����>~�]���䵷^��_C�x�%X�]�"�ɤ%�~�a�a�)9X��o�,�������<�]�dd�>rp�r�%&PJ�Ex��P�M<TV�8b�A�8��d���lȜ=FƏE��|R'��_�bǸBぷ[0�5���~z��>�w�X=��N�������a7�?מ褺Jdc<X������������eK$�!�Ɲ�a�9��/<,����l��6(��� ��+�|Agd=Z1,Q����ҭ�!���y���)ŕ˝7�e�a�>|?�_n����h0�POXh����ꂰ���F�P��͌�m�Ն��a�͗/���e�Z��0�hI�<��إ�/;v�0b�ںy���H2�G]e�f���#+�|����=��3���Y~y>nF�&�UاdK=6#m^�tr��VL��	>�5T�E��'&o��˨�T��:�#�ۢsHf��4&t   IDATH(�6P�e�
����~m�T_��Pvlǌ���4�3WКk���*��$h���M�γ�5AwĠ����r���y��3]v�۵��m���2��O�{vsY��ܙI�@���q���[�h�u��������;�:<gP�j`g�����-gp���cr����)��G����;�y��r�q4p^ͩ��a��|�o#n$끕ө�ÿ�B��|]��,XX�k���D<��9��L�@c` 2�v��F��Fᔏ�'pn*�6�%u˧-}MDL 5�RI&�%��'x�T�4�ހWl�O��D�]P�jn�ԩ�m���l�8D�"�ɾ�"t8���֌X���q��{71���F,a��<Jut���FeMXW�7S�nl�n�.���{?b,�%�_s%�z����L���y��n�E (�N����a�4"���j��J���AA�2������dX��	�؈пL�o)E�A�[�N�J�XeXm?��n�4�	�n�3"�±�`0c�.��V	�Q��#�N/R����,�k0���?"�F�)���l�.��9#��~�Z��G���j��d5pnh�(&vI��p�P��S��`
��v���Ij�ï
�Bi
�-Z0�V�����_#d�׶�y=<�N��� M��&�l�:��y��S=L�h���H�_<��0+���Z���R�G�P<��������E���7��T4Ly�Jh3�Ğ{��r�2�+<��+�̊��l�ߎ4I����
��0����/�<}��@0���j	��5hh@$���	In9��(���M���v��op��x 6,j/�R�ɓGKM6���z���N+��i�]A���2�o���|��K�T,����V� �̙D9�F��60�u6�m�x�W5]h��||�<t�D&O�*��K
y��qy�.~m��y9�w������ۤ0�D�|�E�T������1 rh*N�U�9�����C�xT�|�9y���G_����MW_���)����C��c��K��+���9s���_~W^��-�6� D2���vȌ�n�>ꄐ�M�h��$�<B�2�������e�����#$��J@�f�zq�46H,y���^6�>��*�(®��ȃ�!��}�lI��rђ�X8��}tT��m����H��`lU�Y���ܹ�wy��w���.���Urk1��P�
|��!�H�5����Tt�a1Ir�uXd���{o(�V.�I�' !w<|��@y���
w�ᅲz-ב�B�Y|��}����a���݌�
�k��0�Ǡ�R�b+�g:�R����B�Q~�|��/��XƐK��Jy.1J�a�4m�!�ϣ	��W�|���>ƹ��!t�.U�9���$�,\Yb�k����R�~�h�4��W����`��'WmV�Y y���hU�1YAD��+�p�Os1�V6a8�:Y�
��"�[2R�@�����e�uU���t���z���J� ���8�.(93I0r��9�S�?����t�Ϭsv*�`g��N���矎�o6h|�qZk���Y������2u<QLs!�?����v�8��eV_UT_Y����Z��'���,�����""7|��X*�*���2��D����CT��L��ъ�Y2�+����[T��d�B�<4�ȧ�W�ꡪ1on��u�=:��P)D4�`�6$!//UZ�a�B�ɚՇ�34@�о�]�J颊a���
+�P��e�����<�h����r�f\�=�V� LV���s�6��2���U�?�������	m�j��ZRA�2�-�D�L��j��"�B�eۺM�������ŻdeV�4���hP�r��vWՆ}�	!���K��J�4�
V�5���Y�FR�T LI,��`nq���VZ]��V���q�\y�0@Y�/�7��iC��Y�Oz��h���m��x�]�Ȳ/�ky��j>#�ɋUz��h�¤ơ'a��1�\�+Ww�4����&�=I)Γ���TP3
��G�kʆ�����fPoq*�������|B��4�P�[��&���F%u|�J ]h�i�(X���]4x��62��% F��p�eQ��
�����!�g_xl*��S[�9�-�����+	��w��y�T�oEi�$�^��ōCW����EgQ/���Ac)ws�v-��[�n(D��W��&�ԟk��$�,�{�@��C�ğn�@w�Ծ�.ip�ظ�VX)&�{n��$,=|�=��-x����>�耥,�}�D ?&���H��?�����N:���vsG�����|T`ڄo_f^V!��6�|���=���Ce�C��H��jB�F��
��{v�D���3����sO�A��S��k�D%������t����w��wHϡ�/_����_Ș>����V� FM�!�\s�|�`�֤�t�}KY�õ��@;r�|�	lzZ�$�U 7�fr���� h�S�לA��<?Zv�<C�"�FD����+w�u�<�؋�ݭ�Q��"/�2B���S��}�7_�k��@z�J ��젻�����+��7��+����ē�,���4xt���6q���#��U�N����ʡ]�e�O�I��t^��������>�=,=��8ح��<ѵ�T��'zK"�Ԇ��VXssaB\�/ <�b���6K�������(ws��[R���_9�2uz2�o!��%�MW��kf��b���i����Y�9�^��>CK��!�9��A[����?�ڪ0X�P�W�+��鞔��xn[`�}(���(k����J@+�fځ���2UW�z͌l�E(ଁ��a�#�`̘1��(�w���(�ʉ3��&�S1&��ĝ�S�zO��t�,km��� �Yc��g�
�Y�n/�ٙg`s�ͱ��_�xd�\g;��~�̡u�m�y����t�y�k��;YS�u����8�ks�m�79ʒN��� �?�1O��¼�\��x�\q���?a����x�ɜYgJ ��U�� ����88��@PZH(���V�e5�`Z6Q��,GQ�6:��w�t5��/�`デ�a��>�ʑ�ęԢ;*K?.�Q�1Q��W,d �����LtՒS DD�h����<(	57z���)�мXF�K׈�R3��+�� oucg��MIT�~�e�k�mAST'�ыt&�v��R�+���T*�R��F �28���Bo�A��R�M-z���O<����t�jŃd�׫�yif���DW����z�i�����������X&U&��t�l[���,��� ^]�DɁ��L*Ǚ�}��.��!LgQ�E�����}$����2�����F%�.�9�ҘQ!�ƞ����`T����8몳`�HKlլ;���dU�+�o�/l,�e����%�6Uu�R�y\��<��B�M���I!I��՗�S,�I�5��d�o����I3�Ӕ��&�-��0E�P �pٟ]!���!�]�$���`۫�������[,dXB���N����{�<ehb�ꛃ�>*y�Y�H�r�+�_Ɨ��jU�O"�H���n8�Z/&�������� G��(K�/Y�nU�h1�|47��"��#�?0�\׵�W�/WY��z7��!��2#`�;���=Q|���������Wʮ�������}�]`�a.���Hv6�/>�g�^2uJ-�18/������h ��F�ӟ�0&f���[&�z�-��XU\�Y�l�$�ݧ�?��9H	]\X�|�D-��=����� Lӛ�I8���v5˯��Bsv��=�Ry��%4݄�u���W���9�JL���7+��xص���6)M�����*�Ϟ _~�	 �B"YT�5��WA���ԑ�њd�
s�}L<�0�tfwB�����X��9Q��{-�xn���}I!�9{�F�N��d��>�g�z�En��SB�4��l"V-'�h��h
�
�O8<�jQ�OK]��۵W��K�{�F��6ʚ��,]�Ŕ�H���[^{�c�햻啷_�G�q�<��k��otW�㜯K~��x#�-d�ӎa]�kR�t���Fw$��¼Ή
�)�a?q%�7_�2���	ۓ��`��,rA�RCzE���ņ-�".������䙷~��JΝr��ѫ' �O��q��Á��b�*��ݍd	j�����G��
�S#��ǹP)Д��U�Y`SwF�!p����uӚ&�'�$�MʑU���
�����'�D9��U�I��o�;�`��ح���2��[ξOΓ��;8�5�����A���h/Z���X,��;8��P�/�3 ��sy��G�s�|�Nw]:��3Q�Ǳ���6�8�e�v��_�N����:�����e�cӚ�Խ�oߞA�`eZN��u�(�0r�ݳ/�T���آ2&^/X)U�A����0���ߑ�K.��F�� c��\�CX�=�L�*���L�fU�c,�萤��@j�w�6�|��sƪ��+�tM�n�+4U5 �'��.�B��m�-��T(��V]���P[��  e����wt����I�$��RzÓʕ��u�׮M&gu�� 8p'WvMK�\��ǎ�t��"�W��Ç!5%�U��!�}Q����vwh w��v�G��&Dۮna6zI��WK@��6Tz!p�3c�dˑ���[.�^#b��o6���k䆋ϓ�C� ��beP�h��,�1�T�����$ȼ�\<w:yC�O�R��!���J���݊���B�k��ޙ�Dʊ���.�u�+��V���f/XP� �l*�Ke��c���0WO�-�7�k/�Z����`�����\C����6t4{��m���\~�x�|8G��友}S�AlJbd�D�Q�[(���Wp�9�#�莂��E�%8��CWJ�>���`��0`�i X{+���۷ � t��DkQNQ�\6���ʮ�M�ol��׭ݘ���/���d�O�ٝ�ͽ�|�F:(��ꂩl�D�(�z�����U�,˷�A�}�ղj�o��;oI,z�ttTa��t
�|ߛg9��+(1�A�DU�_;v�у
?~W<cy�֯��1�쓔��G�P�
���$�G��I���?��ǯ���V�}�s�����|��2�]AQ��PN�ɕ��qB�f�Q���M����K/�(w�w?�HL|o�E&�7[��b�|��Bb�d�ƽ2c�hD)�f��s�������aG��q,��d��>�g�{/��\�3R|�WFcBFZ�C�+���E'�m��څ�sUµP�C=]��y�����>�R��멇L����;�Ho�"�W�ʒ��#� ػq�5�%ix�i�I]�4���71���AB��）#~����	�7f�H3�4V&�%_��@���&I�{�Z�כ�$�H4W��P�5,����@��7:.��F�f��}5�ec�l�z'_z&u�X���	�7�3�=�a��ܤ����U��0���WxT��M��%X;,Z.�p�"��Ə�u���*��C#�'a��4E���SfJ0҂VJ�� {/c��K	9�Y}��N�L�%�'A,��#� � Y�jĹ��w���p_���<�����`�&�(��dѡ��>�.M׸�@h1�E9٤o�����d8�s䐳&ʮ;�gv�T�7��p:_�dv�c����)y�}=���#&�z��N��c���i'�m>ֵq���p4���������*�X��@X�Z��*�LG�FU���V�� /o�;�����7qMt�ɠ7��F�BU�V21.Ԯ�FJ�J��â%���b���m�_%��Æ�3TB�����U�>�8��TxF�Q�9�G��V��@)yt�|��p��)-����?'G�p������FiG�xM�W;����gl�JĈ�=��Q��k檞��5��D2��/�	f!�&W�vөߗ�S3���ȝ՞��Qb�6�ʒK�͡�3�6<�d�����P8�t�Q�G\���$�/�d۞�wZ�� �� ��⣲��W�p��"p���n�w�� ���d���Q��/[�_�y���d���+���3<R~\tH��	�WG��6��j����yR
�E#�	�h�]X3�ك�s�jW<��b����O6��y�r�[��CK�
t�E=������A�o��p���}�:i3�5 
��Ns���hh���Ŀ� �����|�B+���8��lfēɫƔ��:&��:�bL?@	�A�:��t�[
�?�)�Q��%����XM�N��u����zm�WZ`K=�H��`q��6���1`��|�n�����ߕ�	[#��~�r0��=�o�y�r����~���ӱG���~�8��~U���|o�����a�'��L�����	���`|��W�ف�E.�~������h�%t5���Q+Фe����g����R��}K!��QH倖�}W���*��<����ȱ�4�lޕ43���cR�s�� ����SOɣ<(�?���~�-��Dw�-gϺT��|��_��na��|��م�B������h��	��n^w�1�/��z���:�h�=�Y���E-�^�r>ƴ
�{��FlP�E��:|H�4�ZW� µ96�Ӭ<�Q�;t<�t;&�	��P*��1�p�Ř�J��[��b��HLu����~�| *��3���;�o���s�EH#����>1!���i6χA|���d��Q��x��.�{�CF,A���A��os�ɗ��#�4и�FLN���X�P�ӿ�񸢉�I&B�[��x&@Y�䮆��C�ieM���������4 �{�=W�9/,����wH�I}�sF�a�gƌ�G�E�
�~ܣڡ̍�\#T|<Y$p5�*�j���`Y� T�]�x�MG!�آ�B�Y�(�kӕZ�ӓ1ό��Z^�н�=Z�د�В�2�e�V��?X'@X����I������,�ݬ���[���GudX�R����8��3?�2���v���J�}��Ek��/LXG����.�0�k�L������y�3sx��a�,I�e&����u�ᣞ�.������L���ra�\�w"�2�T�	�aw���`8%�h�]�tEG�+d�1�(cV�Җ���̢տ
/��6^Z�{H�����2��5��@��L4�Sj�4���-��K�q�nB3T$�)��3�
����+�ۚ$h�֦1@���'���~ !ѥ��,�oʊ!����j���*h�1���ݒ��-t~����zl �V-K�w�ק߭���!0$����Wa��*�U�1e{��yhi��?�UfG�03(AϷ�|P�/Vl_p���9��`4�o7, B9G��L�ֳ�J&6AA��':Ir��iD)!D���f[뤌]�wt/���I�$z�WR�n���F�8+U^y�F�v�b���3�׿�
������);�r�X�\��MQ�zd� ��<
���`4tB�tk�&�	}�h�Yj  m��d�ձ�A`"�5>��AߝscVk�f�RV���[!Š��ULkB6>�L��Lb���h�X����G9Z�w��Q1�s��w*�k[���!"�C� ���(�ݩ��ӆ�V�j��
b�8� a3�j^
Xd� �}ЍPfюX]�7SBn�1 ���&��J��x���e������;����8��w.��J`�Z\�$
�vRxg�	:��O��k�b��v��
�L��B��fN�7�]�#�o>�\��^kԜC�;{(M7�"ơP�R��}O�.\����`�#irƔi�GI����!C�p�1�%g��e��#�x��'�]�Kj���GY�f+�A<�	�Į������j1 V�aL�uF����[���ϒ+/�!��
�^�qa���~.���rؕ&��` Ja�f�� �o6U�?�;��Z�4`eR�3�#��m.�oVn�L�>]�*�-ʒ߷�7	~�T��l�\v!��2������-��{�Z7~�}�����<kÂ�����o&{ӯ�P^}�9��%ݲ�7�I+�%�3y�}�'!�m�A7q�L�8��KO=�4����[���-��'ߑ��4�J�Ԧ�_М[o���i����e+:�C�x|�����*����U��_�TP0����
X;�۵��Y��S(��i}�:�)��?H^c�\z�t�9�x��s��YSϒd�bka�2R����F���<O�--Kz�|���XL�����i3�9�7l'l���u���ٟ窑��0[���:��c���j)���D���_��Us�1pvu��Y9K���{�\e�����}�����֘�<��Ka���tĆY�\�M��X`���:�y���,:��n�W��T�oV;pu\�su�)@�پ��k;�ڬ��$�\A��-�oA�O�gU��W��c�-���t&
�(�Ēx�K���4&�S�>��~1L������Λ)c������z
=�ȡ�L����l"4n��&�.��E�a�
�!Ir>��S���Ys���2��>M��J7W6�:(yMxU�+�d��U�*K-�51�����8��sј]Y��A�y-���dZu�-�(�Z�����`pŲ��A�0�� Hd�n�L���.|��2�0��_P�z@��P�w+vS2܂����M�3�j���G�mo��n(��PC�գ��M�m�%
XCѫ$6��'��g�Z�w��"ئr�؎����%|�l�q���c ��a�6l͔�^��������0�E@$�����A�﷖ស���STKm��VA��Ra�K�6Ԃ�`8�j��ɤ�N�x���\�
J|mt��(7����H����f��������f�*������*`f;^t�z5�ёX���`�gA*M�1+�$��U�o&mV�t�����M@M��bm��v�V�.-GR���w�ޱޠ��"U8��14P2je! l6٥� NM�c!�
` �]���; ��	˃r�dL l%{7�L�|~�)�84�ZbB�UI�[W4�0Uux1퉶� swX]�W�V-1*x��C�N����Nn!�W)+接C%zJe�8�5tc�Qb��ѣ��Fq�½4���Ͼ�q7]�8��}��8xL.�s�\8c�:�*���	��eĠ��q�N&����-�~�P/Y'���쳯���!CT���(9���:`1�RG��l]�2z� y��$��nJ�xR�6s�R'�&��z�m >rz\���;U��@B
6+�!H��V�oT�ٌ+~�	e�]�����-�FKzX���KX�^��s����ށ7�W�����U͊��d��7C��i�d���cQ�،']L����k%گ\��e�>m�\<�b�-$��&�E����˫�}�N��\:�RS%x�ge��_�x�%����.�~�j���Qʃ�U<_����"W�:i}�e@t�$f6�Z���R���T�oiVTX��;�+u�?z� �$_���Q�g5N��GeqRQ���w��0��HC����d���P|��4�!�hl��W��������<c�߉%��.��a�]�cIX N�{ҟŷvK��.���2d�jL�3����.L�3�莴[TX�v/�dl� O�r9�����w��u������na�7X�k3�əaQv��fן�`ʾ���Xّ�}pv&�d ��,:��, h��:�I�~[Me�{C.��R;Hu>w����7��w��ُ����,�m�q'���L�f}�݊Ě����#a?����Z�]=_'���@����;,�����-�o������{�"�l)@�:��)i�ȶ���ve0Q4K�^���4]�eE!+�(&gڬ���_��a�̺�<ٹo���)4j�Y�����O�d�o���`x�%ڈsG_aD�	}(g!�~��e�G�dԘ�\p��VXںծB; 5�������k�Ѐ� �	��dL�v�2I��"�F�ѝؔdѪ�hкJs�����S�g����`�tr1�R0)-�W�'%@o�\t�fP��U���Ԡ�?;ӭ�_ 9FfF'�:b��m]hc#�T�v �t-�}�B]�^��>���k�����-J�P�	�.Rx�ڵ���ep�0ټn�A䌱�岙S̈́_S��W���LBt��SJ��`[a�&|��V�&�O�8�h�RZX�JE��I�Q35g�Xn��UGت��j���OmL��Ng���� ��α� �E�e�:��^4+�R����¢;��$s��i� 8k��b�C	�����ي�mF���?� ��yzGWu8�o�I{�k�bʘ���vwj9S���t�1͖�1����.�4VɕrL'?�?(�K�]!M%ш��0 -(J�D&�ԣ�$��ʐ�h)�:,>0��\~��"�sil��9LH ��6���!�"2���f�z�7����ՑƗ^���v��Ib�����^��B�}�`�ΐ�5w&��p^J6o= P Lҙ�X����rɕ�Hמ}�](_���0�`�v�NX\Taa�����4r>�5���0���S����|$iG���J�RrdC1PV��rl5j�	� ��f:�UN�'�/�  R+|
���((�L���_Ø���QY�2�{����N�~�ey��w�W?,���"�����+�H\�$�������0A� 40���0����cWHq�Qy�װ{!͜�]�i���[�If��=��N:oǌ�@�э\�y��Oa�*�����&)���]��_{�y�_w��O�5Y����@�c�7�fM 5���n=C�&h��ޮH#��3�2�l��hxSG�*����V�s��B$8�	�Z��\���%̒L�U})�na!�������N�rl�R�;]�,Ģ��{w�g��)�s��� �d��s��������� ��;
,*B��6k�/c���)XvU,c�Uo~�b&�s����H��Q;��=a�i{OǆY �d �CT�#M�P�@���-�c��ҟ�dm;0��.ʎ�����K�';7vpr��ک�,�m;1�u�����4�/��S��~縖y���n{x<��� �v�x��0<��Jk���ڼ]��vA���R���)��S��A���-�N�R<��b1V�.As��fA�d�Xm��9��_˼yW˼o���֔0�\}Z$���ƣ%ø2���c�$��@������)Ƿ���$�	��wH8�e����˃����7��H��$�B�O'0��Q��2#��ʃ��Q⇘x24�\���|9��
9ƿ��m��N-��{ ���FfYh9ˀ�c[��Ec��B ��ˈc����1l�P���8�e��I��ј#Ր)�}��6�=�z�n�4@����Y�rݼˤ'��H����!�'x����l���ЦY2e`�$z�5��j��"u�	�ѝ�=��Δ&`U`l�J �.t����Ш�MA�vvie*꽥_��)�61����Y�TU��u����)hRcx7-۪m��`Za7��>� /�)F�r��[e'ALJ�^͠���y4+��Μ��\0Mf�U�h��&Lw�}�T��0�3:��w Ig����;�k}�xz
%��V��_zT�v˞3��L���6?��_��3]f̜�}�*�,�'x��I�d�C``B�>������Z�v��0LΙ:�hǲ)�mۼ	��*閘dX"�4� +�C*�~b��J�s^^��3�؛N�H�S��0����HP��4y�?�yH�~����7�9^ЮG���˯�I^y�gy�ï	�F���x�EsU������'/2���D�b!�I/��˯��1�'zXj�8؋�m��Pֺ	�����rC�	]�$�4��%hc�V��\u5&��fañ��;ln���k����3�le�kmn0��x޻����e��,7m04�%��o?�H�lG���
sZ��AY�[��
����x���=d������ʠ�C)��{��xs�_׬�sfΔ�n��S�Ӆ��3O=i���h!B�b��y�I���V~�<��R�f�@hV��� ��]����9��$/����z�9n�z@7|)�)c�����j�=��k��M�>b��se�ـYW���+e��������OR1�%������ p|"�"�G�ا��zI��x��X�5�e�} ?M�toJ鹿�6�r-�>����:�%���w��1�a�z��b��^�T7����"��UFȱ�ij�c8��;�:O� ��:'�H���М�}v��>�[L��f�^�t���m��u*`�lV�Qiӌzj�`�����_K���n}����d��~��ke��ϓ���Y���O%̷�����*[���FU�@}'��5a���xӽ��߫A#0�܈��1�ah�R�T�V^8�hq��"����~�E�K$4�,Z�]1^��|l,e��������3s�^�ʍ�W��������z�X,-j	������-�����g��'��	I	!�Z�-m��[ww��-ԋ���w�L�qw��w�3/�f&��{����̜9����zֳ�,�9���;�5���(v����"�d�E3fC +�E������ Qm��{Ѧ�0�����a���vh+Vq3Y�X�E���^�ґ��%�&:~W�J�	�[��wLd_Y�ݿ&�^�� 5Z\�$m����Uj�������7	���k��gH�Ii �E&�2Rf{W�=�n?F�x� ZO%�s�2���٬�Sa
��-���+Y�{ ��WT��Ο7���#�a�BL#���ε�
iJ@��y��P���"�p�x�4�|s%�� ����-K���}���wrO�j� +�N��N�5Q�'���. -��[�Sc���ʅ]�d	bG����L�� ��
(5`��oV(�u��=�W�a���g*�~�9����2�2d�A:��O��F��[ Aef�8r�g� �H�၄f���D�\�ų�ظ�v;t��}���V�ЬQ�^]�f�}�s����MʶS2��+U�&7#	��Dg�;y�TJ��x���!b/��۷S������#���ګ�76��g_x�u�ND%/4C� �G�tW�0I�J �Iy�?!�;5������~O�o~���d}�M7�9^d{�e��O�3�2Z��S�T	���X�M`��$�
��p�o��B�G۝����Q���w��(�$���T���<L�64�蚖��P2;�~�FS����8�E+�rl8�35�(�6�r��-7�ISP���.�l���v(���~/ݠ��� �a��cs��2}��1ZD��3;�ۡ]�m*1GcGe��mu��y�x�����C�y؉lǔ�<�Η?�,5��;?�^�b�0͞|�Q�s���T�g3O[h?��-y����/_a��:��!Y3Lwyt7]�0��JWox:Z��Ū�ܭ�Ƹ<躢0�+�8�BN�MF���i&���^tБ<s�d�i/Z�{h�	���,�D���j�{�m�7R�l�J���i��>ͳ��6�6w�9�!�iV (2�є"k��s�Ry������5ĦQ�T�Q�<s��)���ʮ��:�B��UB~ie��h^x������{*��=���~7���g�����`��� ��3P:�`��F���A �����W&�>����2���S�'�留��u��  �dl���}�S�ԫ�>4���'&"��N�*@�� @뿨�hA�\�U�1q2�G����YщJ�ñA�Ƈg�{l��6�3��K�a4�a�[aaL��l�a+���&���������t��5��I<�`�馪���&��������>e�&�ŞB�*&a �tZ�g����J;�Pf&�S��By]������"��V��N�ǟ�b�5��c`P��>gkw�ʮ!��K,�p�nt�Ź�^^��m�iU��m-<�;�E5�jr��
��Rȭ^�@F�_ {�C�f�>�IWR�tF�����aҭgRk�h,&
���pJ ;���K��`��	/��u7�b�D8�Q�QZ@:7X�MV	�hn/�����Rr��n����C�Iɢ��G�V�BF�Q N� ����@��tS,�����]� �R��{�7�u��r�8C�� �`�C���
g1U2�4jj�`��th6�8"ǦNI�
{v��9j�=�q�o�30�����S�Ǡw}��
HS^�+p8�I���ZO��k���m�?Ǭ�Mӗf��[���r�X1�v�� � r����ٯ~�}�3�r;�OIۇ �l@Rؤt��������ƳG�ݼ���6�� ~^s ��r,(F�<^Bgb��|���e+ӎ`?��n8�&��Hj��W�����yݥ�%x�Ѭ���˺����?}��8J��v�U+�
[oz�q6)�,2KL���t�F#$f�
�$�F4iu��D����%v��Yv�_��C�a����҆W�0(�h�R22��®�0��zL��ma�{�kER�jf��ұ���5O0�ꚫǔ�h����A,u�g�� ��׊j6��tNR�LA35c�b����]�/05mZKO����贳��{PD����<�n)����գ�l;���|��	��q[�Gد~�]�x� �߶��������,����s���Wh��1[v�Uv��K�n��׮f7��J����Ӑ~hK%6������ۤ�:7�:��P6�j`��C^^J�Ri�y��I��(~��F��Mt��L�lٙv�5�q���L��mt�Ѵ�J3H*lf$Z� ��l�"�2���Z8]�o	IC-��|��I��ɦ��86��DG�3OD)�UO���)GJ+��ur�d��:(��8�Z췛F�+��8���T ��A:�b�7����z����)�?��>�;??�s�s�0�~�|���>?�-
��g0������
>/�O�y8�%��{�{,'c��A"	�Iw����}��Qq:��]&�����^�%��D�M�Ǵ��N�2��?d��͘����"[�v���8�&Ϝ�i����+2�& �9e�=��f,
m%]d=�w�JL7�{�av~�6qn�c�x�1�1���)g�&�NۇI�:&T:�4��{���>��+�Z�Pi���a���"�Ɓ�h VS�q۾O^A��7
��Z��}�J&���w�V�i��Ȋ�ഓ��"֦����nb~zh�8��m�E�@�!��q�.4T��'�@瞘6t �-��Bz(�
���`a�h ��Kj?8�?��M�x��Iֈ~��Ԋ�����Q`:b��:�(�	k��g�/��`z����(eg@N�)h�Jk��sP�0���0���Ʊ<���0Ε��6HkE�ʍ"mU���������F��U2��g�n=��7Qg��u�zz�����,���e�b~.�Y��ǣ8��h����$wyZ�[ɇ���	��	L��*�"o����J���c	�kg߆��JLQX�h�p��tBbHJ�FðIP.����12j��D���^x�VMG]2݀���c���g�sh!+�H��v����j|�V��n��mǎ��4_�Z�kt�?b�(@<��hs ��6��u�{: ,QlBZj�dq^��F� D������1&����ȝ��D|�ة�ٱ��0U}�	mo�ؕ\�n������{'��G�+�`����Y1 ��*J�s0A%U�c�ъsl������[鑃�M2F�\�4q�u�^�c \N�C'���S�d�#O��VQ��`���mB���;��C෍9��y�n,��Rrfg��8�g���zL
, {��Ju���*"��	4�'X'Pl�v@~)>cqQ��ǵۏ0������ɲ��f�����}��{��>O���0K�]s�]s�eN����}V1�,�!���҈�f,?��# SX��2K%������}о��Z`B�i�aJ��4�0]���rhm���jə�\�Mx/f�Ww�M�ފ�:�n�E�?��ȅ���崓I�����TE�S�|��4��Y�F�QM6�Qtw��W|̊K+�����L�Ǔ�ͤ,�)Eo���c4��0w���S~9�V݌���J��E�ar�K깓?R���Ij�Xt]�|_�L�R��n�!u�T��	����z`����_��D��~�)���^�YTF�	����}��e����a� �A��	���&�9;ٺ�w��tp���?���T?c�����������ȻO'�	 ���T ��N�����Ս �G]k$�)��d��\>w�k�߹�-;R�l[q7#��ӿ�ysf�a��
��7n�U�w9�е_�����Uo�K���	vb�:i�`�z�?8J�b熩j9��m�/�;���W��SUJ�N���U�������W��H�R�H(͆��`�.$Y&Ĳ�D $���Y,ylD�l�����9���R��Q���ض��C�~	J݄��V��)	�#X<ԥ�f �(����'j�AFZ����o��5�Y���-1��jGP��V����T��1ahㄢZ����'���d (��o������a,�aqVN f���m�FCH9H�Ik��@h�={�霬x���
#�T�f�H�KMM����K�
��GlA,��p]{� O�����a�h��t܀u�U��1��(t쌠���:A�+�B* ��-Q+�*;���*8�n��1F��c�mobӱ����F�et&z��!6�i�.��U@��F�e�\W����WiR�B.�����b������Uj��8�dò����FH���XYD�CTދp Tf��00�꠽����eãO�d�-����a�aO���J������[('q]a/b�F��ɤ��c�������A��5l�:"����Kz��4�$8-	�_�56z�����`�9���cŶf��.Z��f�ٳئ���G&c5@�U*,WS������μbg��M�_9x�uE��U�R#4�#Y�3��`&:fX��~s�]v�G���g�O;��m\�� ��E+-�F�Az���c�Æe�ye�;vn'	��vJ�Ǐ�[&:��S&!�Ǡ��J[=�I7�+�S�K�n�kǊK�t�|O�љ\�J,1��*mû�%�������D�G��S��S}S%v,�S���Ȳ��?!g�}̾����O~�}����GWg����m̘!��o|�{�a{��H���M��=�0��S�˲�⠿�H����s��7�6jh�}�cW�Ա�L0�>��{��-kb�M ��n�u�J��y�"���!�E�qMJ����h���:ʇ��rhoc���N:Q��kl񒉰���̌�B)Q��	̞3�ˎ��E�PPr?�B��?ik׽i�7o���[�N�J�mt2�Өu��?�vw���:�U@zǫc�2�ҷ�a��O�����_�b�xV�o�I3>��=K2�";p�>��r���9~�˿q7���er���O?x?:~����d,��󃯯���H쓦�z 6~�[����u|j�ұ�u�j��3ؘ
,,�}�r��̌
늌�`��0�n o���Ըi�l쌉�wT��$�fJ`��	,~�����N�Qq�C�J�|w���2�+,@Qx�yX�r�W�~�^�D���W'��H�_AP����^�uB�8�T/]�l%���	�ǉ=ET%SD��G��H@	�Ys����7�)	�B�cmፈ�ә3�k��BY���\��I�Ò˿�HBXh:1
�S�,t�U/x����A���4u4
X�<'D�S0w���º�_qL!��T:jgb�E,��f��a��`J,�؂�Y2�X��(�VP�g������6J��\�̔t{j���|�[�20yL���a�d�Ð%�^C(u�i���[
��6�k�X�P���a^� ���*gaJ�� �"��c��*�Ų+����nJ�@��ZD�b�$��qu�$]��u�]Q\+�J�">)�R\D,W-
[�n��`EJ�^Lϴ,8�J5a\��!i����`g^i��#ʞ�\���9�u�v�$�1��F���D����'���#�������b��%�]z4��=�t��K5��M�����q��q�	 �&ѸD�:�� �`Xׄ]Fe�.v�-\C���bYԙG�U������k��؎w�;{�9�[m^K_���02D����o
_�,��=�S�������d+6X %
�pt�����h�*�~O=��k�/�;�؊�ш�i�㫍��A�>֢q~�Qr-4.¢�c�Z��AW�o�(9#��}�+8��X����)3�ɕ%���1�S:=m��'�ڪ��µ���r�Ŷb�B{��;l��u4��x� ������׮��8�t�P��Z=�_�&FLv(zF�S8���H���B;�4BcH�b�86O۶;-�[�������Q�@(nN:1~)��H9��t�M�:�Ϭ�ͯ�c^�᩶���]d;6�n�<��]�evh�۰�;��exm����s�.��SFZ-���w�]�o_���؍�˯�؎a�,Z�P6
[`��R��of�����7K�=�yoE����܌�_���ǐV��ۮ4���ox����А�jWR�c�Ơf0���n�Ea��1�UVn+cd�X,/�q-�5:��l�+R����{��-�Fk8�Ǝ��gO?��%�XNdZ��E3�2�����mb.D6�j���uL���W;m䭷\E�9Ѷ���< *!�����,��3m��)�[�c��	�V���vs�2�J���r,�d��*-�~��`@�1��2����H�A�~7�6�c{���6óY�a?@�*�!�uLz��ˆ�y�~0�������,����Wn{����F�Ń�=����_�y_W?���3]�B��E	����jT
���w�� �;� �D�C�� ��E���<X	v��'j)!�gX.L�4�3�V�=���3�s���a{�)awʮ���1i�3<`�`a�	�dVV���"��6���d�Y�;t��azފsm��w#��0Y���?װ��<��Kh,)t��v�b:��&�nD@Ee���6@��B��Yp�˫�m�a�]��a�(��N��c�_@���X��D����ƌ%݁)i������>��`�w�y �$��\�J��40,v����25�7$>'\�E[z�5���(�[RVL��O_w	6-���^�X�����V���t�VS��#��rA�a.������ߏ<8����U~[�#��S�%v�� v�c&��/�2�/��y?�q��4�SOA�CM,�b���DI����fҪ܏e��ƛ?r!�N<�(kI+��q@H�H�-K���R�Bk+A�	�r�m�v`�v�ď�G'���EQ�r�o�Z�	 ��(˦�}�u��j:�������8w����#��x6�`�x�0*��KvHb����MC4Dܻ(�S��2�K�(�da>�]�1�XQ,`ᘯJ��� c����2	�q=����z�?c�TH7�,Y@o�ko�杇a(!�����tߪ<�r5օ����t29����}%,�u��p�Yi �n[���\y���l0t-u<n��չ�1Ǎ�^���L�K��z��Q�c�ʳ��Fk��O %��v� P"�0��9�H����݈�S���4ܴb�ЄV��Kl�`CU���m����m@V}�}����bll~��ّ#y6q�H�ޯ�M�67�%�Œ����|��{�T��Y�O�7���<�wӸ��f%QzE�z\�pI�1ϕV,��N6��w�,�9�f�Z�(vY�E�FU����G��H�6ZfN��t���t��t�Y0`�6,�l��uvb~lp�뼍�����~m��ܮ��x����"����?߉���8�mv�ʕ��/|��
���匚f_�ڷ�XE�}�G 0<�Z������b�'�ۏ~�]۹�-����W�����`���w6 ��y��Ƣ���<��]��E�QOd�`�Ei)#w���� 57����"W�mb;QDXp�hf��d�:6^.�)�`�捖��~������i�R|���Z����Ϛ�s4��w��ٴ�^|k�5�cw�p�呥Z��X�v�向��}n��$Mm��(t|�o�s�N���$ -���I�U�%��};̚��	)A��;�m`!�w���a{����P����:?�A�g~ ��np��y�����Q�œ08ﻄ�������&~�ɻw~��]�z\ݏ���A��x5��Ͽ�����Ã|}h�*��磾� �u����%�!�V����A&�M[�Z1]�2�L��v�Ǎ��ͷ�Q]x�LFf��+��w�ƭGpT�l����9g�}��v�h��q��8]��egd�&�_��A���Zx�s����||�V낹�K3�U��m���`�Xۙ`�$�>�[$ŵ֣I��D��ݔ���H�@��P���ת	�kG\�l`s\��]fi��ʏ���x����e�W9��F/0�ʣ*q�P�O%���˅]�R*7(��E#)������S�#l���)�T�T�}�oG�I�xf�u�J
��J�/�:�S������Ϟ����yk�3mTwRL[ !F>
h����\��tK�����]9��0��Q-������Te��D%�r�*�N��ᒥ�i9��PF� κR	��]�A@MX'V-��6ܱ�Л� p��m�i�gs����*:��,;'��~R�"g�Fv������nǆ��m4e�k/_nE�iG�pj2�E���5�L"z����w�X�)�'�	5Y;sn|
�ń7�E����l(yzǏ��u�1m��_����)���RXTb�g��[m +G|e�	���ϖ�@��@>��0JQ�ĵ�L�_��p�,�1�'F�X�A���Q����r�|r��LSB@�D��G) ݗn�n�x���D-Wu��WC#JiU��q�2��ᥣ��ʊ�	]�CD�4b`�� >����!	4
��wӸhC��l�� �$nzA*�`{]�}���/��B�.S�	dZV�$�GE(��ή{"?���z'�΀����� �x�.E&��ɌU�����GiiiH�F\c��$��G^a("�XH��a��(�Wq�[__e+/Xam5Ev�����!I���~�~��oss��}�~����-��V�E]Z�a_���e�ٵW^h�؈��4��J��E)����V� �9�����E����O�iul$�C�K̡q��6��g��6�~��������L<���V}���=���ax��%��/��:���c̽���WE�ZL��ۤ�x�W�9����X��1�8�w6���<��:���wmמ-6��L����c̉g����ot�V[-lW;�7"4��/�>I]6k�JJ���z?J�x��v��7�U׮��_��5����\���3���N�ݳh�\�_y�;m�\��X��۽��[��,U���2��^�H��g�@ċ+�6���y݂�c��K00��`�N?��H����<U`2��x������Y??�� ��5̝�=���K;����\����2�*%^2������I�X�+�^�&�6�'�p4��\��?�͟,#���a,�P�,4Ǐ��Nx�1|V{l_U�mZ�&��3llz]\I ���\W�p��t>1��{��ڳq�-X4ך0~���7l@.͕��V��'��XTz6%�.{�{��͕��QS7m�*��6E��{��w� T���_n˧��3/��.���mm�n�f��@t-�!�R�g�ҕ[�4����(yX<*�B�+0�;SRA�Pu09&�X���(ԫaD�A�Ϥ�����JT*"8�ļ8a��ܳ�����������]��|[�=A�< Xev�A/���$�����q/b_QH�Y�q:���s�6����48��zX���1 �H:$���7�R��gG�n��sg��MGo�*=H��c`L��{��"�y���#o�sO�׉�i��|�_�\Jm�.tz�q�t����ȁ�̢���JM0�&�Co�Ե��;�a�wo��~�vl�.�v�V}x�[`k�D�@;��R� t�b	��Ǟ�����6g�(�OY3�X�z�Ba9%�׽}"}����P��c�����z�wV�9˷�N_a/ay�>�r�u`��� ����'N��N�w3����+��O�XUH����b�XL{�P����NA6Pi� �ʓM��K	.��*�秕�!�.�.>���g7�.آ�$�ـ0�\l�|�xyf�L�z9�:v#	SO���c�g����[/�[':�8�)9��W�<���w
��Jl
�}Pc�ed�eHne2�橸�w��ݾ��F� �/�+����\2�~�V��럝ͽ��r%9��U׸�2����`�������E�s��w�:`�4�*?2���V�m8ْbϵAC nmh��:v����7�����V�NW���kk���2�p�V;k�4�l���o�V���\��W���wލ3~�M�=�z(�%�W����Rp�}�Y����}Ǿpۧ�kny��cO<Mi:�~���X��s����Q�a�u�o��u���*��S��3���-���w ��k�ƍ�'���ay%�����߰����m��,۰n3�b�}��Y��q�i�a�a�F��g���?{�4P���X�0Ռ�r�d�2�W��f��2%���dY�31��B7V����"�i�ᷢ���s05�`��t۱'�v��Co���"[��f�>,- ,�8J歌!�j�����_��׻1���ΰI�'�}h\{%2�A���eIo1^X����~�����``��#��恩���@,�w>^�n �ּcf�:�����``.�A���u�������<U�|���=�7�&���6�ZM�@��� ����(���	@B�J7�1��B+j� ;Lb�&t"]<�i
����N�����]~��z�)۾q�Y�˜��k�+ۤ�q���66~1�����/:�@���W-�풋3�O�\r��{�u۳{�]�|���d�� �/y�����8�O�(�p����;�i�1e��I,��,M�C�2��rlML*�H4گ4ڳ+����Gk`rwA���j��	@�hrq���a��E�8׾;��� �xB�u�X@YHU.QdI4��	9.�� 2�w��ts}�_%��]�����)r�>!�e� ��J�l��i�g��֬Y�-��;c�*��!6@��F?p..�Me�-o�v�4����-t]�������[�:�T*P���IS��n�-?�	���~���9���ˮ��+���A?ǘy��UV
kgq;6ז-_��n�]|��uι������G�赣��O\w�}�ȗ<��)�NF)���:|�b�3q��Uv�pǳ�6o�BT�����E���jm��C�a @�y���m�2uNe,2�p��YMH�E9�9A��ySl�˯�ˤ;$�kvV�)��;�K����{���3gڍ���[�=�f����~��q8�c���P6)������j�q؋4[3$���;O�l\�I�h�|��b��ET+\jc6�Y6v b�@��i [����,��8�%��	�V)��Ղx�SF�����Y�{K�'��.O4.�脎N
��M�o{�ݵ�4�����A����U�ɵʒ|����m��v�?� *�&�p��Z��JB�]�5��aD�U�+��]\%7�R1��F��&Mԡ� 4���6�Ґ!x��yG���@���P���{�8Q@�N��w;,a��v� �j+�H�D�w*�e~�q�{ȍ�]^�ҳ�����uD2�`W^�����G��X�TbJ}%s��/;�UR��'di�������N���+m���l6&�7��5ۜ_E��sVR��4l�e��\{�ư��D�&��?��^z�>GO��mٙ�6dd�}�#�3�:l��Ih�J�(���l�\Uv�gYd[	�q�}��Ѵq��Mbw��/J�-m\���N�)���r��4?t��%�l��وF�1kø:�N���R`z�I(�t���� � :���Y����A�����g���6�M� _}�ugK���,b���r��Ob,e}����F���O�{uI�N6�)hz����%�` �����<|rҢ_|������ H0c4[���O@��mx 4���;X�k�˹��\�7�����~P;���{M��~��|�N�T�|_�ɿ���{?�Ϟ�m�{�i��~A?�C�0-M<����r�vS$�e<LDC�;�8� 9���x8~-�C�p��9r�e����lhD�]w�E�"�p5�7��*mhE�(*+�"{Μi6	����� {`;�l���v���Z �B��^�G�Xb�g�������>��;ˮ��L�����%�s���8L�ܥg-�Ӧͱnl�s��	L������J٩%�T4W�	H�w�	l�V:����0p~Pw�T1�"�_�}ӻ������S�taz��؅���+��&�ݨ�v���'A��f)m[)�U�zм�*�&؂�e�U_[n�0%ݼoXf�\�v��dU���/+��#&��ES�N��baXд#�"_r���v|G�`'���`ϧE�c�T�i��(�E�� q�6z�H{��W���m$F�����Ik]!�u�P8jJ� %u���F�q�`-u�|~1V��S�B�0;3Չ����4y��*�4�?j����: �C%���P�J���ࠝ�x=�Ҙ��{�!�=`n����XI��RKi��I-Ƙ�����H /*ͪ���m���m6�� �,���9��q�B{n��vΙ��W��F{E��}�s�̨뮗b�g_>�-�����P�%Ӆs}e���*�vQ�o�`&��(:�y ya�g���ST��%�LV.�@�FzDi��w:>�6J��l����.��X�@���1h��]���Y7��"+��ӧͰ#�� �R�
g"h�E���@Gd��E�՜)c(#�ɶnZosщV���R�J����<�D��&0��q���C�	j�w��Ca�<��H�-T,�c)����z��-60��g7f�0h��iA?r4ߕ�t���'-p�\�T��l&�p�Wg�������6H>�����r�A��7~������� �����؉�x�b�7��7vľ�ݯP>m�������?��)��;�}Ǝ�"H�M�����a��J�좢���_��R ��h��z�l�)Lex:����poF ,�+����Y��ٜ��B��Dޫ���x>Zmִa�,���樓N�'�p�=�i`�s}��#h�F�u����a�p�7+����ֵ�[��;�`1����/ �d���7�]�4���j�N�q�;�!����]CE"��d�F�g|�j���Q�AM9q�cl�4�΍�tto�&�J:�����|�P~Ps�%����O���� S�����3u���{?X���?��3���
��޹���,a?��~�T�q��T~�l����[���`p�����4�̞w=|��O>�.�C�0�p\�c����HV��hl�����gB)%�9�GW!ޱ#f��Jd�ݸm��#��sW.�8�	��I���%���.G,��p\���m6�v�a)C�o.�U,�r���l��,�;�)$�{
ӭ,RjD<z�0�;��t�՛��n[66�?����;�.=�4B��X4L�"�%����{8�,�(��D��m�$�����k��:9�뺫;���\�`����O���M$z}/��^��������F#�m��z��zЁ������^�q���e�̂]���0:K[��#RCs�,a2q������.C�D�,�X���J���f���%&��alm�eBGGI4�V�@h�
ɔ��PN9m�,=|$LF�&���u>��	((�S�)k��T�¤�?��:�f�H&v�\4Izjڪ,��%�7Jr%��M���C�T6�hN$O&�����<�=��d>��{'Є��F#;�N�0���v��s��j�v#1�E!�,�N���]��~�0um���؏�s-"Y�B�-�B��y�^��C����<b�NX���A�q�Į�:�����]��k�󜽄Jn��b�j���3��݋�R�>��)��%S�j<9�8:~[���27��P��D8�/���U�:)m'�T�6P���Wz+>O^r#1>_V�:aB�k�l�X�`HM覬��B��ؖsyLp<�����f�������u��D����3��#�c�q�-^8�~���a;q���0y��i�! �����YK	*&D��^��+I��pǮ͉��d�'y���E#�a�di�/��m�6P	 �X�B��r�W���1x��8>_��Ͼ�R%i��VD�i������OU3���h������Q8��sCc�߭Xv�m۵��Zn�C�_z�U��b�����k?���{�2K�[;���^`�C���/.�x'���P����Wו�֍�/�`��8���|�&L6���&ƎUb�z=h��`ܥ$G���-��.:Ӷ����^�
��%��z�G������9?}�<J�Q�c�.�5u�F%����!֧IJ��tw�\� �/��2��J�W٠�]���K�|!�\�Î	m�<��I'Ռ4���(�.�/���4]e`%��
U`7'��kS+�B ٔ	��g;Lsp����~1��8��d��~�w�w��]pW�.�� �,~z������@ݑ^y��@"�~#��a~�7X��`�>#�����\?��w�z F��AX�S�O�[�|�^L���A�����R�ݾ���?�C�0�U�ڇ>�����y�
�\ĆwT���	��<(�2^�I掟N~\�Ӗ\y���G�7��u�)��{�-��ն�����|�dλ�B�4=��r�V$6�<��}�Z�C����G a6c�hۋ�׶-��:��~@U���Ї�[Q	lMy�}�[�	�#���Z;\p��c9�q
Gd��=��k+g#hF�[�ݢ��`a��� ��H�� 2�9q"5���J��N��ZP�sf�Uv ]Fr�v��c��}�r����}���Z�U���������mV-���bJ���h�v|�m�RT8o�qc�ٸ)S�͝��w1�Qn8��Q�4I
�ЩZ�b׃�S��G�˰���"��2S��I�1��`�U`���;�p��h�rm���C�2l`fݔG�QG��Y��F�5$!��FI���Y�J��P�c���*�p�|tU�8^2���,��y�)��Y>��VX�����O`��6ݜ�tS�[��ctO�:'H+�uj�UmE��o7v �=� �2k謶(�d�]���<��:�:hEd�0�>�N���!֧D�I��Ыf�k��'�\yw�\��H�rIh���`�ak#r8ǯza�}�#�ڭ_������m�_|���5�����R��ݸ޾�_�6g�{��B�F���3��0C>V��Þ�r��uS�v� +���q�TV�&��
�Ҧ�,�r�8շ26\7�(�3���(SN��oj�$3D�k3���]I�
��lx"�וY�XF���d5* Z �Fp^f����;�����JC{� X6��tS�l��E6���{���./��ӪA���19�$�K���0z��{�D C�@<�ۓ�lV ��vbI�5)��1��ƌ���p��ag�jd��6�҄��ԟDʠ�S�3���e��f�u1È�ø����F� �"��p��W�X]��|�7�t��M���v���-�w9��>a�l$���ê�z�n�i��������+v�g.s�j��Xݰ��l�`9�4&�9XI���/��FM�-�q��t������v��=���~�dE��o��m�#�o�'1tƙg�2B&�������4���<b�<z�N�?F�S]�*�.Y��m�s�F��ϳm8�7�:}��SUX����t�	ۄ�.�C�HW�C�6sh�`�z �j�*`��,�(C�lT�]B2�&�Æ�� ��U��[��bH%S�MM2�/�2r��}@��y�0�?I���`�F��� �R��j��"��<����,*����E�R\0`�D�s<P����E��������_0��G��{��=�\t���{ ��������:O���w\� ��<�< 4��|���A{�痎�_��_+w=T'��(�g��~pn�N>0���@'r��w�$�Xx�_�&�Ȳ���r�߷s���4�N������[�[(�V�0�gp�`YF���Cl:����{G+dP��4��	6y�Y숒l��	Έ�*k�h:Cm�굘4N�e�c���?�(��14�:�B�˼%K��_B����+�aȵ���6
�2Z����[a'��d��	��ÒD�&��)�����Y�yEn'I쬯nik41�뭬6����_�܅�z�AwF���`�2��Y��ݙ�R�U���4�Fס����)����J���:�[1�p��{�{�1��j���E����v��gB��SM�A�t���;�o����o����r��r;�[~�t�Ű��"�n`G��h�]�h�]C��C�<l?��M�HN��Єԫ#�rM1ݐ���;��p޺��Xia	����������!$޲e�˲a�����6�������:΢���j4l9x��/o�������2 �G��F>r�8����;jY�
1�o���jdj�{��ka�Ck��p���g��[��1�G���}�8_I�ms����S�"Ϣ��J:kc��u�S6%�\Trߢ�VRr�Pn޹�Jj:;*������4;X�Ŋ�� ���g�;'�
�@������ƒX�� NI�+`҆���5 �8���cU�@J҂D���"v
@�NF1n��C� �'4w�qh�d��+��R�������'U4F��
�� ۑ�`RY%�'ΒT>tw����ʵf�x�xVb�_X�t��i����@Y���?���Ɨ.	 Vj� �m�K�����5�#a:�G��EӦW��uA��:��D�-��4ias톲HW0�[qq1��X�	�����K�4i��k���z����"�Ե[��jp�M��p>\���l�_0{���z�]t�
������Ζ�u�͝5�6l�a�'ϳ;�{��6f���K��p��0xr�`,�27� ")B< 7�ڀ$#��w,�uYNs�ޝk*�\�P��M�&�I&Niw��vK �����o�N�2���x����{m�ks����gG��h��ل�gYD�;�m ��bG��?��#!De|X������҄E��[m�y%�\S���
�U1����x6��kb�vPfO�c�+)���NŐv��Y6�,�"�7��@�����_�|A$���9f��h߁�� pݳ=*C�ƅ7���{JI��y�oN�!7�;vUZ�w#h� �>����ey�(l��ǿ�菭�Y��{~����c�������������j0@���?I�>�k�����J���A�=0S�+���c��Y3w>���+�����U�E����H��D��=t���B9(6��eو���+l�x��$ĠY;-��yv��u{�p��	v�Ev.<�N���~����*�.���f[��mX�q�����+iP���{��l�bK�n��6�<hG��v�������o�Ŧ�.~%�!/���̙d?���?�3��^�r� �q�d��VJ\�hBY���]وH�	8O��k�Ec�&��a�'|׸( @�1Ձ �
���@�nG7T�
Z������������c���ӆ Ze�f�����/��#�z�	�Ɨ?a��Ǘ��&K&���F=�Y��wa�W�U�֢�"ʗ?�+c���lw<�����3v4-��)�V��Ɉ��A<Ԕ��v�U+쌅K��@7�K���ꢝ���
]Y��|��V��F&Z�cG���Hm�ȿ���.��
c�T� ��]�(��V~X	I�?�&�)�&P][Qty�)������n��Fk�,-Qe�Jl��?��~�"�����7<�LLu��9S�ڽ��`�?���ؔ��,ذXKW�2)��~,�rk!%9@��G�[e��D�|�c��\��s�+*kaC0���A1�0�.��6�b��Ht��i���ʌ��ቄ��/5<6O�ze�f̆e���YN7P-�?��hi9�x��� o*�u�R��PK#����.ul% Ищ#y%k1�QХðO�}��\�n���i#�)�����~r*M,�,�b/Į�s<)�;��TW�7U�<��KO�뮺Іd&�]���τ=fA��yʥ��A��P��[	������#�ĭ��7���-��	�d�Wd�D��(fe%�NH��<���d�V�O"^b�mj����nIS-e�""��-�^�,I�_pv�YtJm6��z�� }E���W]
hk�N��g�a��	v���X1�����aocG�-e�:c���q^�e��tl�0P=�l���d9�{�J�ɤ���=�n�ص���w���G-s�H���߲�^ow��Y�	������9�z�	t�w��8J�-H�0���� lG�О�]�~�*��E�cO�N.�:�?c�Ă��ͪ:\׼����)�Uܵc��t��lf�����m Ia�%6{�$�w��Dw��v���C��H�f�ߺ�[�H:C���������h]y�E�xRK�o-ll2^f�0Օl#�RE�v�x^t4���D�bU� ˿8�AT0��g��t?@��`��T�Y�o������^6��?0���v�5��W�.q����X����������w\����߃���J��}�ƪ>-����߯?��Y�a'�o}ﭩ���>4xg��,;�:�{☨ʋ���Xj�i/���a���tŝo�^y�m<PH@n4{�������Ut��}�N,ۂ�S��4d=���^_co=�
�W�۳��B���w�潖9f�%�l/����Ax���a~I���ѭ�%���8{c�a�(͘�����;�H����ze����a�<�I��jx�<���R��tD�z��KZ�p�4��	��)�w�,؉�H���>헷�tc�C�h�1�M��]hz�Y*GbJ�!�U�=5'�ȡv�E6��3����:��;�xxc%�!�f͚��y����ٶk��a������̴LJI���V=��mܰ����D6�K���&Hg��B;�Ï�n-U�m����ƺܾ��)���[D�Y;�xZU��� 0Z�ʊ�9����;�}��u�Q@��	��BRm�&ܾy�"t|�I�$Q�Z�~�F��ǋ�Eq2R#`ZNs�Ui�	{���n(ݖg�윅�u�	{�L�a��ج�l�q��!W�;�`SW�6�y�˚0�Bqޗ{z� ���&�� ^7&/�K/z�xJ�8� xj�������g�s.�KgX��ް�a���J��M
�y7V��Q&d/z�J2�WI�8���ܩh��T���6��/18m"�E��S�$Y����B�mt��'P�iFYjS&��d�]��h*|�b�\�[�s�M�v2���R�/=��B��GC��K�h#�C��.��Xdh{�)��K�8�	�n")��g�1$=���n��|��{���i�8��q�ݣ<U�Rb3b"a��X	�йM��@��d3����/��M�)�K���F�*�6�*�l,�������*`&���4���즤�Μ2K��F<�Ѝ��H��]����@��{v���$��`����t��;��G��w�	��d���!;���l��Km�>J�� ���F �B�&EdkDL&&6�.T�Z��(A���ѥ���D�g��i<3尐���Q�co�9h�'Oa#��9+�}�%!����ўm�9��֮}����I��6�>�P�9a��<���H��:�������	e��E��E� ��5e��vW=�G���δ�?y��u�D�<�5�]y	' ��@,i1L{؀��v�5i�8bO<��}��ߴ�h{���}ac�{^�̢�W�b�r����ͮ�>�<�fBf�.έO�`o��,��������@��>�-<y��{]?8��{�0�8��8��������}��w���w�~�?`< :��� ?��̉����|_��4�>6���&�@�k����k��D�^�6�R�Zr�4�J'!�#�O�!�d����.�q�N�D�N:&f��3��8��N��_<,H-�!��P�$���]
�j�)m��fi7W#m��6u�t4eh�*���%[l�8+���f�1;P\b�Lĝ����(��+���*N�ME�Y��ōf��xF�s<�j.���a�ܴ#��8v��!�IC�i^d�����@[6�RQޜ�P���%f���ڕ![)?8)�n�s��&��t�"̏��'�:f��ܥth�[ܸf����{Ȋ�/��\�hR�7!.%?�ܺ[�-у�=�^,²Y�~��?���;L)j��
Ka��'ϭ8:�`��9V{b���w���W\lW`�8n������ ��揾����
Y���?�f�,�aBw"&޹��C;�����&:;�����o��!��ߵO���s���o�k�逾��6�I���|�di(�ӽ����2bb
ʦ��Vne�m��k�l�i��^`M��z�[Lf�m����Fq<G� �;3���T��NroUr�U�V��N��#`�B��I�o���(�̟D9����'Y��_�$6	�̆Ws���q�j�q]���W9�G�{��^<5dQ����vlG��o��kW̳7v��[�Wα�X0w���M�;Mݔ�Zm#��3现��O�tu�6�����Wz�S�����b�b���0��Ny���輺1�l�ڪV�''�[�����esQ���q��f�^%&$Ⱥ`j*qd�­��v!:�����h��$�`�K�\Gl�4a��$��[������'���DDn?*&̛y���O���PYR`k�6h�
�޼o*��4�?-�ǎ��X?��Q��_v*�q?\@&Y��j�w��'�6H�	vݗ�7W�s�������b�s�����!cѬ�~
r��tMظv���zrOa�##j���
X�64�N�v@k�Gн��O����Ԟx�e�&`t=�6����R���O?�y�s1!�_���0L��˟}�qm�`�r������Yi7�tsS�����\��v�Wزe���-���o�f� �Kl��6����gA2�w�0y���ɔ%C�D+fC�ҮJ�bgj����OL@z�v2��!����h7a��J�#5y����ˍ@��b�Ǐ2�h@�:fd��+��ӧ��j���(�ƦwQoa���AB��cOQ��x�^����\ޱ�^�3OGu������<cZ���M�g�O�s�������:�1�^��@ '0��>��H�y�n~��?P��Na�z���1a}VY�Cp�&TMLl����=pｶp�|���X�(Q!��Y^�K{�SƸⲫ�Edj�%2��%���~��F�6�6'���,[f�5��ecy�_�A�v�9��@�<d��d��E鱚.�Fi�p�og�bRN�Nu�	�� �%�E���tB���f�щ�#1��D�rfؑ�rP�̌�d�p�`��eai�KF��v�H�z�PUjUN]h_Ǖ&V�c���z�r�l��n���Ӻ�`c�Zja�!.&����vh�L�mF]f�� ~{����+�Q�;�0y�t��/�bt16R�:k���7�YD,�o�쫶e�*��v-�F<����v�|n2L;yr��SbB�%�8���9}2�/�^�����%v��t ��J���Ye��9��1y��яR�����нg�o<���^�;��.��:��I38�{i�m���6k�{����4.<�":�m�?��;�Ǿ@�K��"Xz�� ���O��졔{3({���30�̛3m��ag8��f�]r�U���s����v��?���KB�|�$�&�% ��X 4L���^�l����b�0G�5�4۵� A�[i,j��i�O d����L!͕�,hB�jeEF��iė�0��f��k����Ćmք�����D�w`�ph��T*S8x4ڨ��օ��D�Q�������d�0�\ݍ2N8�@~�X�(��zY��(�+��Ԁ�x�~���HJ?1�D��[��o��h�T
�#��@E�/O�%�E���Ơ��3c�8��9V�X�>�U	z�d��7`|�xw-ߚ�c�U��Xs�m��}y����$� �8*�n�J�t>��ViQ����[ư�؈��!�L�����4W� ��(�	�9�J�~���Xl���Tת����smh3�(�EY�,���νG��Z��b�F�wt�H�r*�F�y	�cG�������e���ڡ�$��X���r��D5��.Xf%��[�ړ��O^����f��߬7�&~϶76m�s8��/�7����nS%�ËΜ�o�A���Y��U��d���W-ڗ��%*U��&�X�Rb���c�|��=����$¼�`Da?��4�#��N.�.T2Je��ۭ�p��!� '���Գl��	H �p��U�����k�̼&@[J9T��thb2�'�T�,�d{��Ap�� '�T�-��E�?�Opil���L�}* )���%�������d��Į��@��`�w
LҀ�k����7�`{���~��ww����|
lf`wx��̈́�C�
�;TS�b?�1j-�=��]���8�,k$~�]Ӑ�l|wv���K*�}L�0㦐]XC���x�t�߆�&��7�s)Ͳ�f����o��R:K"�Bt~]�EGY4����d��7̒y׵өSJ�����F�=Z��.2Vp���H>R,���Eh|�G��vR�j�A�6,��]쉺��9�p:��^F:,���.�s`g��=��mW�p���ad�@�"CV�)wv���"��F ���v(��F_�ޢ��J��@O����H�ӽ����?c���$f�X��Q��D�����+/�c��5q܉h�Sl������tR��B�Q��DD�x��m,�8�V�b����ί v�ö�#���nя���肋����6�K��e��.�m��u �J���[���-�m%�-;v�������۶�G���%�RW����f!�c����p����C~`)��H�%uÎ���9{.��f��N�3��~�yj�iR@Ў^/�4Ya�E(\�ԃ(A{W+�C�xY���u��L�p|/��4��ACA��89��<Bi�pn-�͔�q�'���N�d�0�$�f,�S��EI`,����g5�Ӎ ������֭1[��K�r��m��/[��v�6���.JO�
��GJc1�Rp=����c[��J�x�qPZ
l1�k��)X�JPp�=@��.�-�u0y�����H�N 
3�ai���`cR����" ����w`Ր��i�7�z ���,����$���,���L �lN�o��z��J@`G�M���9���1wn�هs����ޙ�\9�ۙ11r��f3T��>S�4U G-�4�PJ�]�H_b}�^��X�a��A7�q�7�����b/���9A`\�+��Ss5� ����rN<���R�#�/�����Fʮ0B�F� ��m�u��.�r��޳�أ�G�;\젺�ц���Ԝ����O��'�m��=Cl������ϵg����ʋ֑�&�[ �?�y�G_��:���ꈜ�JI�a�a��34�,˗+3َV����8�~�SK�]t�������D�1�f�����N��7=��%#D�!�S����hq�Ͷ���XJ��VBlѹg_���"���"Ǖ�ET!X+�a�Za�ӱ�Q�د6��q?Õe�����59�.�����`��~>���{��|0��w z?��<{'��w�z��\��k�`e>y�#�������?�낵j���߰�]O�������w��K�=O�	��Ӌ����]��{꿗~��dc�w�'b��P�F6�=*C�������F�
�_�����or0�X������z�E�ȵY3&ٛ�;�˞�����[Q4�I��� �2�N!v���{��[��o#3�l6D�����/Z[�T˝d�,N2(�3<�&��Gͷ#��C(K6��۸$vl�ee�T�o�6�E'�6�/g�2�G$;Q��.!�h�t<L����2p�o�|J��")#��Q�P���<Mt��U�x(���*��<�����U���d��:/ܶ.�̏=A�v���J�"�Oh1KLpIL�� 5u,Eu�,���E-:S~>�m�eZ� G(~h�-w�8;�S����B�������W����pf���^��U�Xܯ�lZo��	�CLR�e%���&�сɗ*��*�]  �#���y"y2�l���$�l�7sp�ߒ�P�"I�qum��3o�{}��<}�e�F#nj�	�8�!�����~��oc50��"�-j 	9v�'>K��8{��U����ز��L�mϺ�v,�=,�7pK�p�,�Q�&��iw=���/]j͉�v`ٍB>�E�����F�u��bgO�h�f��
�g��9��|#ff�3ݯ,$��R<o���KV`�mE�V�7�FV�IN$KVI��6�O;��=����;�ž������ ƥ6l����)�Nf���T�,���L��ls`��)�v�:$3a4��7r9����Y9V%Ǆ�)��uS�# �M����ð]�k?`Xݒ�!��ٴ��y����������)����U��&Me�a՝v�G��t$������*C���U�Xf\�4��!1T�
� �������I��$�ZW��`}(�=O�����T�EY�\��j`XR����4h!<'Y���oe��;�H�+r�h�U�U��%�1�8V�U'�UQV�4�l��8�$?w M ��ʦB�R��U�X��4X�ʼ-�Baқ��舣��R2���3xo7��&�]k����z�R#!���U@���g^ wP��g\��֍Ɖ!��6:"3��tq���O�����n1f:�g���_�)�H+!�t��E�%�h���b{�ք1�)�)݆�2���C����B7�b��cAB̶=���m�P��Z6$at�vr|1��t�v����&ظ��ݔ�k��K��,��"۸��eX�0��12Vc���٨	�I�'UFz�n�R��(����٪`f���Z�&���8�����r�F�Px ��]?��^H{x���?V��{���,�yTO�1�����¼�s~����������<@|~�������kp�h�ٮ��j0�����d��ǻ�Q�Ee��>`�_3F��˾��� _�i�$���zW��ur��N�4oD�<d�FK	4��Y�GG�`oo:b;Ƀ���3앝�დg���Q��v>�?;vn��l��~?z��F�2�������ZzO�U��h�Ə�s/�����!�Q#��t�x�D�rd��1:�~��z;�7'��>v�t;��������}���Â`t���i������Hu�������������	'�P<��ji��kuT9�����Y�IN�ܻ>��<N�/�����0N��� �إ��g8�4�X��杔�aiz�s�P3,��R��<��̳1d;f�Cz���-�2o����o�09�!H/"`���`�8����v�f���(�9B��qɍ~(LS,k<;uؒ�FWB���N�:|�"�ǏK�i)��1��o�
�i�]�WP8L�Q�w����i49iv����W䀍��[��fB�c)	���Z{�Gl$e�O�|��D;J��V,)��|�͚�	H���Woş,ߎ��������<���v7��4؊K��������bk�ژ>k�eg��fAb��j����_:��_�o�-��,wx��Wb�V�AY�}_y�
k?��VLjY�l^Ý_�O��c���2[�h�-�h��ݴ����cV��IO�H�` �x��Ϊ�Žf.(f�����cS�I+�}-�<�5n�A�s��Hl  9�Fr�b0��­���Yg��5��hF�6Ѩ��i����͜I,q4��/]�]��da��>"2	�V�	fJp&��D	H�;��(e�*ܾ
/6�>z���E��qo( ��h~^QQ`{7����G�̅��?���3O�d7�%���Z�����희]��.�z�/o�pe�wf��M�Lg4}EqNz�䪮�PJ��(%���	��,�}�p���*��t��Fr����>�T���C�����t�����݋%�f[��i�ډvJC%���ת�UM7�4����2��Ļ)���I�t7 ��p��@y���&�aڬ6q�+'�t���)+Vڟ�O�AǥDB�1�.�l�=��z=f�� ���&@e��,5*��Ǳ��6lc8'�
J����O���.Un޹m�.+�5� "�8��Q�$���<��Ng̰��\"ȶl��,נ�q�8ȢI���QT���h=���A�t�?��>�&�4?��#���W�7��qY&��~H��%9���3ڐjs��b��w���T���8���JX�����<�?&�2��٩_0#���u���6~V�{�`����3m��\~�_7����L������`p忿�k1h<��m��Ȇ�B��u��8�fI��lN��I�����������>
���\���PK��!o���6v9�������#J��^x�&�i�7�km?�E�v��+l����<�u�x��kd!�^�N���f����B��%�p��������#� ���xX�0a����}�>�06�6��׾��[l�HtEL��,]�v睏�d<ˮ��"[�e�lJ(!����B�Ӎ�'����Nߦ�&"u
u��!�(X�&&�p/Y�)����:%�����^ZZԴ�J�&���P�^���d�C�F��j�2E���$��ix:&&��|Js��C�^���￢u|�
��gz�ڏ\Ϥ[jo���ņ��I�QU^T�6,��gG����0�@�qP
4O�J���::"��0n9t/6��l�u�&r���p��aDη;������E��e��q=���7�%�c�m���pO���n����}�.G���k��_�u7:����;���.w��[�m�<r�{���6��CX��N���W�h�xv��4�Q	������g��c[(��#{�؅��؝��O�[��3/�*0��t�Ԑ�5�,��.�<<�
��(�����>��aK?�.��{k:-���P+(���,`��P�ʱ���뻎P���	dcK�f�-뤌���4X-��Z�b6(���]�v�So�3�� qT�I�v��#�g#�k�a���w0�7�M%��x�Ė]�]�H�iA����m�$	���F �X�(�(�c$c:��^�o�Ze�hJO�q��(�!����Q�Ah<V!�0����\�a�b�Ʒ��϶���T~�[�bFi�j��%�^��Ne����y�I��x��`��)k��2�nCuN���oGM�ןg�)��\�ձ��įKJ�lZT�t_j{w�|`w%#�*J�(9��,=���k������@�:T{{�$�w��	��^���l�����`����`?��U48��и��8|��eyv�}��,ͯ|�h��0��i3�X] �����/��׾�C��/�o��H	Z��<f�xN{`�V�\h=��M�2�V��!��`D9^�M�<�]�Cq$]�u4�65s8����a9�$"є=�ʆ�@^W��g�6�.��H{����X�[I!t��r⢱ ����)F�b���X��+��"	�K�e 3�����
3]�B>�b����<�����$�������r�3�q�b�E�}]���Ԃ���J������<�z��1�돩�������޻�쾿s�ܳ��>���I�>�C�0���X�2hk��];�n&��^�F�$�����Sքp5f� ��=ۭ�]sEu �寻�yҮ��2ۺ�m��3�h��I��b>X���p2�*l�O�i�^������<`	SmȄә����atA���LGD�ExC�m3Gu��Zv��rn��O����ß�l�cVNgW;�):��pM�,d���Š֠��?��0!i
݄11�nw���s�-G��eB�@�S��҅�0�����"o�p�D���Y���6l��ƨ�/ �u�^;�v�Y�8�$�X+��w���h�x�$�Y�ǰ�����<:�����N'��5۲�M���k�y��i��t�e�>i�pk <����D7dyU��iA܌����#C-�n�Gy�X�`��l��bKQe��.{k�V�,����˗Pu��]G�#Ui�(��@�mݷ���M,~M6	K�HJ�o�ۀ�,l�~�H�0�=�9(,Z�)Æ���%;��^z��Ўqi��*C���VkM&����Mh�nYi	�U� >'�Yj{�6�?�^e�#f���ғaLz��"�O�z{eO�!�%�x����!���#��c��m��+�K����x�}�ۿ���/�1�N�I[��Zqˋ�_��[!4%���W�e�d3��5E� JNK��{Ģܓdǹ֝��m�Q.f�_X�`����A	<F���y��0�埏���n)��q�ف����&O��h�Y��K�C�F�h;���0ZM�C�϶v��(�O��V��Ё5�Cy��'VYc< ҅���|O16�}�6�x�!�!�	?9½�zv*��~kROin�0���~W��\�˔:��W.�D��0�-��-�b�<N4��	�!e�!�+^�
 Y�L���v�����ҘFb�µ�Q6,�Utb,�)�ɾD������v��<4�}��r,�lS�	�mS]'�7w��;�~I��	�v맮�[>��M��$8�i��o���w��G�s�d'b	#K����	�a���|9ny��ҍ�y���G�駟��}�K���5!�+X�8�.�MX3��NXx1S?����ՖH�d"㤉l]��t"ʍ�EEx�qD3vO;}	�wD�նح��Ɏ�n���I��[-���q�]�B��M���6����k|���>�����`��b ��]0���TG~=R0��ց� S{��c��c=p�_Y�?��g��c'j��<ؽ�<�A~�T��IX�w�j?�|3@����Ϝ} `����� L�N9�w�vC����c�l�,F�����O��a����t�$�Eۗ>�)�H���k��-H	1+��[z9M�]��(�Q�N���}��?�"�ٳ���˴	��<;�V�gη��\n��ǋ����j�>c6��^��G��������~�2(�p�l��gη�k�%������S
��_WQG�"3��lYЖ^��w� �ϱ��(�������c��M�d6 (`���c>8,`�+ 
W�Y��uҋp���0z?sW-`I������puNL@�,�葹��[�o��D���ɓ��H�d��W�gH'�V�hH�k ѱ:�;U�\F)�m�QJHB3�$���uR/H��>�kj��T��ʔ=�i�hA�3&_�:�,�L��]�[��]NL�zO�%}���K h��$��� :|ܵ��S�q�Pny�"�A/���Yǝ(�-�Vi��r;K8���U��|{Y�h%���hR�)����C���ұDI���/�3��&��K����f/��ֶ�L9�e���iZ8��'� L:��ƃ�Da*�3�2L�U�^��B݄!x�đ0��ܧ^ @8��B�F�S��C�'�8Ѿ:�Z(3%����5��	�̕h0J������`D��Kɦ����H"k0�p�Q�bh��̕s�[�0����R�L�q��y=�ck;Ǒ��p�0R�F��B�%�f�D�R����l�9]`�.o?��� �L�Z 4�h�h�FwkaQ����g��K��2[�/��Y l��鏷�kW�E�c��������=�\�@�a? �;_w�C`Ua���h:���a6��b�E�Y%6 �0J��h[���D��X���q�����*�U�������_���c���?a��[�E'M�o?�)����}�v��k��$���o~�KJ�� 3?��w��U���yLW�ј�4�*���n�D�,�#и��4%ݱ�&8}��?b�x�]��k�<7 F�}��jr��O��❎�y���A��]�ײK����;!߶�T�ņj�C�
FPN�j��f��Tcy>� �9� �#W�'>�&����0t�ca�/����#x��O@�B	���(�=���]��^��@ k @���*��������������z��{�������Y߬|>� ��h����.�
k�[���r�凄0%�����$vǕ6i�H�`�%���,��EJ�B��S��l�#��quQv�4z�Xډo�W�	�_|b�5�O5b1_�ή�ÒrF��x� ��,E@s���G��_��-�W`��XL����q]O@ws�'?�BGI����'��B6b>�:��$�n�(�,HY ��R)r��d��FE���H�a,�����~�g�4���6	ܒI;�W`-t`D�ԄH���{�r��+:�����S�@8�g�)	8�Ӳ�VmJ��F��I���{��n_%7v�V�Ed�	�bI�����n�Ń�XJg��+�[��jk`��,9�GLjjم#���&�]u}=��t�J���$i6��'�;Sɞ(�*�D��5cTU�z�P�mjT����qIWp���4w���J:�F��p�t�[�X)�އs�aU��Zn�����7�`q]#�\�h��	�t��8[�^@Ȣ�m}~��H[�O��	9��XkdQ��q�C�U�Бv��l(�2��4��9 �T��B7�=u��z�r{�w�1<�p���*�0-�D�p�H���!/�c��j��; �u,�V]�qiG����X�1*�1%'�mH� d��G݂��9{U�k�h+cQ���'Ƥ�RiH/�Z
ަ-�Fֹ��8����!z-�L���AϼP=�Ct�,��Ωt7Vb��H�5	��d@tڥ��&g��6����Zj{i,�a�e��4[I�qK�0o�������go�����ͤ��Z�f�,��U�W����ɦ�����,s�z��8���@���L X]�*E
����5��ؙ$'�H4`
��/�`�-�dգ���"�	z��,�M]Y�q���G9��>(6 ��FIRsh*�»�l�[�^mg�>��a8�\*ۑ��и�`B��;����}��c�M��j��tb4�Vrρ�,�.��tسO��7^�Xw��6���&3�y��T����M�_� �8��݌e��R���5�:s��s�"�NK�i���*)���Lj������+C����iY�:�`,���E�A6�t�q?:��@ܑ�xt��-L�Z�R��2�r%G�_���S�}�Q�gF�����	��~�����3T~����@G�&����>a~��k
f�c�����t����� :�5����u���ro���_�g}/:���?�C�0
�����B�p@N��P�,*��709O�B b�Y�x�D�aR ��9��{w[�ރ��~h�6�L ���!%"��c�>��%�5[�8��5�
hˏ��A�kvS���A`�a\�wn�j�q>�ꃖT��"\�Sl���v������}�v��?�c?�.��\�TP�Q�g0��H���-M<߃=b����~H'�a�u�2��#���X:�:: t��a.�4��N���h��B�M���,C'B�N��=D �bB�ck�l�+���i3GD�H���r.%��J"��r8�h,=�JP�"KY 3�&�Z:<��Df2u�i󕘂�QSE��" �],�B��y�bqQ�VB�vئ6v�ٙd@ƥ�8�`�J�h~�������0v�bݚ�X�;�*OH;��<"^�z)X���TWꉧܢ�l;e/M��i�T�B_Z��Ӱ�/0�e��lfCV�~��7�u� ex�����d;p���l���GK�Hy��\|�K��.�B����ְ�U��?*	��ÐP���Ya����n챝����O����:�<*��u�S��a��m��7��W�@ΑpP�+{�TB����M�L(�T˂�qK�[ԃEJ������u��5�7�jh�����oh�Q�c�j�r�]�}�_�w�̪#����Y��I2�f��N�_�زt��w����N�r~VWAw+��$��TU-�ni$'tP����|�G/�y�����_������F#I4�w+�T~��-	�%��O�{�|��5�M���K��J���hyeH�.�*�<*�Z߹X����Rf�d�ۉv����rF�4� @�twq���jJ��a6e�Zܓ}4���3�`哌{?�>5����˴����]���m._4�����<�o�8���k��[ov݇?����Ql����ɉ�|Ɏ`��N)r�`�������}��=�`cX� n�&��H���>	<�40d �WY1�|�z�m�e�9p����z��x4�o�f���(S؄��F�Y%%x5@�G{z�š���}۾�_���횡b���J����p:����܃6�2���9-��yw���;=����gEcHN�rjlw��A�f��KN�������U=Ƨ��K?�������ƶ�g~f�Bc��K'�~��<�����v��'���	�c����������9�qʂ�w><S��/,m�k��	a���<a�8�'옳�Ra��Xx�4�d:֘aCFυn��w�x���@Wc��ʢ���&1$�&:���Zh{�%�b��S��79z�VE��4��{:��_����i=�`������t��'?y	��͖�FtxB�H;g��LH�<�	s�옕�o����C��k�$���RXi�hj�����?	���p�V�3gE,��	%ԁ���+�EU�S�ש��ʢ%/)��kL�8��I"
����4ڳ�ӥv��v�	�m89�jߎ HtЄ��
p`�ag)Y���L@w�X�%#<7n<-�Ă�s'.����l1�ˉ�S��;�&�f����k���ħl�I'� �C8]76k��H�u�&�e,%��*�]4׿�IXv�b���L�X�dx)o�f�4�Fp�M�5�`�$#Ը����2���(���Tv`��|�53n"�41j4n`?�-�D�	��N��l�"~���*V���d{{o�mކ�Q4�Eb������_Uy�v�{��\���f��4T�e���ТT��ý��q~Ř��5b�z����,ц��r�a�`?|�l�-�X�NJ܉,ha0�*k���Rq7c"�����`�q�9�^JӅ^Reif���uHwC)K݈��(�1u�Q��Y�l�>&2�Z�`,]'����Nw�=Ҹ��~h�ukc�I�i(��GH8h��ԂW�ʋ����3�?�>��a�˽�u�1F�<�=���%������-���H��$z���դ���/=�r��D� p�
?~�F���eg)0-ݢ|���fx6zOu*J�N�7��41��$4��1��$M�W��.��"0/E���^+�(��hu�rok�ܼ`�r����vţa��CI/�إ�O�e�
Ū��e.:d<�z�-'�D!Y��d�;�N������uܻ�mʔ1�yڰ�(>b�vފ��O@Ȳ���6���3���ӑ܂�1�X��_�5d�2T��c���s��:�sK�s� 
@�����+0�ͤ)c;Յ�(C6�93�H�(�m���ZM�4�F�O����Xb\)2`)o9-6nV��6!l�����ځJv����=:4�׉���\��m �2[��|���������~V�>�}n�wm� ��{p�����kH�,��8���?��@������s����ߵf6�~����� -/���?<s C�|:Ww���;�BX�s��ͮ�)��ۉ��@�Ŀ�	,9P���ْ�J NZ�z�]�[{�YWa���ߙ��3��`�\@һ>;1P�Q�]�%]����"�Z��bk�Ũ�-*f���pT�?����BuU���ɖ�.J=��s7%�)����%�^�a �Re�p �� R����M[y����z�����҃Z�uR*�è�1)%����S/lb����a�6��PE�D3����X���,~=h�ja�a!��=�Rd"���X��j�i��T����T��a{���ddR��~���Y��%)t!I�'x�*c�j%g2�^w
w_Z�����H}
�+X�[�����d���3}�]����bz?���M��������=0z�<ˑ�Q� a�c�ċI�N�k�������4���x2�!��,\l.�Æ���壬�t|�JK@}��˞X{�j��Y m�v�te8�7�� �D�����<��h�X�j����F���p�0a[a��� �t�z��Uc�!��D���������	C)p���a�Qd�S�]�b.�&�^�W�Cdf�i����u�}��)�����TV��J
�L+o�R��g���11q�uq_�@��Y&l\&��,���Ĳ�n����hk\��;�=�r;oE�� E�m��n6�Y���3��%�-�0���gZ�-�ޮ\�Vh�ʎ�,D��(6_��N�0ޕ��4��#V-�V��<�������#em��Ue�0����W�T�9S&���x�p��0�#�*�]ހ�V���Уj�P�Tb�؛��Lm�G������?	���ߌK��C�����a9������bl��%v�����^p�Q0"�̜FI\H6�E�ݰYjC��.�������?��q��O�0��5�T��D^���.��D9�!A9qi�8	�V1l4�t���0�MU�䅎�6�Rli)�0�q��k��ǟ����ǵg�>�}� �����l}�iS�W��@���t����~���л��k��3S}kb��	~�l �U������!�1k����y�q�/����A���x:_�8��,��:�kབྷ�wN�M��4��)�y��3�}/pl�7���U�����~������?�݃�����`�0�ׇa�|KD@�*�
�u�ie�l����PvFQ,
!t߱갈��!�lDɱHd"�ω����/�}G���,�W���Av r��ӑ�(�{�9@���=	��1�D_��c��!<��8;�v��赅XLQ7l��YS�3�iě�X�4� ��q�Nb�h P�� `��@8V]�^���)��981)�/%��KS�=����r��X& �ҵ�*�@x�ڞI�WI)蘚�����%Q+yJJZ	l?�$5/7���4S�T�EQJm #��7P>T���jw��H�R����єl=:9	�3ӕ	��,�b�+6� Uɱ{�&~	�n�K���%cB oR�c�3�>Z��4����Cѽ�ly� ��>�(�C)xZ@T%���m�����=�iT�A�g��E*� ӊ�&���/�\���a�ֺx�pX>-R8�k�����Һ��ӇH?$,�n���Y���i׮2۸n�ˍ�qX:.�tLu��9������m�aI	����y�1�6Sa�r�p(�%�aS<�b=%�N�S#d�����~<�֊�T8�	����k���42�0`�FDM(�kyY)Ϊ�����\�B()7�eaB=���IYMa����(uQ�TFc'P��g�G��D"�j�z��V�Í�\d���?ҰPccF�����X�Viud��6�} ��+��=���>�~�ߤ��Ih�R�ƪ"��j r�I>k2�L�5�� e2YM�/vS��s&�<�b{��1��D)������<~�d s(ٮ ���/&}*�,#=Ų��]�q�K����>j�_��58%��������F�[�KϷ�~���Zʼ���$�7ov1o�D�m������ow��oNO8e�(�6y�}�g?��^`+�[F3
��#l����6#^�Mb����ߵr]�+.���z;;>	�/�Е���M���?fl|��S�_��>-��A.)���5�b�5)y���ډ��c,L?]���8��dI��d�S#�D��_4}I��Ƹ��:� ��H���>����
B��~�r�¼���)~O/ﳃuY�i�d�1A�=�`�?}t���T>�������4?����@���������yd ��?�IG|�c���`�z����A�Q�LN��XӯZG &�B�����v��2��Ee���8�Ä��#��Eπ͘%������6ʂ��Y�'d�, ���{���pI�|F������%�D��10B1b�|	�e��|�P���u�0:�����',5=����Y���CL+��8��&F�Z!��	��x�L�9�&c� `f���a{}�VK���ä���#Ţ���wE�h���,m�vq
��9�1 ��Y��>Z��e�P�̽�:kp����������\���+3Y�#��fe���i�X�	�ޱ�EEŰ�H<�Ҙ�@�(T�A��1�AR���B0��h�����3"`�H�t�,��̕N�n8�ť`��q<�r�J|F���X�V�1��rl8�`X(���1l"�
Ev&��hJ��J�z1>�,jr����e�6t�gLm���,�EF$M�'�[bv�fu���Nqc[�euUZ�b^��mz��x�����c�+��;��ϞMN��e� 7��OL�h���aW\z�]u�"�6�1T�;s�~�S��??a�w��=�tE�Z0v�D�z`�,�����>���A"� �1�Y9���'�<��d��HG��x��)T�J��Ÿr��{ U��
��ݸ^���n��i0�e�n=:���
ˤ��Fٻ���Kg2z#��V�Fں�p�\y��6}�H�#�?���0"�
m
�?UؽH�(� _�.~`�X���ɗ&P�i�Ā鏞Q�W�9eNq���y���PL���Y@������a�����yj������ W�������͛l{���±���M���H*���<��ܻ�_|������Sm��͌�:��2�Ӕ�3ik;��7ּfo��ڲ���ԗ������k����`F�m&Y��ǎ�� �ӡt�b�¸k�!�A�Ьq�H6J��q4�퀫L�>y��x��� �����N��͏�Fž�3_ǡ'�`��������}{�ߞ�ǟ|����!،��M��,WؓO���s��y�m���jG Ws��q͏nL����������9��3K��1��Y�2���
We0�}�N�wO���c9�㝣�����#x�o���[?�D�z�����``;����N���v���|h�bD\V�JQګ �f�� ������)3*��K/u���۫��_�eG-&c��4�Č)�ؘV��e��<�Uo]+��j+E��H7�L�.�����+ݎM,��8��´[
����q���ab%���B[[�=�X8��Z�l>dc�`��M+.�cQ��E�����r^>ʈ,�3m���!�VF�h�D&�XJ1t��B��kg��q�C;�xʃ2<���1�rPy��tv��`���i�eBJDs2{�<:���m�-Ee]Lj! �H�M�X!v��mefP�"���Um�{%@���#�U*�􅶨��%P�P�,ی�#������������o�̠@o��;8�F��FF��[�[�kqn��ˀ=�բ� v_N��}�=��8�*���$�'c�������ܲɍ#�0׭��e���3���?��a�6�"����|��V�D��ka+���t��N�]e�1;�n�Б]q��B��缲�@��FNi��%v�_�b��&����Ѯ���3s�͝:��zea׭����?쏿�e#J�Q�L҇���t��&��ptu#�e���^Qc)D�b�چp[i��- �H����b4d���b��4	�`�	��P�G"���q�q����r��r�8�8�~�W+��75D4�yi��Hī�����ar3y��?�͙1����V����	í���Q U�b(�%U2��r���I��fg��n�tNer� �ɇ}��MuJ����<��J�b��1V.�3�el�=�%A�8q���N�1�2m7�Mm�R)��k�P_ơw�I�=����A�P+.`�>֒�#hy��aO�L�S~g=��l�l�)>��X�v)��}����p�}�cuMO=��^b�U��UW]e�7����N����?go��h��"�۷��r!���+6V��%��|�#�IPRT���787w�Y�?n������9�DK�X�F�dsnU\1��x��1�R�m���6q�iD�Ͱ_~�=�\�r����BLf��kb�R�f@����:i�bN��=�I SG����Y����oi)������d��������0Z'���3p�@���%?��~��a��?9�����y��O����^� ���7 p>�N�C�0�|�#�!s�nv}bZ��
E�XRYc���St������/��9{"�WCiM��i	�tu��A����ˢA�DF�M�O֐7A�_��n�6��b;z	�E�N�^l'���M�tSz-Vm3z�1Y<�	N��<fZ.B��
5��ZB{C  �1��9�3}䆫Y�����&&&��J@axB&g�J]m�`a�#�'�n��F�A�CRz)&�N�iH_&���,��L���T�H�E �ԎY�����[n�˽����W�DQ��U5��;�0�v&�W^~f
ww�Y=e�Nb�"�{�B�)�vX���Ԁ�^�1���ǔL��ʒ����(�"�����ױ.x���@��2���v� v���c$�8
VO��2���H�JU�\%P&�Ҭ�-CX�ͤ��.4Pm,�*+j��Қ,�a�:�y�����ۍ�]��\k(?h/�^mò��>�y����B�8�*���nZ��$"+�.9w����C��AG�D����!�9"�>u�m6,����i��N$Zk��Tp耵-�ng-�F1�MU�Ԍ/�l͢��VZx�F�f�U�0�8�qN�ـ$$G[ɡ}N����j�gՔ�[)w��@��:��׭���S
�݌�._Q��*W�H�,fP�#���E�䫪�\�y6Ԙ�H PH�WI'j3�8�C*�n5hĪ�3L��NI�W���x����_��TlCs���䘍1�߆#�Q�����p��G}�O̡�O�C<O�/����Ա^�0n���sMs@,�(uGJ�t��Q���V��q4!Q�,D$��W#�W����;���҉�\� ܫJ�Z��,(��PV_�uE���Ȣ4��É�|o8����Jd<�n4���Sl.i$A��I9\]�_��g�K滒�}�Ȕ��Y����?��B�w,,�hۃ8?&&�u_�f���������� �8�)o�����g:Ϲ;����x��Ȅ��n�A�L5�4�tRK�AMFj<),(�e��sͳ����l����n����K2�.���3�`�Ip)�:ޣPY����FV�W�'�6��8��P�R�����S)�0��Щ��NƄ�gڧ[u'����A�������>���<�;�S9���5��"�A���~we?��:�i��_:�����>V����}h檐,u|�S�I������TGe"�:��<�4{��=����ka)C�;{�u$���a���nVIRx3f|�S�#�o���Lo%��tZ�yPq���~��I�����&�/�s�(���E'����]{3C/���BQ�-�~Iw�B���Z:�M�"���M�����DNd7ݔ94����xj�t�@�m���k�	�Ùx�ړX�����
�у�hG<�����u)�7�Uk���x|�ͯ�QB`��F`K�B�w����v�^;Kא�Β :����(�18m�� o�\L5����РU�b��(MY�P)��d���BIЮ��)��wbaўL١͒�A���]����>C�:�Ĭ%�"脊�R(G��[�04���7�V��	ۅ�;e>��	��QZ���� �N�@��0n"�7�D�D	��v ����J��r@6�+�"]I��0��U�(PY����M;}
]�\[X��L����w���=}�Ŵ�["ǘ3t����_��3O�ǟ{�Rc��䐴d���|���u���ۿ�P ���Ȍ;��;��cF٦��]l�/~�m����D�=�"t�����&۰�������\,?`��ŀ�^�h"χt|p�0��3�Y�\ Z�T�e�i�����uq����>�ȌUr0ٍP>U���p���SJU�X�&:Y!��b�U�mJ��	�����A)�4Aq����_0���u�]�v.�_YI�+]O�0�N��@S��D=����g�>�\����\�����gR:1u�F��ƕ�u�S��J2ڿ6`=*cf�n:�Z=�n��A��]Q�1cdVJK�;�uY�Mܜ�sh�貪C��XSN�M���Bʿ��0�`=�'��
p��ٌ�C�֏�J1���T�Ts�̘C��yf�9�Y��'?��có�qXuK��*)1��ܲ��}��1�^.��b�)�
�E��=�ʸ���Ɔ턝W؅ןg�}�j@Xݛ�ߔ���86L�<��2�3OWq[w�y̙Ͼ��mX��V\|��ߜ����&1���v�p�ru��uM�`�to����Q����Nu �W�<U`�<���� ~@p*`���� ��������t�u��ʽF�	u���PO�xN�u�z�ˊ��/�9����ݯ��	�_��]�Aû���XK���Z���@X��$�F"�v��j(-8s �2,�ʘ|�0����^�45J����(�^W�X�ʫ��0J��h��Nv�m��H��[��nhs�S�19�s@��z09lW���h4Du��w��(���'�K��&���cz����W7�Ug�r�R�J#ڧ������Ru��~�?�Ab��j�a�p|Q��i�a���A��&��1AL!�t�ݎN��P>1{%����tfC�Gæ�< �����Ce�A��zl���n�k�9Id�+�����Tf�bm�ȴ<ױ��Α��`h��ʭ�I(��C�K�K�K�)=�bm�igLX曑�Ӹ*�hѤ��5���uK����Rh/!�ʻ�BD���p]�B�j�¸�m&���8�=�t2��ta\+7i�_kf�iBx/Q{bj����nT�����'H��0����Y�z�����5�7�4��v��S^p����2�f(*&�i�h;��%��aV�<t�Dk�fѪ,$ڧ��6�l�ugYL���-�3��V�in��s�,`]�kŲh�q�9\��46t�.:s�MN�c9�S�;�@�\��N�"d^YS��,f�)x�2����_%�f���R�1��>}N+,10�:)�wv�;��L�<o���i1�\�fcOv$2���;��1�5 �v67�U�H��Wb��W_}1��������-�&�b�ls:��'�P��dǽLcCT����p�+9��H�P����߽��������_�F�~���������f�)\��;�RG'JT�瓱)`�3��݊�@��n�U��xMr�Fm :xM6<�G������=�#K�ne��Q�d,�ʑ�#�.�+kG���������5��oZ��M�>��G�m�~ ��xt^h;��L��j`����f�U^�d��V��}�ȩg�=�䣶b��%^B��S�<D[#H]��	�O#?�ϔZ���s�ڧ�t�Pf^Ȫ�����w�A����||��ط?�I����xG����J�K�$jMy��?�F�VS��)��tlʋ�����v��f�/Z�^8�92��B�.K�~�9!!������K�=tW�������
<V"xq��~ ���I~��π�z�o~p��l�8��ؿ�{���gx��T�w����]�8���ۋ�ta~'�w�Wύ3"�ϼ����.���z�� ���������=@|}������m���N���{�������L?��ߣ��.� ������ �Cvdk0��Lf���yT0�]��$橎\�%��[����_l9Xb;� ^-t��&N������{37�L�b5T2��*���6�]�oN7:�8:c{Y����h�EK���]_S�oQ��dġ���%�S���皀���|;u:%����ԩ���n���VO@�e�����o�m��Y��DSF��V�2��/1e�g��M�T1V�09=!���Qw%C�����x���1[[5�R�b�h��,v���X)�H�	�FtP������2"�E-�\���J���k��$ /B�'N��{��e$�S��>���UMd�	���^	ɸ��حS�q��i��N���Q�MÔ�����]�e���d�J����&|�������F��v!@h^/�DcRBI�X��w���'B����bր � ��9��`�˔�ЎN 2�=�UbӈuI�gE�s�Yx%�}�
',1}���8.�.^��ri��b�����@�5o�`k�F���n<@�hw��K�ʴ�3�����~���3�<sY`�\x�M�/IZ���D�<��[�^ec��m��	U��5��b��Ev��)�5��d��]?i��n8�a8��u6�g?}�޾�6�]��_��rT�=��k �9$��6a2iY� ���,).Lc@e�d]f r��t�-�����Ɔ ��q�/<�q���N�?��'����Qn�=9� h8z? �.5��5���,��\��/���g��bG�����߾�{/7�{?�W�����;=��/����`O��(��`�Ӱ�{\'/}�˽��Ke1m0����� ��z��2([�����@�8���[͸W�>Fr�����V�j����9����F�'-�*�R�Mىc6e�T�c�����4~��R�l�Y����nL6�G�V�Y�"�%�s�mԸY���k��� �E���Rg��t��3^Z����`.��Z%�������6|�k��ʙ2���mㆣ8�TS�g�Ħbh��0h:���?�G$���SM�#4oA�*��<��-A(T2�ץ$~ϲP����=�:�\ [��X�Q'�{�̢鴎�q��,)���%���7ָ�{~_n�w�<#��L:�Z/A��O�����jy�0�y�T��w��~w)wC�t3D���@�1���+�����^{��c����F���W	�O��;� ���r%��8vO]�~J��w��w�	m��;�w��
J ظ7�;�fܽ�W�z{�ɝ�:�}lX��{ �y�����z�g��c	�w�`5���y��5��8��a<7�1M����`��'�Q;�����9S����W7�y����?v�U�t�k��(�h�f����ހ^)��K��.��8� �D�K6Ʃ������FX��S�XKu%���Ԣy!�/��Z��x�hb���(-M,:���jv���f���#�ŗ�fW�$�XO��L*�5����=[��+��1��8M �ԉ$Xgx�W�ʁ^ǅ��8������� �L�ZG�������ä��� 0y�K�^�TZRF�C׊�e11G1����#�����a;*�&~��4�*�⎞J9�[�*���j(�Wф�ys/��K���k!�FhY�7��.u�ɀ�G�T�C�բ�a���v��l'�����W���+ b�s0���nB%U��P@�Jv!L�΃��0�G�5eK��`"���T�S͟�+�Ѝ8��^��{?}J�->�/���^Xm(	^�l�3��l���uw!�?v�f�<�3����j{���\�@�׾a˖�p�H!i	�v)(�L(ka�v�X�V5�o�=?}%���Y\q��Dg�f�Z؅8�9ݵy��8c�b~{�H�*,nx���P��(�;�����gpu"l��q�f;i��+�Ĕ	(j�M��
��1�������������Y#�XE_6����%����F���?J���o�Q9a#0�ۙ�*k���ԅ��7iy�e߽{����1�^�;�w�K��>�=@ރ��琘{�����ۃ�����O��x��͌�4ʸ��O���QlTԽw��!�W����_�p�aڦR�桲q�y 1ٵH) �g�'@�M�7y7��c�ZKJƜ�1v� �MB�-���C��ཋ��4���g���`���3[����V\>��S2_hn�$]PYo_��5<�qVgw?��.��2��O��<���SdM0�0�-t�gO�M�浳���)�R	�z���y�� �2׸SĳVv3dƭ�%����M`�J��M=SK������&O� ��j���!�)p�+��Z%nW�d��s��H�.`�*��w�B0juC�W�
� �����]�����c���e����ܓC��{z�y?W�0.�yI0�?���9/��=���;N����@e���z����̈���{�L��n��YM�_�����y���?�M��6T��0ɘ�R�@��ڥ,+ Z}������O�Fں�ն���(%�@Y7�y�z�+ƃ���+�T��#��3RA�,Ca��4��B^Yg9��'�hr� X�LFc�aP��l����B��D�]$�n�F�d�i�%]�D�ɱ�� 5PnS4Pf:�n�����_���5�HcЮ���$��GSs��
Qn����F�&��|�+�r�-+�Y��4m��q�.ԩՀ�>]O?P9���&�8�^*!ţ7I�9B�@1�#��w����ZXD�bS:`��o�N�`����)�]�ı܋x9ey�-�Seh��h�P�Q�-9��I@O]1��T�����v�r�p��JV��D8qO��sNpNn�@���r]4%�H�f0d���Z�*��`5r|�.˼M�3m���,jm���h��}kl1.�s�M��W�a���O�1�>���i{�V��̢z[��.�`�M=�*¦����+���ޮ���'���1 vC��>~ۧ���ǔh�ví�%�~q�O�$��6���4s���+'t����oz��鑵��k[� �w�ﵳ�γgͥ l��X�mٸ;M-�'�� Qr��k�q�`#�_-Z��@L�0�C�]�jƀ|�B�O&ÈU���7^g�S"��~jG��t��p(��:���K
P�&�?�0�@ k�)����x���z���~�}�=���z���@�aC�_��Q��J�v�
���L7�쐍u�0,��'M���xO����(����Ɣ�)���E��2C��Yks�Xa���_yc���N�'���LXb$t�쯶?�����{���c���ÆO�o�O ��Xe[v���K���c=ns�OS��������yA-�w���[��al����ʜ���̘+�򐋾+��`4�b��y�~������d̡�DU /)�c.`:���^��8�oڶ�r�N��d����z޻�iՑ�k�(.1wb��_��--�ꑝ}Ů���Z�#��]��۟���`��` �χ�/��X��F�{_��R�ｃ�?(
�
�;� ��^=�wM��� FɱX����s3���P����t.n������=|ϫ��z}�X��]�u /���vHh�!9��zbѭȍ��]X{L&LE��U�x�Tf� �:s�Z<���/�5/���A[�0#��a��5�M�~!�~���(�[Yhm�X���2K#��9#����d�iCG��� 
&�$v�݈�e*�B�*�2������ГE�=��IHJ`�Xf�͜j�]��J�љ�Ȟ}�5<���
� ������Ll����d��H>M��.�3����;�����- Vt�++�)k).�	��v0�N P�4ұ��UB�X&�\J��`�����7� ��vD�CX(�$��j�S�[]_m����5j�Xv��@k:N�ڹ�8e+Qo3�a7������,��*�������;L��2n��O&j�� ��Q��~��c�z�NJMr=�H�]��G"s2�� �*�1G�-�S�:;3���x۹��k�;�"�s����\C���fΘ
(��_��tCn�yg�i����6���q�!�(��E��>u�
;��8�����=����a�l��B$�Qf%�ML.ݖ��Lt������0嗚�R⧆w3��zZ�{셗_�b�J���EH'���q�ph���t���Fٷ�z3�����0~{�\e7\w���X�(V2��/̢��1"3Wu��C5&Atv�,��h"g̜m'��b�R��K.\F4�t�ï~�XǍ�Ѧ���\qFl7� <�N��:0���I�w� TZ�%��(&�e�RTP�J������g#�*�E����3�9����T*	�t/VXcZWҕr��>. m]\�8�Ƒ�,<>��X8���³Fwyu61��#��s��U/��b{��s��a��ئG6`m1����he@���]��+�FL_bm<����A+��T���8����s�e~V�R-	#��v"���l���W� 9�
��A�=�=͘=��Y�fr�O�5��㻃�Cz�%�6k�[��o��[ ���ϸ4�I4�JF�N�J���|�Ԋ�-4'��Az?���T��[\�.n*�+;��3�E��^x���? �P'c[��` l���E>��� ;	@qo8��ț��{~��M ������\S-za��V?4�Ƣ��(ˡ�f����c��aK�<�1$%���<�>z�$�d[<ϡr(}X��}�z�W�����u��.L6߸�r���?�蘸b©���ė;~����(���*&�z R4w�ʗ���HI����at��ȹ�'Ѵ9]U<Ҟ�.{��Ģc��G��W�o˗.F�@nZu,A�̓S��} Lt�j�#_�e�a������L\�S�J�ݾ��yy���Qi��7�sra��,�3���%����tÕ�q4�r��ټmeL{��&����f:���͟6w�˧����+j+,-5`6��v�h� �ƌĬR�E,����e�B�n5��a�d�,bj�Wǔ� t��
 /�����Ґ�%C(l��::]Dv2��O��*wHw"o3�w�r�%�����k����ٰ{�t�~s�Y��q8�_o�7�>��[��h��q�y�dF���6a$^F�l���l��������f,8Ӿ����s���U/�f��u@�ؘT\�|���(�4b�l�c���E��.=�4N3����]�ځ�����ҟ�B��'���l���(5<���k�8a;�cj�m;q�����c���D~a]���!������p�4��]A�0�- ��*��Pl�B�}���x�eK��.�����(q�y�&���ɓ �y ���Bt�{~��Ș���ě�_*<����)6J���S҄�{�h��CW�@����T��9�<5�`�ґ��q
 G�M�%�R�6r `�e9C[�+�g�\4����:�@��7Lw%U�:4�bP��M`Ú��� �������x��;�=�tנ�7��C���3����Yӽ��<#�X���i�������9�1��=�آbˣ᧱����X5��c�	����:�e,۠���۱�I��؂o`�Yz���%lt?bo�܁q2FF���F��U6�U�5��As�@��V~��
O-h� ��A�����X����2�7�NV6� c�,�Z�:��[ ��c��������
�D�Z�`������);���Q�&- �O���r�l�`��:��7L�M�hc��L��(v�1b����M�+�n�:؇.X 	���;�ƎH�i��v�YK퓰�^�)��O�����O:A}^~�M�4Ů����������dS'���Xzv��"C�K�����D�d�|�6:BweVx��6s v����D��n��>֦^��Mlޱ��{������e��2~����s_;0��E�3LR� ��q�[�����5�F��e���.�]0�	1xII |��vβ�(�ô��s�>k�)�L;�DO���x�	|�rl6e4��a,ϽX8 �!��C�2�g�yx�W^}��0�s=Õ_���>U찗^zڐ�������/��s��y�Am����C�<fSR�ڴ�Y�R��o�����hU�E:7�Zi�|���tm\G)h��2�4��Xv��t��������ic�o�]�f�=`�����J'bjL��k��R��'.�Ƶ��ڭ0?��h��n��L�[�+������}�Q3��x��Gϱ���F��
[��:�p�15���,���)Sm���وѓ-lU�5����}k��h�=��+����&�ɸ\�l�՝s&��*���)��Xy���w�"g�b�7*�~����]��E���9g��ʱ�� �h��A3��<�b{"切����.�r�[��"���F^�l+�:�>��a4~HWf�=��'���\� 1���R�e	��Ev*����k�}��ם�?�}�G���a�?)h���H��:"���� ���6��4�>t��:�ơ6)0>� �6�J�@�U�K�x�� b�P$��־���,��?lϦ�6{��b�&��h<��F�ޟ,'B�H�H�ÛLJتu�R��+�V��i&�����h��4���jb��4�)��r#.����ݰ�I�x:6���ǣ!m�ٌߑ�Q�"QM�R:���=k���k�ҸK��E��`
�h�Q�i)���y���αal����2̙�J��Tl�e)L~n�ubo�����?�"�*����1?�	^���_K��N���<��������Sy��~w0���4n����sp���s5s����|��	��R}V%��a0��o��XO�^�ߓ0���@�� _��Qvc/�:b�^���ub���L�/"�Z����}�Š�E5�����J�[>z����?�y����do�'�M���s�r��3ΦT�BV�|���=d�GN K�x&�0:�����h�!i��M�����f��E�T�]��a���l��] 1�1Mm%{Q�CO�r��Q������췿��e�/����e��9A�LX3�ت�A趴�������؁��a�fb9r$��uN���~��\�lT�M�4ݥ	(�Fl��)+ح���͛��7ƹYoݲ��RzR���>�y�I6��)�p�.��q��7�K.u�� �g׾��҇�G���3��c�{�v;��e6z�PJ�%�/��;v��8U�դ��5�}�[Jc�ݒy���K��_`�-�`�����o���ƚ&�v�1�|��\�����O`�7���=JwW��r�-V�Pb���l\t�m�<����B�U���5ܖ~�#8�o���Z+!�|��%�BΜ1�����PdؾB�������^qA
`G���ɧ^�w,��}�1Jޭ�ԟi�a���Q*�:c�e$���#d�1�'c/�#�-GtJU!�v��Y	�t)|�����b��u�&�	H�ì��+�J'��*^j�Ei�:z"vF!2x�-�R(����7l��3��Kٷ��=�>e��Ȃ�� �2�,�Fd���K��Ei�_��S�mtޙ�9�@i��t�����+s�?�r"u� q���LqC`j垟A��_j�Ps�"�$��ˡ�&]�$�lņ	ȵ��qZe|���6�?=���$2�I���~g(����_���<�R��v�>�+?N@<�� @�X�g(zt�ͬ.�Z$�9��Q�&����^�C�47�p��=4���:f�x�Z�k<5�;$��FJ�1��H���(R ��Py�'���m�[� �VLl�*�bN�Őb�\�#z�.�W���X�(Ɇ��"a�"э��O@"�6i�Rv�{
t"���:�% Њ��s�-��?�2�3����z��@ Lc�?���N�R3$޸��}�=?3�_��zg�R�����1��`� �='�>��~��]�S9V�5�1k�>���>����W? ���ɋT�����8@(@Z&��F�C�L�:���{�lLe�d��i�++cG����OY&"�Q��>��Ch�6f���N���6m�\�0{�7���(� �UŪ��&J��K� ��ض�o�f�����r��S��*V(J��x9_+C�T=���ƏG��Z�+��o'�2c��"od'K�&�d>��s�I�g%v�	:N�ݗ��n�����\zo��$w����<�k,����0v�{ɋ;������,��6}�t,^�4��:�ͧ�|����(�6k� n!,��`�����Mi����E�n&@E�̙=�i3�Y%u�ʊRʓ'(���U�����y���lDߡp�z:g�ƺEI��YYT���ҶP��������� ��@�%�Uz��.��U�)�|1����Q�����-h�t��c�AL���X����/�P��>q��R�Ozܞz~��I��~n���|'�����^���~�.�N���v��n�Z����1N� ��(��:l58�˘�&@&�]�u�{o�Ua�;����o��5j��z�<�sq�ϳ�;���V�ʿ��Q��{�ɇcI$4L�ѓfQ�����E��!.c���lἅ����c���M�v�U��l�4��z0M��J��[�*�:+�$���_������?s��6{*6,��<[ETN6���%�6�WUcjc+�2ʼ}C�7*u��7����A';�==�%�����ϓIM;��8���2ҟ��x�8X�Cޢ�q���?�L"�T��K�⩃��-��8DP֯��q&LK��7�d�Ħ0�!�M�ز4,-xd���uM�q�m�s�f��a��|�[�a|�L��}�6�59�̞`����97I:QXюVX)v�����8��ٗfQ�s`H�J-T b	WB0Gå��%��.$ j���;�G��w;`�f||�mݼ�>q�Ul��O�Ժ�f(���ƻ���e1���x�ӲS����+n�i��k���h�*Ic;^y��K����y�T�Tc�<�\X����l�wس`���?��2���@��>��q����ܛ�����0�_��;����?�����I4��d���_vt�շh�K�������c�/�z�蝿@{�Y�J��x� ������L�} ������?��g��?�s`2��C3azo��>� �P�X|�W���؁/]���~2t���?^i�=���F;o�ٶt�gYA:�٧��u��q���u7�d��̴�&�Ux�9���/���"k��o��ӵ��ޱy�e&"'�1!1�&�����"Ŷ`�+@u�sOF�!���ݖw� �Q��s�4��q<�⣗�n�1�����t�Ա�{o`g}m}�qw���C	��kPh��ToKo���Vo�/���Eqwww�~k?�$'C���{����df�<��^{m�Դ
"RS[�.6�d4FmlT�#t}�*�鵷��o�D°pD���x��9�G�ZZ�~R]�h������IsR��l�{����{�Gk(��n�&JP1�2�]{�ho�^B����g�4-?��a�$0�Ʀ@Tѿ65�V��m�^6�_�lz���[}�0Q�$�&�T��|}4D�M�O%��V�� ��J��R7�JK���|6�kj�|�i"��e�>��� ��O�8�� }X,��=�	��qS�ٯ�v/�> ,�e^h�;�;!H��A�fR�U ��_[k��خM��b�K��-�b
HI�8�s�@�|σ�рy��|�l1M�����v���o���Y�هn���˕v߿�E+�P`��^ l� ~�h�k֌G�vS��u45���V�S����Kl�����o���W��[ �}�1jxE*�L@#5+�Mu�ui��f��څ��:�����۾]�l�"+E�I��l7�Jl�4qM�������`��6	^�b`ڄ5���h�|;Ձ^N�D�3��q�-�*��X~[�с�-K�4���U�ǻ�����E+*VUCK($� P$�k�N��r�Ym}2���$�P��J��cR]< �{�����-�H|�.{�g   IDAT�QO��c���lCFM��Ιc_XdM�j��L��"�U�0i��8T�C���?�&��Jkú�'�?��|u6Nl�%�O\S�^@��X����972
t��
���F
Z��"#�$�\��{�}e6=o�`���^��,���B����]��צȩv�.k\X��IᏎ1��* :�%�M�(��d�"~��m�9��� $@���@�r��v�SX�{��� �a���Q��-�\��AX��GK+z�*TY	��ּU�������6)�YSW��{���P���Ð0%5H���8�<}���f���y�4Rb�>t�]�kr>:�vؙ_��Wnq�M7ڰ#��=�����Ch}z��+.�Ysϴ��ⷊ�I�dPA�M;m�x�t�Y�٧Z����Sh<L_4 ��Ay������o�d_Y���U{lSi)��Q�]�<�����s�Mc�TZ5�TZ�����ge�ِ"6H������y$~0r�? 8'�� ~�^!�,Br,��㰡��%�0d�X���\� �mǬ�'ڪ�+i�����a:�l�&{�#���A0~�=�ē�_r?��n�[����|c�
{�UW�`�X�����l��j�,�kIGv�T���a+I�FQ�_��$��
��q8hR���S'���sʹ	u &����I���V�up�B�q��r�a��W��3�������a���X�����'�a�0�C��xEu�7d��}�iMUKJ��>}˭ �X�F��:��{��)�����X[P��g�e��г��w��k��K��{eSj ��뮽;
L�;m;եټf�RF����O�����\�;k������)�<��w��6f�>��g�Ʃ�e�nZg��Fͣ��!,���+hDEQB/��|��I)�d��W4h��sS{���J�sc�˽ُ�@)��g�a�Nc?��O���k�����ҋ+d��NA��~�"v	�b�"4�C#��<��%:xI8��8Q��Ө��L��"E64 �6�f �*e�,�jf���I����OZ���{�'�4����n�Rw&�*"X��߉�'	��0��U�[RU��Ҍ��-��PA����
G��.g���d�T�2�6o\n��d\|�|{���
 �.��):R���%�Uepu�~�:t`��`��v�*e�6AQ)��p�.P�3FZS,��Z`��dG<TL2���]=1I��Þ����"1Q�D X��FF��a�4��[M�밑ij��0�麠�[�6�cR�[��X21`
�e%��gy�:'������L;ꝏ�u�"٘�ώ���
XNk~��@F�q���k�vM��A�3��!����p�#�[ ��a��n��ﭮ�!��ٷ��.a=�@ �
���I!sOOm��7�OpIX�ǂ���6�v��x�T4�YqA��4}2��9l}vʌ��v�}��[�W�u{��N��2���=G�Z�� ���6۔�-;=˅
���e{�m���S6��7��B�9  ��ꞿ�o�����͗��"��X0b[ʬ���T��v�	�z#��tx28�My�e�.��z�������	G�T�!�a$;k�	����`Dڷ�X��2S_�H}ʡ�w�·q���Ǜ(�I=i�f��Z���^}�U4(ݰ�h�S�6���[��rRbM�igS�G:��VՏ���Ϙ3�/�6r 4%vμy�+��&���D	����Z��*�z�0�Q�ȸV�W��L�ao,]���ۄI���/b�b�h��O>IJ���}�R�j*�v;΄�7��9���� т��S��J�F����r2it�K t)���uI�}�T��ņ�&�'�6�����g7}�6}�[�������ZАe�U�klWS�vV$��/~�.=�$���K����|���"�`��)���`�q��z}F��I���^~�ٰ�	��l��<۳o)�&��
m�� q�ݪ��۶��k��ϱ�~޶èL�6F��^]��D����y�6{�Յt���^Sݤؕ2�V�*2uW���b\Ơm��b�d"�ˣ�� o��qrOw:ʤ�k�T�68e�z��
X"i.~��!D��0?²^|��
	wRR`lSR(< �xK&١���W#18+@�Q�������m�ԳU��rx�a�=P�=��%��"��@#�";�ݬ)۩$7f�M㞊��Ҽ�v��'��a �e�ޡ�#C���i����*)X�%�B����LpN���<î��|{S��zR�	�A?Q��� ��m�fkbC�k���N���*	v��+'v?%� (��.3fU?�06�d9����K���K�B(�[�k�AW?��-3�BR�Mh�N�3�f�H�,c�D׉v��Z� �O�vQ��9��Zۻ�G��u,)L����G~i3}��7�ԑ�����*F�pJ�M�;O�}�.H��#�#��#]�c9��^`#�_.������H �pl���H��Pp�#�Y�s�Z`�����۱���>�53aG�����9!bXl�|�0�Q�����N�|�V��[�ʋ/�K/���
{�_�y�G>�A�䭷��#�.B����o���j��:��8e�c����Ġ���cl4���������Y�79�h���+Z�������.�<��#تmK��f�šU�mM���$� �|��-�a�IA����Z78�f��)Cc�v�6s�T*���
Ԭ7���i��Т��½:�L�[�?r��hCǐLA��;�~�G�Ң���`]E���@��S@���<�x�����m��d��엱�&`���\���G����^��x1��q�O�cͤ�7l܂��� ������R�|6#T�W[3UK^_A:�P�)��ԑ��*��n�8��<H�(�	��F����  (� �)&.�R��jkҌ�,�N�0�s��U����q&=�&ؚ5+�~�Vo^k��y
ƫ9�v��T)�l�;�X���T����I��߻���,�Λa��1�6F��5��Ttrsmݎݶ�����N�/~2�b�6ZL=�j���^6������'8xݽ��~��;�0w�議��O�����'��$S<���س4�.GO4���R2���P@������L�o���-]�6R�zH������j� ���H>��׼�b?<��¼���mu�pb�ݜ{KK���>�p��Ii:�А> VR�oN��+<
"(�pD�TY:�T�r侫E��!!uP��<?˹]KKt��7���ˣg�2Ys�!<�cP�+�����ѼL����C��$RŐ�����hڶ	a�_Lϓ����#�'&wy��^��ƹ��E)�F�
t`��\m��dƬ�s�եk)>��N�e��!�����s�{ˤP��`N�.} �(�>i�T #]�l|H?����5N�S�#����uP�v��S6�~���p�u�y(كT@��eH	:Г�b��i�jX�B̋s���+���7�� ��[`�L'�Bz0��o�uM��]Vk���ąt�G�a7q�)��U�X�����Xa�f���D20GD���g�-��N��}�1���p��|��1]�@�p,�?���=��-�}m�iw�K��;Pc8�5���]��a����c
���M��M�J��JD��
p��y�{l�'��Ihs��Qe�WH׌6��Ff"��D_����T�t�p��(�)�&M�����_�9���;�T;c��J�Ĥ�k���E��jO.x�tfpiɝ6����{���!v��o���kX�&�!��gg�8�&My��|c��$�'?t��*Ȱ֚���26�1v�cO8HQ�ny3��w���!O��^; ��$�O踊���T��bS�8�+fC�ُ��`,+$�VZX���Ţ�r-3`��^H��^�~ҳlp�xQO�����Y�F���`&)�N��]�2�Ʉɒ3��M[�Dby	�U�P(;p`�d�\��-'Е��8��6zՅ8����@�ئ){�:�K����2$�^��j��9�{L`,�
4���Z�mD���7�^���Sh�hV��?�>,2б<��l�'o��&Ιiũy��{���7[tv.�I6���,kh��Uwؘ��l��x�u��3�������ʇ��j�������m�vb�i/�������=��m:Ǳ�|����?��m���>��a��N����݈��Pi�6��2(-!5��ؾ� =��ȢN�	;�`��Y��P��$���|��1��9o�M�2����0����d|��|ȠbSt�l��V��-��b��� r,.�w� ���H�Ҋ��|W���ͨ�͢Z�
�+=�����T:%��|�<�_�7]��jI'�i�k�O��*`�Cuk&^~��1Ǥ�9�����,]�:I��R�IE-��8�s=i�,�\�R�SRt�b�Qw
Kه�1�Tr�-}a�]uյ�-�lG����K(ϑ��տ
�4�;��j���j�x:x�~���bQN��R�Q5c�"�C��/ٕ�̓^o;�yu3.�jJx
�h�"��6)���]�1U���0���=���Ų��6d��D�jg$��
l�8.�3�`j��+'}e������|�f
o��
^���V�H��a��DVn,:9�&�xE�Fo������|�[ͫ�]��1}Ap�u?_{Q$0=���@��` b:F�u�g��d��f� �`D;���P�Mxobg��	ꁫ�f�ǹ�H��ߒZ��*-=�.:�t{ᥗ���T��ͩ�[n��,4��/N�K6��S�H�����.�RM����Z"�X�Q8Tg��|���H����y����;��sO��uZ�*��w�eӦ�u��B������f���|�B�h0�aE�H1����om��b�/|�vی���sN�0��=�VkA�I曃6�H���M=1�\��Vc���d	�/)G�,�-TY%�x���c���P�H�߄p?�jE����k� KD�!-��M-��&�'1,���][�KQ�6=�t�>�Bqq��G%�Od���d�K-vB��$VjA��"�x>;J���Y�z���E�ȵ��ʄ5O7ym���F/��E�\F6�>nJ]M�-���t𠡌����쳉�f�w~�S����~�f���y��v�Y����O�ʲ����w���U6o�\�ݳu�}������тi&L^vn,��� Z�$�S�oKi���RU�%�8��9v�sm��/�]���ƍdӦ�����&�{�_�4A�B��[[^mk�4f�xQ�K���E�T�f�&Ǡ/��������z�X��>ڈ�l*鏕���MpPV��l]e���lĐ��Ͼ�7X��ƒ&J���4h6i�0�����`^�[<Bw�@J2��s'ѷ5\��d�W��X+HD�!�Aw�W'*�<-��%܎�Sg �LA�52>��,Z��p�U%�(��07�3M  Ҍ��̹����'�+A��WJթB�|�)���KH�qIĻK�k'�=�b��3f�\`�X$ Q�+�����]s��hkU�d��L�+�R긃�0n�h�2��0�^|�I��YF�[N6����J�t��J��N!IF�]�2��J��Щ��������`'�52���X-u����ů��1�|l�A�>�zg��%��b��9��"��$��I�3S	��[0f]O�-�b�'Y~Z�I�o��sKf��zD������~ĪI��xM�a��=���H$9 �����0�9V0N-��'R��mҿ�M����nͨ���^�o�=�����1�^��@�y�ϊ|ޱ�����з:�H�80�|�.Є�Z7�d��v��'wT��tJkF�"M����DW�u��!zυ�������´Y�����Ź�Ӷ�u7�����bw�}�]y���Q��쪏|ؖ�A�f�ne���,��e��;�FS)X�FC�����*��'+ݻǮ��J�0~,�z���V�X�b�N���V�T�lX��ʶ�E�>�Hn���6�r�T�! ���6g�ɮcJ�miG������JD�5�����E��6����鰏X��9��x�F��2�^�VJ�3�3�cG�@CB,���t,<�Z���%����u���Nb7Ra�8mVr����>�B܆���,�U�&��/�!�J�*��ף��ˀ�ҽU�A�j�
&�(%��E�"{/�ҬI����p��{�C��~)����]l������e��>D��V�%rKROKh�<���c��W�~:���k&�[V�0[�a�}��߶��Q�}�����$�M@f����/��,�O���6��v�I�l�%'ں��ڦ�kI��h8� w�[���i��b�W�m�y��s��s����q>�6��vޙ�8|
S�gN�
i����m�Yg�Xҋ{0���Gj��?>{#�����'߰����@���i�^8�*w����̲�Ӧ�b|󪹏�g��&�!�mKV�"��=v�E�l��,{��{,���Ez���}lb2���f3�Ő
$�-�)
�녂C5��#�� Xr�Wcg%�&�����m�3b�, T�n��:%
G��
�Pi���eWZ$U!��(����LcK��`Rj�k&�z�8�s�����K�#�@�����#���o�q�m��zu_�B�/fv���.$�UENN>)���ڴz��>K��aCp2l�mީaU��P6ԫ���bze�#'}fkk���o�ݒ��Һ�s�j;��`���SRUd&RY�h���}L:��},VAu3�4sk:�����-��Av��e�F�*̛�,޲a�-*���mD,ލ�)U�5�ΕTd���t��H 킟��㝱wIV���06���W߆��ʆN��LՖ�*���l�e% Gҩ���0����qo&M����`C*,j�Ҫv�7w�����:�fh {6PS��!�=C驠:��"7t-���tO�k4�F�_	L�*���E2n����kh�9��x8&&�H���p
X�y'{��
��qD�����}h+]��|���{�sTD���!��_ۣ��G��z��m`*{���[��#�20_,_r�Gx7�}c2E��u�#%�R��DRS�l���N��Ͽo�]�]p�9�wz�q����,g�t��Go�vh�|�.���Y�s3��������?��K�ۮ�^ô�	9�μ�,7_�:�ضm�a��j����%���l��ݖ?8�V2��.q6�ݙ6���g�}2͑I[�f��W���ϴ��^�6��9.dI�Z
Q�c�?3�@;���&M�C~;/����)I}F����x��"�具��s}��?MfG�X�0��L���<�7������xD�������X�c��Q�W��Z���A���J�6c�|�����_�8U���q�Z���o~�+{_���� ��Ψ����@h��c�����f���f  I��Z3O#p?��s��ӈxl��y��l�X`W�G'�����{�ǆ�َ�\N����IŜR�iq��j�g�D$E��d�Ȗ�~���H�Eh�i_��G�iC����9��j�5[�Qa�gu���a5�a�������kq.��<Ͼ���ݻ9�1����_@�1��H�_�ט�� )g|���أ�1L�T	�� �%aP�/�G�O��:�A�_Z�aQ��!>>��K��U_��H�+���*�P^x�Me.�br�K?�3z��$8� �k9ޏ|���i���ОJ[�^�V�!'�E� �Y��z�h����=�e�������T9(u�3�8Ӹ���r������+R�O<�O�w�v��=��`m��Ft���AU�UR���I@r�A�껚�f�~U�	�9��c�|͜`9����m�hHK�Ռ���Wٸ�KKPzPb|BU�r�'`�GY �G��|���wͽk��J���L�G���#��!�B�W'Ou}$�@+-�Y	uH�@���:֔ԑ���ؐc]ߊQ	��c�A������g+�x�G7��ua@	��������f�i��򚣽�q�0�|8,��i~A�?64ʗ��+��F�_��;6��_N�$Br�/<�ʦ���7VP�]L��i���?I���X�o�p|.kΤO^���WlW5wa���d�9����(��_x��A���?�g7|�ZKE���i�����K�����[��w���B����B8�H����^%�y
�˷3�_@��D�{��a2
�}�\�t�]y�����:�Spj]�t���������%/B��A"Q�"�"�6���;�~��'�Ƹ���L����o��_���z����_��Tx���b 	��f�x���\�f�I�j]9�f�T��y��q��a�Vەl<���^�۷���l���ب\F�h��e��hꍦ��Լ"�=��k˱�h۟e��m�(�Ey6q�4�K�-�%@G�MD���q��S�,#���=y����_F�x6�K�Ϸ5�ϝ{�Y7,�X�T��Jßu����~���~���ND��\ �f��0f>�M��7Ta��R��G��a�IƷ-	����I[Q����=���B��Zaz��&�Έ-�4�"�F�K�S�K8��V�n�Gx}i������Gt�V�j=��0f�@C��<��(�P��x@�4��hk�S�v֓݀�<�V�@�1��tb���d���3t��B ���+85f����3v����C����i�ԃN��p� 6h+�Ă��0͚�G�CYȈU�Ϗc��o��]}�Y4&�l50���>��� `k�M�kL/EL�Ϥ � b���%�
K�(���J��=+%��^0s�Ktg��uU]|�փ���8d �s��U��AE�\�t7�ni�sP���7̘��v+|���ɯe�r4ْn�8*x�`z"?�g��	.��>2Fow>�X���>��ᑮ�����{u���o��Ϗ+�����c���~�q�����c���.@ݒdE��F�Hj���O�=f�,�����=��
�[�|��}��*X�r�,<��8��PY�d�������7���^yM��`*�_��n;����~����,(�_��~{�5֟��D��'��4}��>{������kI��. p���o`�d���'R��\���4Wi�(t2|�O��o��dRp��I� h@K��$G-�}7���}�C�����eZ�=����J�2�	,ڨTRt�tExc�*z/>a�q��$����i}K/�]{���gLg_Z��L[���^_�C�HK�۾z/c!߮��Xھ�t��٤�V��fS������	nzv"��F������R�B�k� �R`/���6`��4������w���SsM�=�t������}��ˬ2�쓦x����I���6�묗�)�"����g�ng�x�=����e7���0`�hhd? ��4���="���Q��=�bb4�j� �4e:b�Dq�A�/��2a@kvq���JOC[TM��*���S1+#�8�gcH���S~ajh���`<^V���"����#��ȍ�@R��0u��N����q��א*UW�X�d�oQv�ժjM��fO�� � �ZG%���/�1%�}GU�,aL�dĚ�XI�N*zٚU���3����#O�h)ţQ�R�H�HBV��i�F��۫�ۤ��[Є��?����6uH�E��3� ��n�￙�+;���Xs�l��MZ?�����H�5��.$��j�&P��.X�NR��򺃆mD�م�3�9���D�f�ӆ@�*�uM�}�Uf�b7�& ɘS�M��ms��
9޲2NL���Ia�X*Xf�9��� �͌߱������-=z������xm"h�5�B�w����T���:��#ƹ��d"��>D��nM>i;��bny�q?I�-"�/��l-a�Ek��Ĕ����u?��i�4o�����	���_����[���
g�]���o���2�S�����o��54�Iu�R�	v͖O8a������]e��[����'�ܮ�^I���Wڂ�_�{���2����͚3Qh������X<̘9�ٍŋ������@Pz�5QoQQ����-�A�R�^Z����\�Ua���x���K�`�J����_6Ӟ^��㟏�g��E{�k3|�1 �L
2Z�`�r�P5�H��$$�R�1Ap2�S��R`//|�.?�\���N�
�T����q_�o]�5���qd�p�פ&km����S;���O�r��I�
P�MaD�mv�S�Q��m�_��76�L�w�i�-����zᩧ��td4)�(����<� �g�ת�K锐����;*�ܵ�+��$t�=́����@L7Q��.���"U���]���=�P�?QG�$���0;3�5�)����A(�C24��Rm�$t�wgN��K��Ō1xԡ���v�pJ�su���5�̾�Z^���H�/ ��B�X������ F}'�;1r^�YF� ����*���>HC*]+�
���D?�g:�4Z����پ�����r��{���h_�	���%	�6���Z�w�tU"��F�T_޵܊w]MA˨���ɧ��W�:�Bhck�uDuya�@Re/� 6Ŏ%2'�a5Q�a�¹�?͆��F�"(�����=��2R���~/3Wu��S�r  ~+��h��[�87�=~��g9Obl"����*�E�O�E׻��{��0��� ر��k9��t���9�޽W٩��k`>�pyL��q�0��B��D�aA��Lk}��O�EG:�C��{��|�`W�ܿ����93줓&b��ͮ�䧈һ�i<�NWd�T��?󬹶�fҵXN�*LE8߂g
�LW��-���}[lOV��|�U��M��Z���
��S��`����g��){�����t*}&w�U����qQl�=��{,}Ȏ{qo�dq�=�𣤛v�$�U��J��[}����Pį�fyY�C����Bل@�6餓N�,�
���%�հ���]fg�3��y�äUF���2�̌�8a�H���0���(EQ���Yk�1�;���ç[c�.{�;�~�R;���mΉ�I�Uڎ��m-��n�"�4q�]z��l��1���e��R��fث%�.en����dC���^�d^z�v��3e��F:�{�����VP,��n�Q0�򇏶u����X7�7����Y�졿���� ����c`V��,����YX�6XU�Ţ�:D�.9�d�=���R��Hw�]�=M mFb��e.
cG:Q��H��UOz*��i��DPk��}-�Ę)��^vاR��ЍYnU���]����7�D�1�sz���^?�qIMK�K��d��^{ �Q�G��c�Ƭ����m���~�F�(����4]�V ��*$��`DL��c O�"M��rM��<�b��Ux����
�]�j�'43��Tѓ��+/��v�U�_b7����>u�YN��"#�'�_K�����|ҹ:�^� ���9���
�_�=�i���\��&g�V��T�Ko/}�X��)������P
��?u�z�rCe2C�&�+#20����)5���ۑ����F�~�s2c��ܿ �w!�vT�rL���yp8Vo�L9Qy���#�7�B�쁢��������/D���Kp���a^�b/����"�,Z�TV����>D�=D���^?�T*痾�q���h���Ǘ1T-������nƉ�Q|�}��<�Ew�	Sl7ƢI,���񟡭u�a��;��S�>^SlӺ8Ǐ���p<M�������`4H�'9w�m�_cQhD������&9�(Tm:`:09�jh��'����Ì̜5޾��IwTz�`�"u�6����ǿ�
x��îp�C}~�WM� z�
R�b ����ک��l�����}�4;u�9v�C�ۖ��NzR1�����/�8����Ӹ�[�$ �UI�GJ����6��oӧ�J���{z�j>V���`8E�m�]7�:�l����V�lШb�~�<۳c')����k�T��O�D��wW=�+4�Jn�,'`�~OEd'i���ظ;��9�o���O��Ko�]Hc��Q,Έ���W�R4`í��X`io�����^��FI2`E�I/��9d�ۦ��U�]� 5�$���^͛��R?��*m�ʋ��I��Xvv�WV�����7FFڪ
X�����A1��\_��T�T������`���K��V�\9��0_�B�����m:¤��� ��B�jkk��Q��U�Q�=��4dTz�Gb�paİ��Cm�Iԯ>���Q�O VQ}wU������fʚ�0p.´u����$ھ͝6�j*˭����Z��zabIG��S�m4-��0M�<�N�<ֺO�@��%���/��5�@�x�#OR̴�&�$S���J����#7�Q�&̖Z�/ȗ���U�|�#�,Ƃ�^����2��u^j֊vQ�Z@Kz[]���-F0�"*��X�xU��t�������0=�h��H���M:�Ǒ��ýopNon�30�y���n�����#��#��p�i �NGa��y�{d���-��a�JC+IP�T�����%��D=�֮�c�$��Z{J�7�M z�a���<3۞c��X�����U�/U6�+i̢���Xl/]N�<J�ыh����I�&����Q���_�W����Kϴ���bc?��}��k{,6kz1�������z��y�$Z���E����K��FO+ ���3��;E��%a�t�%��x/4a��!�hd�S�����7���t�w,�p�^�"��#�4n��xJ��L�	ZnO�	h�P�g���l'���mv�x�ŵ�o��w���y�FϾ�HSH�������sI�L��o��dط��eT�*{\L46h����l�������>q�E�ȸ�{�
�>r��X��bhh�c��V`�0�]�v��t�Y���]�?�RI7n��\9�n��W�e��P C ��8��[��clw"�N�Dm�{[{��|�|�h�٣w��J6��05MU�C���l���a^��U�v	�"�������"��{�"i���~4��Fis:�E�H�9 -�712��rsU� P��9�EW{�D��X.��W�t_Qh@㰨�^�L��ҍ�x���*shMVG��R�������n�xi<9ˢ�.7|Y@��G{D���RZi�����H�*���}���ꯚ�Q�@���@c>Ͷ�
�=�ذ� m�F�N�@k-�!���s~�D<���゘��^�M��Z�$�3�G��.�®��\���[4^�c�����˝0�:*�Yo��9�>���:�\�CR��A�������(,������8.a��0ۃ=�#q�Y�`����j��cJ�箽�l:>5����/`*Y�x���Y��;S1T��X;=O�@�s�-�:�
4~�Z��M2���gd����|m������M����*8	�uGKս�a���p�/L{�+2%	o�~�Ǒ�����7l���
_��}���s(��]���A�@6r���{M������}6|���N=��U�'|�#��K+��WT��n���+8��A��Y�-7�jB+E���B��ڭ;�sW�5&�Ў��	9֡�MU\	Q�Z�q �l�"��v�;8�P&��SR]i��wذa�Vpz�՝�G�3�F�r������%k @�mwc��遅�̲�,txQ��[��\�����HY�d��(�ƆK��i�d�k�sS�̧LcO?��Z+v�2����?��]y�, ��A���&�k����O�Ы�4��o9��JX���8_9����u��89y��4Ć���*�W�?1
��K*`N;�l�食��S������3����[��}8��%���!ND��.�/N��4�6lfIl�%E��������v;r����+�(P��a����1����h�m��n���/1Am�\��&Ξ�=4�l�d�T���}��-v�%��D�E'���f�UhO̴��\g;7���^X@/�������l�_n|�Mv��s�n�!)�]6}�(k�uV�~X���*6y�-򫊥����+{�-F*LU�2��Y�Hi���@���6�(�;�3D��]��a���]�#ҽ�}P�#�� k	���+�6	��{i�xPt6E?�i���M��A�L�=0�Uem0���G�W�C ���@��v:Z���pI*p)�J�Q��Bַ,z���А���W&AhuM5��1`�Fᬟ8ӺS�~6�a��@@���q}�[�$� J�D�逶��>[��%+�A��/���6n_[j���6�D���l�'|�F��\��>�Y��P'6�R�z�=�Zey�)rA}1�DTy�����&��4�Z+E�B��j���/�T+����/�)U�6R��N�U���i�����q��'c���:O�7e���؊�V;�����cU"׮í���?P����3v���#�0��X���E���o�`#��� ����h 5����z��y���h L�X���n\�/����Ђ��Yk�>�D��<����a�g�:f|��I����:��X�?/.5����-9o8�ze� 4��fʥ�0eLd��X,Q�|�eվ��"�l�u���;'&�j��u�����2Q[-}ǰ!Cю�c���X}�k���Hy=��"?�VG��+ ��_���.�VV�DzmƔ�^���Ro�ה[���4j�0��.��rۻo�G�aQ�X�l�7�)7�à%2�y�s�=yz$m9��
���H���!���26.�:�o�g)>F-����� �瞶��l��*Z��B�쬳O���>�|teh`���.��t�&��AWu�ݏY��aVV��U��PUVB�������[�A\�۸Lr���jj�P��=��'���0h=�(�ݞzi�-xu��*h<��#%�n%!��*�����|Ȧ��ȥp����1�.&����l��	����n��l�衴���b�����8ٯ�����n�R�~����]#�
�h7e�+�&E��p��í���ּ��:�Ŕe�����z ��EM}Nu�$�Vګ�M��3h�y�t��T!��	���)��yk*zH?�bR��ƣtXҚǀk�����G-ư��4��"��0��?�>�D�����(�J��\���+Cn�J��6 �BUG����dґ�vT����E���K���Cj�k'��f��^i@U��ڣ�1�5R��&�[֭Zf�//��C��fm�b�d�/ <{���4���m^��s�N�/�!�Ym���D׸ԺiC��x��h��r�Щ�kH�61>Wu�n��U74hp�͵O`�&�.I�	�O�]	�9UB�K�S����׷6��	�)L��J#�7c�D~�Fn�a�~$�(��#�ǁ�u���ؖ��#���@�xӆ���#����ȗ��<x��F�p�*����l��v4`v�jՈcx���}�E��H=b���m�B������Q�Z����8n�}� !r�XW��2��4s�d���7�u��(��+l<��!�⩛u'�+p�ƲcA� 3�(w��hcT���n��3�a������t���϶����-֚��h+3ʽ<k1@,���̪ь�t5Pу�E#�(Ki��J��"��� ��'?�����Sg����6�أ펿<f�'MDOt"�w{z&<�ߊN~����0p������DG;��ꝷ{���>Q�4��@ު���.ڀDX4$�ZK�+���z���^6�a��K�*ޞ{q=%�e���γ���捔����I0>�\�}d�9�m��yb(d�	����i�.��} `E�o0� ��Cp?���sg�WT�ȡ� ӊGL��y5�glF����+
��Ip��N�C3cMĄ~�VM}6���4M��"��~��[-����,	'��	���O��ٛI��r�)�ƧF�nĩ�l*0+V� ����� .)^A 6N�Y�p�� �۽�d�����Z�L�q+m{����+�#�K�+$ja%�X'R�Ib���JcJ�G5�nƌ9����	��#��8���b���T�-��G�}��=��*�@���y�ox�
J% �:g�nO��h{k�!���Jz�� �ƌ�{b����c�� �	R���}g)�6H^͇�S̡�6�w���2V,]Jp����\>:]�+�M3�xx��L�^tw\������F�sO�eK6��'`��	��;�~L)y���P��� �cC2��6*��6�L�&uMe�����@U,���_��@'�^~^��*u��}$;��(��Ϗ�<����;
Kv��x����}�{}��f#�j�;������?����9���7��p<s�pA$�v珞?0�Gc����.���	���N8�~�H0�]DZV���_��s	&�#�$��H����q��qP��[�XUGݔA�ť⸜i�q,tD��2��,:-Z@M�5�(}��q����p���4K�E��"�r��AŰ�t�޵>K�fI�Ť{�}��G����K�e3x�#�����������	�Ϩ� LO�x�Fi��m�"�\D���_md^���h��N�L�lzYzZ�(�;t�9H"o��(�X��wz����c�����H��?6�q��:�n	����^���F�HZ/!�����6c�d�3�${��E6~҉v�e�ڶ=�ĳ�q�g��r���ؾ=5p��e�a�w�bC�*eLm�6���S��N�X�<��**����C9��W��+l�^����f뤾�S2�:k�>���Z&�-������@��6b說�^@��3gZ-���N��w//V�ϡ��i��h��,��)N��/�+^� �/�>X$i�r������2O}�9�}�J+��T�GvJ	�&�L�UJ�7-�^��c�ӟ�^-�ޯ4�u�Yp,�]G;�=5q��Z�I?�
�
�h�
�t�9��@����������[#��	S�(!�J Bf���D練<h
���DP�DU�\�.���̤�v�G�C�J�gꅪ���4�c�Q��K�o+�Ve*(�:��B�UPP'@��^�@�j��C|	�w0N��}���}%�y�j�0jf������O=e5�M�g�h?���ĥ��\菦Z=Ն�-d.ёdc����*���X @�S�o��S�)1bJO��PS蒘L��%��J*���Ĵ"[Fe���d�(����������:u*qs��ڱ����힮.^	1S��4��k�����J����!� ��팡#�������c��ȹ}�����N��ca�����-Y��#9I�{$;9���pg��{+���7�@8��]k@,�F�$�Hx?��t�����U��\�x�諃dc;��c�h">E;���V�8���޲��&k�Wj)��Z&�\�z��,�TI����r�YbJ��V�F���ټj3m�FP#�
�kj�%��y ��� �n"^����M�;`(����M��g��oD��0jy�?��S!�r�j6�No���R44K���<��#��	h���Am��	pPZ��]%��(�9�y:G{ϣ1a�y����J}��|�3�7?��y˘U'��"*mO!j޴��R��4�����j1}������U�c��r��슋.�)|����*��?g�f^c��܂����ր�����쥅��Eﻀ���i�2�&��Y[i�}�W[K}��s�\���_=m{jJ	>��tZmĘ)h 1ʄ�2r�U����ĸ�e#�Ӊȼ���)� bŲln���������8����?�� H�+Km
�جUT��8�%�Td/�D�mo�̿ń�=1b�
H��'���G�]֊}�a�*-$�#FLc\�X��{���B ,:�_J"l�,����K.t�����QO��M��-����M�/�5�� �n���ή�}�u���^4��H�/���?̠Io$�]Y�;`�D��c�;��>u�at�z0�孥ު�������J@	���d0��2��^�O,�sR��
�b<Z,1���$��Zu t���C�K��R��T����)��8����U���f���P౅��Y�/���V؏�d�,���ް<�DLV��������ھ|ۏ����H�(��&舉f�E�ცRV�#!>���SO�^�w�1n�]Wp��ۦ^��s�6QcR@Z`t떭��m���,�=F���4��1]�@�'���w�lT��y��,-n�s"�u�B�ۅW��va��1%}��=�!r�@��C򁁇������q�:������}T|�Pf�?�?˩T?��x#�w�����W֙�Л��$GyO���������	ݻ������!��������?��40����+4�H�3|��o��.���g�%�`�A6G��Y��z'���x��/�E�Ů�ܩy'�@�J�a��Xx� d-P�1DQ9h6��Wa�FT�Z�`���.�Π��.l"(��q����9u����:��/�m�]���F����SDu�M��!P�YK3b�7��eˢB�('���iVA3��l�#�\I��
0���d�H;�EYUE��6��,"���ȟ�B��xUfiR� ���:4����k<0j8p�}n��.��^�/4���a`��C慊����b�&�������L����Y����"3~@��]0���=��0�YD���׆�+q��p}r��OZEȾ��FMHx����u"t=u�@Yh"�xI��� y$Ud�7�F&������i��	ʱ��2*vw��W��M��:�㾻���?�;�3���O��d��_���t�B;����^e��`��x�l��˖�C����ɛ-���>��������܋lɋ��~K�Ec��F�F�0���oS�s'��n�ژ*��c	<bT��8%�8;��ldqƳ���QTB��^^3f�X+��DO��WDs�zQ�\c��D������^�_���o,��]��(ln���gc�Q]Qc��F��ȯ)|=}3q����1���y�"�>�ߡH AN�'/*���Z��J�2��P�],n�b���P&�*�t�ڸ����Q��e/ 6]� ���f��R�	��]�E��R#�n��}3L� ],.�*��!�qj����n������[F����L�|Ԅ�c������Z��((�w�~'���.@��݉�t�����S�k��^���inQm�"�.�,�U�+���Uk��XnMfj�3�q���8��J�KJ���E� ����&� !����tQ4	_���Y��7�[���`wh����������+��87r��TgF%֑AI��Lo�������`u0�'�,毞�\�����ºe+��E��Ə󂯁�wP%4�Vj�e�=��-�G���c9X�ÀM���$��o�tm����/���RU����s���))�2Bc'<}Bk�Ww�o��oF*j!�Z��t�h+||��  @ �<B����!���J�6�`��1���oB�-��_�}�!A�Kd�ï����-������z?�>��v�jI���Dc;A������P`ޏ�`(������U]'t���{�8� l��|];�{�����a��ݻS����;Fed_O|LKl|,-]�q��Ρ��HҎ^��m�Q�h��$8
+�Z�QRn��6~�x��~��mcO�����v�E�l��3�?��	��F���Μm�9����U�ڇ(��l��4��pqgte�|�4$��2����Dɚ��J��̃<��JK6��`��}���1�V��6��;�>�7~�bOg�fj����C�93�y\�i��D��v����
 �;!�c6ѷ�J��T��t�0�<4��^�[?�=R�$�ka舐����HdshbcP/N5��f���G:�K*hE7!&#�G+��A����Y�J��:Hq��!U��e:[WK��ǛN6�J��T��!p� j��*++��L2�UJ.M�4RD�b$:�,�v��� @V�};����nRd]�
iz��@eϕ&G"_�6T9������ ����E^Q3o���	Q��<B.���F�������:Q�ۧ�j���i�^뾬�6m�k+�m$�����v�'��J��HU�mA�|��jg\t����"[������#�W��^�#[l0���?�]�@���؋��t�hȤtJ�3�弻,Y:픢�Ō;�O,+�KR�x4%��.=��*�
�����/���m�s6c�L��߁��(+�БyG	R�)|��M���iJ��aõ������w��ǍFs��֮Y�6/�5��#�*�scc�������.�z�����P�=��QO�;�Mp�7��������{�E���S\�MTҳ�k�~%���)�4��\�Ru��{E!�$''Յ��h5�'5-��Ѯ݇kC�> ��	��:�҇%��'5�
F��x���l��ZH�E%@L(�Ҡ�����`F���}�R(����"�5S&�ӗ��&D����ЂI��sVKf��e��0`4mgޤ ��R!A�LsW�a�=����ƞ맍H����v8���cN$��&?'�"��W��L����vL�W۝�?�K�u��������� �ΣU��.�����j#}�L����\K�1�?�acYk�	|�b)��Nؾ821�  �5��j��Nw��xH�c@4�=� 9^.��[��T�kM`��˙�t��`���(6F����*xIf)ݞ��YP�	����X�İ9VԽm�]~�$�aP� �q�o΁����ڰ�t�=�xפ	�vJ^e�{��w?ɀ-(XѺ��|jTy~Y &�����2��:25G%�é�� S*��̍0��gx�H�Gc ܨ^�V A�A�[ib��AV�{EFI�"|�j�.�]�7a^-͵�x�ٹ%�ć:5p�J��sC���>Ɯ^�,�*��T��N��{(�I!&�'��󵕎9����X�JP�1U뚃	�0��z�<�.\ͭ�94j�@�9�A����^�}E+�/G�"ܯ�_Xh�"<B�K����[� �k���Ӯ�����l����K���u��q3aZWz���Yd�'_�ܣ}d,�mÀ�������� �&��b��-6�8Ն���$5وFGJP��N4��s��j���h��o�g�����ɓ�A䜊��%3ښ���9�tH�|h����M7@1
}ZuC�UՕ������l���Z̔ᭃ��	��c�02|��R�e��X�ng7Ⱥ���x���h�������"*]LĪU4,G߳u�� L�����m���`�Ӥ��I��S���Ag�����ss�I�\����}�Xi�����g�ꢴ|�F7ler��������|��1�F"� \�z5�`HRY�ٰ.�x�OȗR�N�D��uU6n�X۸q#� ì
�#m��^{%z�����Os.�|Q�&x�5W9��A�W_}����lWQe:~�{�':���b6�4Y2�U���p^m,1vҜ��w|��`�(��!:��"�&�U���N+��� N�a��c���>E��Qd�����	'X9�D]l"=э����g���j�s_3rl���h���}ž�����'τqʷk����J_�?��N�2q����wS�M�2ϯ�Q�Qos睄�)|?��i7&������m�xZ5%�ꥥ^��lb�(�֮��l��},�tqHI���,�nI [J�o��"�o\g�\f3'��=贌�<6_���r_�bz��8�k�Psc�"�����A����*����``�o{HC�#��`�\�ګ6y
��\���Т)ۄt �6=TI��9�P1J�i��W�`�o`h)a�@̹Rn]�����<]�\�Ԕ��ϗSzL ��Y��@�@��xMs#�w��ߜ�Z=izEʳ���]�S�����>:	�O�+�)�,��$���]=lN����p�#�F��]���ׄ6N� �"}���#�q����XwZW1�\�ME֗F$Ҿi�ؑn�^��%���@��TQRI��M����6�m��R���B`��'��@*Q��[n�S�dw��@��'���l��J ��OH4��S��ڕ���,���Za�:�.lT���V�)�/\Z�0QNJ�9��5��cd�VA)[XX$Pծ�E���#`����!# }M���&�*$�tE�g¤�no��>����-?`y;)�7�q����̟�Xr��됟�ϾC+,�\m��0/����diӴ�&�[h	�P!�K#A���6e�;ga4�@��V�J�n�(��@��;��!���ao��5��-���Tp.�K ����vYy���y���B<8�&1�������80��H��1��je&����}����&�G4 >:4W}f�b�fr�/�QId��Tf�K�@6 ���:����`��f.YW{
��Fd���S��o�8� ���|N�ß)���8P
��0Q�'mJ�y3dZ�tn጑�Ujl��[@�Sc�5�O���g4/�H%��א��R�[��s��9;���|��q��`����ԣ�I3���#O4�g���A�H��%���NF(��L�O��w9�}'-��^l�-_���O�Lt�M0�
���[l��A	��=�Kk�¾�⤡9�"�d,�E�D�k� �d�>'gB��$PY	{����RK��Hee��r�4��Go��&[��%�9u,��<�����π��ǭ���,��f�|W[��H�n�XnsfO����<$)�m���9��o�Ge?k׮u�t
�w%�Vn� k"}�}�6���?�鍈i�l+W�X��RZ��&]�͛7���S(3σ�hC�K��WPP��R��T�\��G�g��QU`k����>��s-��CM UMԩSquGȽ}�v��*<���}�V�w�)�n0c�o��6e���i�\O:z�)D�v�=����v5�U�  �I,����y�%�.�#��R SE�G;���J�w���#F�ӛ�(l��hj  8vw�ǫ�qG����&�c4�|�Ü��ة#]g��+����k/�e��k��og^0�C�{�E�>c�qΟ�x���'{���ﶍ���>J�gM�h���m�����0�r�N^�g�Z���k�z�#�HR�f��biD's��:�m�����9R�[�fQ��<a��S]j˗��O�Y�H~־��/����-_����,�%�Ww�L�Jc�l�m�4��(o!C��|��t-����2N��z���$�T����o���Elꥰc�,"�ؽk7폰�����M�� P��7-�}�����IA��N�i�a̰	�oBn�D�bs�K(�q��?1l�ꠠcQ*Q�oO2 W���VD��M�SzV3���}�u���ȼS����#�4h�P�o5����@���.�L��4{ٜS�b��Lz��1��9[�f
9� ^$Hi3����B��C����׮�O|�cv�����=[-�u`���6iJ�͟6��r��0�c-���u�a�jW\r�M=�Ϡ�\E����K0�}@i�hw���*�EW�XKH�F������yoJT�%a�K�{tw
�k�%�䐞���n����Ѱ�i?��a��B��65��$L�[L`"l��UiVUm&s]�&��欢��E�s��t�b���z,�&F�~�Ҙ̀5�u��ugڴ5��l)2���zo�1���˓gB5�K�_�E �k�c��y�I1b��7����s!����Zbj�tp�9D�i{@m�3���8�Pz�Y!��K���*�� ��C F=f�1n⭧8o��u������3�<�K�䪖@Z)(�	�)]�.2H;����EJ��9T� 	&&˩��kMʳN|�`��)�Ij��K���9K��b���&\@�c�����G���������p/E�.����)䠪W���s��AR�S`ʪT(2 ����쉈H�;:��2�27fdd�>$%mOww_Y�#:� L���7�ƨ�h�&�yS��jрKn�����D�
w���b�bl ��MD*���V9-"@����ɸ��N���C��� |r�cJ`A���.�Ӧ����RV�N@a|z�Ԩ ��<���Rn. a԰�V�c�]u�%TjvX9&����5�eC����B�(ǚ����ů�b���5�ȭ��� U��X��&���4�X�!�>)�SRR�0��� \�E &,���裏������IIp�����4���1t��ˑ���?��l��6�a6|�P[æ_U�@�k�/ф0&L�a%�+𓽇��H��m
����=�>h��-��9t�0X�uΊ)�Q��ꕩ���s�%�+��55�(�ʧŤ�-@��m[=��τ��3����C�YJ�x��;�5o��nYJ�6���Kl"e�ǷR���M6�)S�o(�Ӹ�F�)1O9&��o��FP٘Oˡ�{�ܼu��|k�@`Y�XT�k� �q����g��ȴ*�B�'d`Ex�0�N9u�{��5�N�5�&�ɣ���"�;m�x+��G��!3`1L�o|��Ц��9�Q�{��A�V��rlK��<R��iG3��B�H�� @�O˳r6���T��6�8�����/��ʿk���~MSө���EU��-�.�a�@��T��@�V�NXYY*��+l2 ~��[������9�l�����k�ЂE<�N�WhE�J
$��2^ *��+����Z��t����85"M��^��H���<kD	@R` M��i;���;�L)��,"�Ԕ�)�a����T�8��ɌE��H=J��Ȧ��,-��V�Xt��6;�
�K&u�=��M�S8�6'I�6�>���w�j�;����Ie��i��>q��k��@T:�b�DZ��`u��RҎ���7�߾��?�":6�0u�����b����g>�Q�W��F�h;�I:�*_(�2 =�H}���^�N�y��>�o/kcB�Oz�򣓳�p���,N
�D�@4�	0w��p?� �Q=T�g�2���[��:H�Z>�4:�4����֢kD��ƵK ʰ�c�t�k}��2�e��6��������:)E�Z�{h򮘩�y䛯�C�dj�
���X�p�`XH�/��
y�µ�����I�.	��
R�ٮ#R�]�W1К�x�a� b���H�(�`#dr�B|��u��z��tNa}�@��Jo�����5[��:'1�\q%/>g��4!��p��h���8;�Gp�Ih5��u��uʮmE��^~��Q3��m����9���y;�g���|�x�v������yI��E�	���#�<?�`S�!�ҀZ���⻴�����V�W���ա�v��R������"�@���^ T:F��g;�4Pѻ���������RK�R�c㥋8��A��@-��Š�p�dt�L�h~�e"&00�� b�)z�iC;��HI�"R���lM���}܆���)�]�e�5V,��A���-���i'ΜkiL��
��'R�?��e4R����䗡c,;`�Y�+��*&�,D��]�RB�%���jo �S�n#�3m��8��f�D�C�f۶�h�r���T�2� ����&�M�
	b���@>hp>z��P�v��no�����E�cɒ%�<i`<���s�xi��n�����;߲ */��RPA����e�d�Cl<n�hۏI���cp�.���j�|R�7�t���5`{6oD�,'�x��6��k��O�5[����\�1��$N��f�M�ï�F���XGZ")���V<���q���]�q��Lhoڲ���6}�tg9�`�br6R���i��r}%�^ ���[|�nشɵu-Dﺎ�$��H�[�� ��1�q��b���lҴ)V���i���j-V�k�y�8'�W�]\��V�V�dk���.��^~��ƍ� ==7�f�
@נ��Ċ�D��J��	��g-ۼ��̙�q�ۋ��[1����N�!�7�(�f�)��i4���à8S�m<Q�d�����Q�Y��oc��hG$�}Jt��/i����s�2�V��o��)ӛ}��-7��@XB�ƃ2�C��¶Z���:�����Ν;l�Z�
h^>�Mv�4���ZNv��u�ky�Jjɀ��"EpO��b��DH{�i�(;����E0"��Y�(U�롍�M�pK�J`�ʽ�b3VZ2Z�q�Q@�(�L���F5 ;�TP긃,�ҕ]�d"*����w��� %�[�h^���.�� n�9`t��^\P[�h��K��CZ�j�1{%�����t�ѭ�k9Ii�����`��+��z����O٧n�&�/[��1VZU��ʦK�_��6x�<�Fyj�g�k.���:�$
���M-@.��:�:��9�g<t4�1���h�I�^�~�3��T�7c���1q�
H3GS�%9A"K:�(�����m��ִ�^���.�}��!����z���z/~}�h�Yˆ,	�+�kf,��
Sp_�.)�Zm�
XŔ��+��U� D���J�	�EU���qTĩ�B�*��� ����MR�~�n�$m��>\���Y�B��|���=5�&��=�+"@)���g�B� .��x���o�7j�ο��GJ��;�+v�ŘS��.1T����d�.��`Gd��Ζ������F��D��o[��{JK,�?i��1�d�R@,˜Ǥ�h
9�t��M��6��宏ɲބ��Ŗ��k'�`��K�#���m=�$��q_ `d|yA�C�*'�T#�4�� ~,f~�������_زG�J�^���}jb�,�����xF����+a�i���Z���A�>Cŝ1��ZńE�p(��͒��C+&EKpǤ�b��U�^R[˗���[�RRW���'h�`]��TD�%�r�݈AC����fNb�Vl�4�]�:���!��`��L?�<���K&��baI�	�Z���iC.:����'�G`o@U�����?����ɧ���Z�R�T%���҉�D�7�S�C$�  �Bg��Q�S��A�O+��Z4�Q�!L��哀EL"z��2��r,�0`�1�ٻ�N�{*7ҋk׹1�&S<��𥗸n	6u�t���>F->Z[w�f��"��JZ=�Ê@�xE
�����e���֬Y�����l�5��a�4�t|z�U�Ғ�W�qVD�6l��mv´	>�_\����\��<���j<��F*�TŦ�z����֎�ȫi,̟X��+V9@H�uQR��uҚ)
U$�+��J�õ���1�|j���@"�����[?e'̜NO���g�'R�7ilZ0򰱈%-�/B/����������B���u�4�Bdy1��3Q=���WP�Ct��vֶ���H�
q1�Kz.Q%�=�P�V��
��m��a���M�ۉ�N��]{�tw)�X-��d���b�ң��)`�����f_��W���c۶c�E� +P��)&��C5Ul���6=�٨�NcQ���A�iq��v3�7�ܹ';xڷ�6_���g<�h��ڐ�)�R���� ��`�L����܃)��*T�����2�0 �Y��D�[�).��sl�dP�q��y�c�
�t	Z���� _�q4��XF��%�M�h�\/��V�lwp�U���<�����X�]_�Y�6wUk��.��!���(�z�Aiζ�����b�U�4�듾H6%^�d%0Iq�W_�}���|�W��]X�4���L�i&���%��	�$�H��6@%�����\Z�绿�޿�Q�ʙ��(�NH��q��t��p����g��"�S�E
� �w����ހ�-6;�l@f`)5�:IWq����QLk0z��������O|���8|v�+V�t�k��Gy�j�9���[_��/ߋQdM"�$�_jo�ױaz�[������o�B���|��*��r�ݕ��H�(�_R���b�'�/U`�#mb ��K�k��Ұ�H�#(������4>����ɒ;'�z��*�n��(����3>��A{��l�s6�%�����Ӧ�����]�L#��������|ZY��t��k(���Ѝ� ��.�Q{���@��1F'���d~�W�A��@O^p�Y{��v\UX���Ŵ���f��`����q]٧����ϊ-/�lN����o�J�E�,adj���i�h_��5�$8ė+o�����w	�4ƺ�N��Y�>�8t�?�6�F��
+�GO]�z��'� ��8-=soSE.��{7Ѭ0al��T�#d�.J;7��ʺU�%PJ߇K2 ��J�G����]w��ֿ<��B���h
������^�����+.������o�����:q~]�^�1�tdz��Q�`F)����-��s:-P��㋭�tc��pT.����|�͝5����~���-C&�,}P�0*g�>��4�#�zza�a�	ۉZQ�6�(����W�_]>����R}�^���I'�d{I=i�J&ZVl�	���R�s5���z��;���RњILO7��6�t�SGՖ"3E�|�V+K�*�W6
C�9(��Z،fҸ*�v�F"�"��<�12�D+Z�U��^�d���o��JJ���)���|��~N�ZKW���R�Y��IS�\��Y?�f�E���%˜mS6^���S�/����T�P�gϞs"u7Ql)�,�[^pb<j8�^J�C�1�f*ᾨsU�)e\^�Ϯ��b;u�8"�(�/k��� ��MYlUm��?YX�ԓ��l��� �� ��*a6��H�����V��YX���H[� ���(������j��6�М"�Ÿ?��8�gX~:&��Zz����-)+�r�Zt-:�RS�iϕe�?C+��6��N���5�I�9��}o_c�����v�m_������i�:
XF3н�������X Li�p�.��ھhAk�E��{�|�J��c滛�����*�TJ��V���������W��b��-`�
�5��F��-[��&r {��� ZKyd"��E+��|`����� �.&��ϖ�Y�(1 �����C.�TiSѧB�l1����e֬��چMYU�"P�f���j5��|��}{+�_� � ��Gض�_�}90�
	��e?\A:�D�g-��Z�櫪��BAs�71<��n���V����������% �OX�um}�bݣy;�����6����2�t<,�
��:�n�+)'����ta��צ��B�%A������0�!ϐ�Ǿ�*lc̆#w�e<�R��Kv$��ǦQ@e�Q��߀��D���z��T���`j�V.���Z!R�Ax�%��4l���FO%�����sv�Y�����Zhْz����|���F�
X��O5�"$~�	��$M�);m�W�Y�KÀa㦱�%E��,\�
G; �=�l9�e��؋u���������*�W�i'�T!J��O2*����+���f�
�z�~bx�T���x�P�
E�%vO�땍���m��C"���[�#�+\�(��]{���cq���hd��inAT߃>Z��ߋ�cP�b����&M�ig���eo`���3�$�N� CQȞ�Z�Y�")Q�6}FkGOe|R�v�\��74W�g�ޛLu/��tD��F�E�=2�e��l��ȭ�{KI}�ѝJ�+�2�c��r��h�����u��5%��
��v>���6�������-��8h��%j�D�.�ckc7����ɵkH��Q	��e�# @�I�dChk+����9�Z��E�OFk��]��F�w-����H�H�����L���и�)l"�+l���@��xu�����j u��Qt�L� �H�H~�0��t9F[7�55��zimzq�Nf��PB�_�9U�$����iC�M��<���sJ#v6����`�r�RI�/fI�Z� �6�~��,f�m�b��$������&i��Ih��pߩ�&n%JU���mA���	��x�T.%-Q듮 3l�p�oܰɡ}"�HIhB�n��/�f��>}�o�Z�%X�q�2R�S������d�yV����j�ZlȠ���*#��6e~BK��hOHm����L�[n�ɦ�vL���A��g'_��_���7y�$۶u�3���b�Ӣ*�;�7h��1���I�p=�G�u{`�
m�AV��e7~�S���~d��FM&�k��x�3cV��icO�亴�hZ� D�Zb��ͦ���T���OJZ1��V���;6�≅6�.u�	V�i�U��Ђ$�3��smb�6v@�,�6��l%�C;۽�ܗ��C��Alv[W�� �ẗc��า$�GqV^Â���Wo����W�5����b �ytw(�ڍ���k�EZ)6cI1C)--@��Mb����� ���,\it���7����"�еND�k�$�wO�g�D�b"Hu��R�C1�l#Q%��X��[�QF��5g�Q�9�#������;���619�+){E���� PrP�,�����j(�!��8Ǩ�%�)�'u�U�b�|Li����@A���б�����U)�P�B����/�B٭�l��r����Q�7�������E��Qɚ������>k���s_���u��t��.'��@�
������u�q���^�{�� ��^�W�+�λ� ��<�wm��D�GƓl^��NJ]鳓�@�[Fu���U��F2p�@f��56���М3�4�q6��J�F�s�v}�v��"��@���z��5dǞj;�̋	���ŋ{b3mriIӳ�-���YUK�#��x�󙪺�ԟ�6�fq�%hWN���_U��y���[�0�$�W�]Hs�����Ja.ɮ���W|�����/�E�n��<� ��/PGz�M�̻V X'd/��;��Ap�`���2�גc(u�xT���oUŽ��S��o�Xzi�I1�Rh�t,҈>1rxu*x�2*�p���]C��@$�L:D���{��d����sݬmQd���g�Ѻ~��A2M���!م2���I[N�v���ϳ�{֪�4��ᭌ�*��U�r-b=`z�ؤ�Ҩ��_�F��q�̆s��\=��i�c�h�R�/,@P򎰑)�'������J�ć�]ơ�;��dą��\N���oT� ��?bTT3 ���������}s�b3�*�a��Ќ��A�F��Fڊ�u3iEj�4swW�"�N�9�]����|1�\\����R��w�2�ո� �����7�$��:c-;��$�z�d��]����D�j�(�Q���3}F����N����Ι�|!�`�9���l�T�1p�7H������5$��E��w"�	�0���/9-��6���@á�N)F�R�>��XHߡ�T��ڼ��MSbBE�,:���,ۼi��Rq�"�����i�s��T�+4�N�qY��!P#͆�N�e�fC�y\(i�$�ׂ!CL���z��W|�)=(�����^~�e�G������/<O��P{}�
�ݡ<���|�Z++�q�Xh:���癧^t���"Rm�ee����dff�5� �v�Mh�dT07��&W����>���� 2@1|A�q�?��3�ĝ�>h��:��.���h�G���5��`ڛ�7��a?v��i�ڔl-:���Wd�-���GJZU;�+�,����LD���*�`3`�%��&��3}�U$��XV��ӢU��x�ǩ'����g��c[K�� �1y�֭|�+�%8�e�o���Wǵ'b�Y���4*����0�F��w��~������E���?�M+7P̂6�ZJQ�6r�[1 �Y�Q Hc��_��y�m�EQ7�#�
`��^x���s���T��L�>���N�w�qj�tb	��F��(� �Ãl�^��A�*�[�̕
Rp�8�#|�9Ұ�4�v����=b�e;!�&s]��;�a|H�y(NA�d.b�Hȭ�t?�4<ڠ�l�r�� E�V�u�:�©�0���-�:���U�KG�=J��.��?`��O��k��2��Y+i�@c���~��ҫ�c�~��~�Cx�ͱ&�������eL����2��b��8�����V�-b�h���ZNA��={��m0d"8���v��IE���,��ܢ�h��`��Ж�ܲ	rF���R��`�N9;S<���~���)cn�kkm��z���m��|��}0��lU�i)�zN'�n�����{��c�àe�O��^ye	��:@)���3*FI���"� �x���:�9�$�[etT�#̥�ګ�*�*���I��AZ��O2��6,5�)(�?댉ؾ�VK�FE�/��ú���]Z�6&���BtDp\V��S ��އ�A�h��+�w9#�ú����Ks@�A�]���i1�x�q���熛h+��<�{2��jƠo�j?��s<�>��yF��P&VZ6^��>�^y�WC�;���寒pp݆�9Ib��5�3N�,�?�Y�G���WJ��,�ݺ�n"��[�0{`��}�J�uiѥ(ӸF@��L`j)�t��Gq*
���X�9�y�GG�r>d��ZLg��.�T���,���4�4�uZ��)]��s�ɰT��'$Ǘ%�&��������_�e�A�.z,�iҍ��*�Ey���x��j}/�(Z���,�K�Q! �O=дj��.<�
���E�&@y&2��xb-U^�RM�w?[?H��P�#L��H���Ƣ�;w��K�mb�N�v�I�VcZ�$�,��ap*��Y�ĝ0V}�,[p��B@Z��h�	@����$3���	@���,��� u�{?��!&�tZ]6l��W�z1��
|I/&p#�����HmA�J���D�߯EfAQ���,�nB�*�X&U�����DTpYE��x2Մ-'��d�.@^K�N��m;��(��*"���ޕ��xVmYT��qXFk1E���[`<pt����h�aѱI��Pæ !�6KM�D��K�N��� q�!������-��V�m>n:���0���J�b�sC^u����(VkX�q�ؐ�짿��=��cvߣۇn�����GXDc�uVP���&}�Py��oاt�S�V�<	*����H5���5��Z*lJlo�5�w��BҊilZuT����'���-�$�=��d��O���x�Ŷզ����/o���gv���fO�yS�Z�g��[����m�9���(/��~�vgd����i'���C�gF���*�~��O~f����m��f���m��X*cnP6,2�X��]d�����WZUo���I�U4(�j�aXYlu�5q�d^J_�Reۍ�r~y%4W���z`G�f�'O-��\�F���;���4�z��Hqj�h,��Q�"R�� ƽς�A�T�A:�y��Qx��.��ߋN��4�h��`a����XWA�*�:Cg����+H]2󑿍'
񅰗�x�CG����J�Xx)_l���%��� }��`���6,��W��M���l�gZY��x؀i��j�����@�5a�-�*G�H��k+�_� ព��!��X����Mf^gR���b���%'3����1Po%���SgF
�G�K�h�֩�][���z־�<�����fv�w<��k����d�l�g��r���e�JME+%��Z�gAV�ղ6�k��T] n��\:/�:� ��iRX �SU�Թ�[��Y�'-���h@�d$1���8������Gk|s�nZ����zc.�3^Ǐ�iyx�i��a_������}��
駱Q�������z�x��DCR�cj"�q@��A( ����R�d2�	�w����q����|"�%I��k�~:(6��YΈ�Pъ���!h����*��r��%�T�ᠵ�֮^e����g���:���⩭�>BK+F������XS,������P��!ڰi`Lu�:eJ t�l�z	�Q}�,�ih�UO���z?��ǃ�Hҡ��ӄ�r��r%�,�� �zƒ�
�7/{�/�op��N��X�����ީ���(N��zH���f�Pi�sC�`.J�,���R�K2�����DۼW�y�}R�Y*�e��I�]GTJ��xX��|Mժ&|�hג�V (�^Z������,��ȯ\Fp�������2�:D�ݤA*�vYQ���^�/*=.�3|��j�j	ᱯ�`�9r&��6"����6m�4�G�M�z�I�����_O2v��l�*�� ^�~H�&� �6C�kІ]~��{	作p��%i�/&��e�W����)Il.Z��� %$
`�$�s��/?(�7�3�ח5�4'*U�uh'�U�͌���Y�Ka��_�Xج3����k�	`����_��y�>��>,���S�64��x��]6 ��:�Z��I,��R]��gT������e��)-�i(�xRR�����B{_���{�筋
�h���ɅhNhM�q� (���b|���m��Cz:�B��-=�BN�M�+�>�?����!�TUVZ�W��Y�v�I�y{�͎���>f��xp��n����a;q�o�f�������){a�#ة�,p�Q���oɦ�Yv�wص7]n���wm�J<�m9���g�m6"���9"����?�~o����O�ǧ�?���k73�k��i��#u�-ס��^�����F(�b�Y�xZN�JCʃN)��qJ1��wI�>R����2`\S]�sw���T?큡X�<�b'�0͋M�Rh�T�|Ȕ�����z�O�	j��61��ISʈ��M���l<��QU�]��m�ˆ�k/������;�
@X���{�WpM��Hɢ��A�V'�G�2;}�\[Ct�Ňo��]��+죟��=tCmls�0���fћ3�T�x֌^�d��l�jk�HE�i����O1���v��^�B��r�6k,�m�ʹ4�M3\��.vB�72���`�IeU�sO)���Ng,֣�LJ�c��1��l�0XY�\UA���!���%�߳���!M��b}Օ�L"p��a���X�̫(�
�����HF~�����e}�4c`���CX~�^�
�$����!ON���F���x
X N�7�sAZB������e���'5�/e����d֛�n�C�M"A��wz��&K�y6�5[ư����Y��خ�{Akz��9��:V���ێ ��NS�" ϙ��H�1BV�;���J(8л�*઺U�K��=�>%VP;�������險�ӝ�C}\�6�s��J���Q�<�ԇw(�tg�V�G�����;T���R�MF�u�5%O"X�@T_FZzGQ~�!ɉ���:�ƣ���/[�KB[LpM���mB�K����q�0��9w�z�i���5�JIJT�k0Q��:�g-)~N�b���H��"S7}$�2yeR6J�����0.�� [	�N' Ս��}T�JoSҽ�(��ІU��o��&Z�}��і�U�H�9|�4���'�A���?�M �ʤUI&��l� �u��M,�F�I��<�d�!�UUڌ����a�Уi3�F�p�j�k�8��]��Y+̛/:8	h����XhDK��*0='��&��w�8�ɯ3�P�2N��a`Ii<�z�!�q���p~�i�����q�%��%R�k���2����+i�vr�h�"Q3�I� ��D��5����x�5,�܇"�Js4��9���e��9='�T�&���g�wǪc�@^�L~M��p��H]�����J����x�tn�M�:��E�p^\Ht��E=x��ܵ���>^:���.x�@���Z���x*�vYvl�]��6S�Dt�?ݖ��f_�ޟX;YX�3Zmީ#-	}�ƭ��('G�"vR���� �ո��@�k��G�&k�1��ظa�6yt�-~�5{�T����v
��ɀʆ�h�^�|�} ���j�6�i��&�e��ί�_m�������@l+N>������=ӿ�~��G� �S���j�c�.7�-**v[���"���a=��äv�s�.
�T�H�F���D�b-w��n�s��5����̦�@i�t�%J2�\�4���B��A�!�x�i1_O\7F��$yQ���+���]hc���I���ؖǖ
�}��3��� �{ ��!v�Ou{g�Ef�8�a�1����M��׿�>��������{�;����o����x
�Q	@�#�?/�$��T/J�� �&�Mr�ub#��u��.&9�ăw�ˏ��"X�!{��Ǣc�t���]Z7kR�r�n�7�	�����D�q�r�C��dPͭ	��	Y��b���N��|��O��|�Qs�V�]9�/� J��.~.^�,�*;���*����U0�}������F�R����bu�'�4�`�Z{�׈�����sɈ 6z��׫�v'k_?��Y����W�x��z qs��5-Vkö]�����M*2�0��2.��})u��L�YH��
Q~_���0�r: H��T��i�7��&��b SҠ�捘-���K@��9A0 ���p;]����u�zn�9��(�z#����P��L��E��>2A%X&)�?����|�س�Y�4Uo��v�ȶ3�{������c��>�]z$zuDe�K�y<os� L� ;y7�U����t�z�Z+���!�7hA_,Z@6�c�b�`��
`
��&玽8Z�_ES�K�E���/Ħ��	���E���`P4R���kc��KZ.�D��$�幤%$(lF/їD��ED�T��%-T�\f�*W��X��H/ ��Z�bi��K)QԌŌ�t���H�AE/�1
ݿw��)��`���ٳa*j}c ���49�}��iJ��R�� ��I�y��|�B>(ǰ )hQZ@��T5YG��6��A�i��]��&'n�(��N�;t*Q���������1 ����lXt��*���U�U��w_���,��OԲ��*헁k'�TR�-ܗ�Li�Tt ��@� ��9�JU�H J唳`A�7i�`��|����	w��� ��lO�c u0��%�m&�F����j-�~�˻`:��K_���?¾��o�k�͡C�-7^��7���'I��?r����S,�q��xZ��Vl>�e�my�I+:�~���l,��t��(���_�;����%L��~�Y,N4=fl��%7n�h[���s�/�]*�~���BL��c��iT��и{�]J;�o�V�T���������Y�,Y���O��o�d�������?���N#�B�W�����A��A����*��$v*b�"��V�8}�"X�j��Z�2���/b;r��<��F�TՍ��N��ZO��D]�m�����*ߙ��q��LNu,�\�;Ҥ9�E�N`\�0!��VX��REn
�7,���RD��N ��9�7�K�+�ߵ=���@�<�\���ab%�u�����_s�����͟��ǟ�۾�m�����	
d J8�	��f"`^5`��z�t8���[^�q]�Ku��%v�I�?��U�������%%�T��(�I�2�y���L�6g*(�)G(�]0m�&�K)�*�q��F[��[LNՄ�-��ћb�f��y����zE��=����<"�M<�^x�i��d`���j&��۰q�P�.�a�k\<��y�`���
_]���AH�4y/F���0	��A�)����N��LB�.)�#{5!�:v,A�Z(U{���A����Y"�b���H������6�ey���gu(4�⯏b�.Zɀ\�>�	�E�k՘0��!�+�re4�]�q�v�:n��u ��J�  � q0&�ME Zx�gC�/�.�R.ڿum����{H��mߤ��m�X������y^p�|�!���j)}H���� ��>��� MZ9� M������aʒ!jG��-$�ư�gVc_唙���b�تJi���<P���(Vԁl���B"�Q�)���T���u_y�1I���y,U��D"���
C�S�$R������,�d"/�$��Z
�zN5��ү������ض��!H���U�^!���>�WEOèV;� R�ԣ��S��7��@ 9��� ��vI�UK�/��W\��Ti��w��M�7�C}%������ ��ؑK4w�7��k�t,l�jH,���i.ēVhh�����cZCT8�]�G��:���0��`��,
|�9�1h�"Z�s��%�i4�eW~i|ommpfb�h����4�^'{o�C���|�C�MP:3Um*+ 6�� :�M7��LW����L�W��w�,�)#��"A�ڥ�ZXt� 7 �G�guU�mѫ�ه?�1[�jF��l�$�i ��nt(e��o`�D��u���z/m���s��|Pk�P�������y�[!���,�2�Z@�
#raMG�
�v_�-X��c����C�7υuU�3�9������|��J�nƉ3�+�Dر�]N��cieL�4��A����OQ�h���҆+#{�W�7��K���`���'���t@x�*Vg����.��`�U�F��<��^?|	�Ȥ�݃
s���X��3N 4.�10n�R�y��aW�c�>�G)o��*lBԪk��tȭ?��;m�b�U���=�nDw1R�~�%W��3 ���n	��;	�����G)o��ސ���@�bd���<�T�.��-3�EQ��iH���!x���0O��>;�	��4ǭu68���Jo
����x��O�b�ڏ_���aS�M�������}����LRuQ���T�5���=C, V^��56"/ūi�H�������6�B�t[��X��S��`q3��t��j�t��	c�ۼ9Sar�ne�K�n���A�Y��5�ss_%�\�n�x��2Ȏ�eͭ)��Sf���:[����������3��8�����k?�P�˯�>p=�L������=�࣌���% vT=-6Lk�>C�=5b�d�Fݜ�5��B@����{"3�B(<fB@E������"b����T�� �3*CU�� �М�5c�>�IF^���>�D��x�B��j��n1����q�GP�Qt(�qxp�hn���@�$5����#�L-��it)�Ϝ���ycq �U�}�+D��W^p*���$�+�pu�	����iQ�|Up|����=�lE^���',���� M���BXQt������G�)芣*ܷV	� `�<�/;��i0puWT��2Zm�2�𻭿�g��I�x0�MUBAa/��oܡUN�D2�L����Z�tC��v(5H���:֭]MC�M�C��y7�\�]YA�a�Z����P���X�1X+Tc���fR@�t3%�I ��B���E��-&������j1�����WC�!�L���91f�-�5L"��T�ا�Ɠ�9�����7���h�[n/���.�����eI!b���"���'#L9�kCv]���&��)��SZv.Q�U�i���R�Q�J�ѲS՜C"t�6���(Z]{���^}�{u�"oq�UW��z�=�������X�;�\�̢��]L�L��p�7�5b���I�uϢY����.D J�*:L�<���<� =�&�駝jO<��������/,$�)���x�#	��6t&�7}J�
}��R�UJ#���[[@�"Н
{Tg��_ � r�ق'_���{�>��Klp&i)�B^"��f)�a9�|	�ѡ<z�=V�6u�����ˍ���z�����������U���j�9�D���� ��-���Bz6��y�$�6)���9�۝���(��]`�zv�r#l�Y�lg�+I��QY�eG	����<��'�0QJ�%e�����ZI�/^��>����o��u���n�����q�HZ�E,��t�)#���m��_i�,����D}�:�7N��RX/��, m�d�b��s��B[4�E��[�u*��VVFi=�打&8��v�w�.B���ƨ����!Ů-T��zP�1���P��M��C�4 Jj����h�$ePo7�4@g'`�	1�ܼ�3S�''�6ƈJ��*��2z��U?:!�߅�}���]�����	,`�R��SL�Z��g�̪���b����^Y]��ԏ~�6��K��_��=���=9�][m��n|����ݖO�ܓN���y����+D�p��������'����xȦWclg)�	��u���$��ѥ����=�=JA2�Pl���Ú4�g���n�J��K6�n>V&�ΝI��}.?���-�
�c���TU>��w�"���?�!>���>^{Y��z)Z0�#��ٳϰ���Q��1�l[��F "@
��< ����rCQ	˵=y��<����
�e.��d��1��l=-d��T�??xt�7)�-{�2"�d)b*hX�z�6A/^g��Z	�U��'�����v���Tm�G�
d�=N��(�U)��rQ�g�X=$?�끻�s�b�����t��;�Ҁ���[8��6�6;@�TĔi~H&��I��A){I�<�����h>sI_t�}��lo��YT����b;��� �'�O������h�U%��Js��5�����f��5� ����j�)VТ!���L4����R�&e���jA�!@����H�I�B(�-Ze�0%�[��F0�ƈ�O�k�>H�����2�c�`p�������kR#G��c�_����(ƈ�`V�H�/'-��m_)�<|�*j��V�0�1��\�*E	��xJ��F���ngAOٷ�Z:i�0��ca��l�t|�`�����^��)��h��,p��߉-�=��:��P8̠��rp�Ck�R{�V��EQ�W���Su���]SO1���H�6��T��&#�jo�#z�'?�w�"�����p���]Dt?UUq��0u{w!\'-���K�����9�*}���U��qeUx�lY��fΚaˈ~)F؎�X���R�����4��̚�tр�6��DΫ�/���	Xlټ����/8�j}X4��5
��(���@V��d~����颸�_"�=�8ʲ(6C�}SJ-���{0��( p���̌��,���wٔ	'��s�ss]������/�;��G��-{~m�m�9H��̤>g6���Q����ⳮ�:��?��%�s�����w�c+����gL�:һ�6
U�H�������X���R%,�8&�?��!I���z���� q�h;H�'t0���>Q�W<�v��}�����:�����۶�glD�P�tJĪ�����Pd �a��1��ww�J�0�4m��훜9�>c���F��-[vx�w���F�B��i0^j���NP�8:��.� �h�%�
�Q�3�<!p�&�`��!3c~_����b�X�]�8��'I_�6�C��1*�5A�	�Zծ)����,0i�񴔿��V��������X��C�2^Zݬ�
�d���Ob_d� {��=hG�.C#���o�.��n����=�\�R�ജ޵�	���چj�9����/���w��&����J���N�mݽ�EP���AEzw!��(��,;��Y����P�T	��s*�����O�t��ԩ���q���(Xj���8��j�E?�&�0;Ū���~��͊�|樬V�͹v�6��ӟ�,]*����u�C��s�:Ӷ��d�ix�U�N��*�gg:��ʒ����� �ZB6r�6S�����h���ǆ"@#�b��!/�`�H+�ࠟ�8	�sT!��u�oŻ���0�wP�h��u����뻛 �fy@)����l@�z]i_�K�����v"9�9�Ë%��	�'SdE��	曞$0�o�U�՜�_�_�V;Hb�����[����6�xn� �������_-��iV+$���_w��6o���"����^G��x}�V�P�}']K栓l���� 0}u����$�7~�q�0'�FR��� rL�p�+�\��U��1�7
@��?7���tM�X�=�3����Hմ�{Gu��VZ��M1�h�:��u��,�Y9������DF^�����U��;��v7j���+z���IO6�jKqT�}FK�<�Е9 ?^�C��%��z6���H���K/�x�<���>���2FA�[̃%y�L�4�Ml0U��"X0B��_��	��`X�ï� 9�5��r�`�	��Sh��� m�r)�_�j�e:��j��ط�[N"��3"�|�w�7VcQ�v��V!װa��[�;������yy���&�F/-G��~/�rh訨`Os�B�3�����D{cŋv�g�`% ������vKD(mB("�ݚM�E �I�L�d*�T:,�c:'`��g#G���U�1���W�ݼsN�F<��c(�'mY4�/֨�a��L<���؞5���u�]y�$�Ơ��M�ټ�B�K�`��^R~�7^uT{�7�Sոn�~�M �|�/�h[fXB[�Ք�ؔ1�m�M����g~�(�S퍵O���n#h��(ن%Ğ=�lB��,L������h[��X?�p�.�nE#�p_e�������h7~�s0Tk2�� G�v���I�	��xҘ3�j�㛀��$R5-6�׭��	He�dz�E��8q�D������idO7�T������e�,͡Ҕ�F��od����r:j����,,����Gh.����>4<1\�3i������A��դ8(��{��+�k�8�}#���O��e���v՛�I�VJG����2�Ri�O|�V������N��8`<��D0�bm�b��B징����&��C:�f��mT�v��
����ާ5`B��I�h���Э�	~�TE9v�8�la"���8���h��λ�ew�u�0�^
k��[��س�bSÚM
`\�z2r�`��]��JO�t֚��� �����{,z7 ]vT�Ͽ�j[�����G헿���x~����] ߰�O�i��������b�`��	 ��  #A����sn2V��̨Ӱ<G�,5tw����$p4���iv�+RsM{WL��F�J��1������ZAm�r�T�M�i>v������P�'+S�+��
Z-�������T����s=���ԥS�0�pT@������@OLY*1r�2����8@̷��{V �S�L����4���(���f������a�ٟ��kp�'h��������D�V%�v�F��u��D�Y���Aؑ�-�(�j8�toq:a��!h$yd^ �	"0�4�xO�����Q;�
�����Q[X-J�Ħ�J%\:�{sU���I!b���i��D�6z�D��Z�@��Uڢ��0N��T�Z���#�$�eRx��H��DԮ�{���JZ�B��4QI{L��B��J1�]^��L��/1��׮[g��~:�{�xsS�����9$�:M6����������z�b!=�o4lIY�>C���v@����ٹ4Dg9�Z�����`�]z�%�6�^C���-ˎ�d����r�O�o�0���\��J9]K��tPۢK.�#U�`�x��c�I� �"�G��*���6D����#Lhi���n&u:�ؘN�ױz8��Gz��^��~1�H;��^n�N��;���/�BX>�&�=�|i�-�@uz��!c��sfS�"m^HQC�œ
��n4&�w�@����93k��e|���^��C����Ϛe�h�Q�@^.��]ѩ��OZ����18e!3���ؠ��ȫ[� YhGbd�BP��-�D�X� ���v��m���.U�Z뗿�Ӿw�g��}&��JvnwO6�!9��A���)�2�]�a���wh�"f6 �H�`)�,!�P���KI��b�4O�	.��,��{ֽ'h��#+́Ғ���8d
���{{O9����M@ ,(B��ZsW����������O}�_A�\���B���r�G�&������~�����.�n����t��<�l��ΠH~�ۨ�x�����0ѝ|%ag� ʇ���p��܏�7i�. l&�?���"Vu��l��5HC������������]�U#��a}��KvxQV�݊r���}�ӎC�\�����m�dƖ���J��G>iw=|�=���#4�'��,,����?���6|���Z*�?z�Y6g�p\��m���;4ݒ�,.i���^~%�8f�)�:�RH~��9q�C2.�+%
[I۫���D}�-a8�	
\��kN(YP���'��`̷7��1�w� '$�	 MhO���cb�=3��J!�u� C�sT�C�������a}�>@�>�����<:�
���q0�k! &+$�퍿�Ԥ�m��n�{v���㼎�ٵ��=�����I�\8n���T7�t��g�y����VMP/��q:c*.�q-�*�-zzc0����p��ݟ{��}�]��n�|I�~��fd��?y ur觼 �M�������S\/�Q���P�����\	5Q� �����0��`S@��T����%��b�6R}�YD�O��|�:��"�$���R��UJ�&s;6eI�s�N�H���6T��S.����Ls�zL��������4�s�d7H�	<(�����k���)*TE�40>� `%}!��F�2�Ԛ"�jEa���i�=g�l ���Px��{�48�L�'�qFm�ꑩ����͘�nߵA��7x�ޚ���b|	�����U�,S�뮿��Ǟ~�ILp���Qm���0jEl�AKwi�J��w�*2.|��m���wg	��ڢ���tz��&��B���G-YJ+թTo=���m�۹u�]{�en2X����3`7c�7��'�Y�����І��w|k���̤��^�yy6�4�äj;K��m��`cF��K�'^�S�2 �޿�N��e>������р����_lW^�A��=�Z=��O�9�:bmG�N��[?��}蓷R�>�~�G�;8�+jM�RAp3���f[Q��k��_c�cH�K��3����#<�q��T�vيE�X#�ԭ�~�~�S~�����o|ߖ/~���b��>���Ǝ]�%#�t�dx���U��jV5�W�c>�P)���jv��C�K�8Ӧ���%>� )E.��Ov�u)���
2���Ŋi�>�_���;}h<�=�c� p�0ڬ�kQx�
�s�u������I��� L�G5�Ƅ6���(���ٍ��c��]����ӷ��=��+v�WېQ�����o0�T
.Z��}��g�	N`A�8��Я�A>^�)�A ����&���i���޸TTzƂ (�Y��4�cAg \��bUm��ҋ5`ɢ�� ��j�!EY��3}~n�#�B�qTJ��Q��s�˺�d�}��� ˖��,��Ϋ��V�i����yk��3�����dD����sM�Х��G�$L�ǟ�A����Ā�+�^U�k�P!�'�ܵ���Ar��}\��Rݺ���;�+��)���9PRzE��#�髤��f]�������&��s���`���'������p��  ~�k������p�p���@���'O6N�}�\���?1r����M{8?s�	8ט�J�� υ�I�4�}�e*���8�	ƫJ+,�0���C�Н��`á�K��~��s��Bw������R������i�T�CҔfut������~��a���h�캵�.O�yY<���>�uw%�u�[҆Ly�h�8��eKl��.���w����i����VZ��Z�0i@FJY%��n��1>��mi0Z�mE�5R��3�6d��jP�2�r�΂ɒ��M� @���bWW+a@Ǻ��OK���.�#:�%:�e�����ie��kc#�����'Պ�+\�3O�!��$��e�����R�gC���`Ϧ/�<�T�)�{1|b�9�((d�w
t
+�ц����J����!m�#��믣��~-$�}�2����ܳG�.*��̙���-u�b����JI	Θ5�ݳ�+(�x!�b�����/0afՕ��}4��bE��KՙM��g �����83]d��9�A�m۵�2�u�$v��J#�#��M���a�����fgM�MkV�?�о��O٨)'ZÞ��ɸ��K~�>�6��}�	)�ܑ�X�K6[ن�x7��I�G�x���o���d��*�X�p&�,�iAB������M6��h�<�{m��
�1�LiGZ���B�D.V�ڿt��M�>��[i���w�۟�n����j[�/�v�6��EO=>��>SA$��uuP�xL#� c]f�նh��1��FZ�#��r`&1���k/��"�����ռ�c�ˏ����μN�2�(�I&�����`���A�<����2ν�6�PPx�<������ig/p����z�`V�h�`��`�?z�-��\i�ؗ��ז��z��l\�_��i$~KMX����b��7Ё����|�u�pZQa\��IDk����i|eP>�E�$��^l"I����U ���n����E�XU�N˱-��xBMF0������-u�t���z�*�׍팊�iHH�PHϘl�#�ׅf�s��_ak��~()϶���,B{�=���{),Ht��9��"֝4֒Y��D5h.���i���)���6t��h�;��;	��vJ][�t,�i��0��'�u�0@��F�$0$+A�pP�� ��u��"�]�}
 L�W���*�X�r��:$���'�* >"�W�>����׋��d�d�!i����~-H�If�@�����P�R!
� �HeL�k�n.��1lt�wh�y��Y��?)��Y&����=���1��"�޴xA��3�b�ݖ�04�{8	�⭥U�)�3gp��фO|����=�N81|����{g�PG4�}�@�!��0�
љ:�@�!-Ot����jSU�V")�6��}�x��ѿP�՘Q�-_��>r�,[�O��ldc�ڷ>%=c����l'%�L�X����]��.�l�]Db�l�td��D���P��]3S�'K��q���B����Q�tvAv
J�*��މ�&�ג� J<�Q��\߷�70[�0lny�#����|āي+g��Nډ�h6�d������z(B��2���
��; ���㘱a�������i&�Ν{�$Gx����Un��k��D�ͱ�n��hA�(�u�3��IUЩ��0KJ�i�"L�MRf9\�2\�����;O�\���G�<�䁦����Փ�7DLK7�{ ���ʞ�7�Rx~��_�hRml���KOĊ�����ؾ��ULňB�1�ǳ����V8]��X{�����/�j��Ke!l�B�2��iԾ}�˶s�K6������)̥�Q��_���PҞ�m;���k.�	�����G��Խ�a�-�|�K/>���#T|�a�9������)m��6R�8K�ϵH�F �~ɾ*ڛ�۠��#����Y�x��)�w)��Ij����;�;�m?Պ���]��o\k�|�c��?�T�f�e�S��B�UE��[��pjD�Q�Z�<R�̟��ܿ��]�#հ��@�ޕ�L�+�P�oY�(U#[��T�NF�q��}�0=z��a�4"� ��N�. ���}FL�$��G�M(��&,|�u�mXl���ԋE}u�)h&P�����5�G�x�ָ��Н`�c\Z4�6�u��'���%5� (��GN�����o�e���WU�7�tc��"��|�gpt���n�L�� �B�԰R��akI;����"�Ua��k�9���?\�H�Scl����ȃ����ˬr_��,jJ1--�,�W�6�����V�[Su�uХ!�i�Z�j�Z��ጳ���\'�i4l���z���F�R4@ʴ�4l3�
Ձ��d:h��F�\g9�&��DP����19**S��90�x]�&�]�>Ȗh��uj飿i$�-��A}���V-j�h3����SoP�0�g�+#l�j�1�7�>ܝE��`(�<ը7*x ��:d?���k]v�'m���dzŖ��I��Ԯ��4�h,C�Q�n��-�6f�pZ'd�������ٯ^LS쑖1�cE��?�����}�2�D��e�]{`;�)ʾ�L*UG#�8���y�b����&�dtO2��\�E1H��ށ0ZAC��/������a��k�F�A��p������=�=��VEQ�*[p6O�e��9�톋O�m�س���������z;뚋����΅ˡ�q�U�R�y��9��O�Ŧ� �)QD�M:�$���7'�j�|�YFQ���T���P{ X�I"Ww�EpjQ4Ax�k����g��;��L2:h1G���o}C��E�tM���?p,f�ȹG��p����~}~#���-��.��.8�roU�~�6��`�$�Fi�gͮ�4�eȟl�J&Q�0�H�Fg���6c�����~w�G�2���nߺ���ͣ�4p	ѧ҄Dt2s��ٳG�!��HOnļt�y�{������,�k$���Itt��"�,����>ѶWu�FK�,�΁��,��0UQ,�9��I���hw�`�U�5aT���n*Yl��z��8�O��+W��{a�����;u�۲v%�d�(m?��?���7���=���'lΙ���sg��/o��k�������g�������`����s4�vҦ+����wI�3j$]h�[Y�h�͓*�z��v�À�����/�]��e&�������G�2�Ԗ)1 졓�m͖U����}�[7�'?�y����g���j�����b�dlL �TJ\������B���(�I�Ja'�W� �� E���l��t�Iΐ,X�,��`A�ݾ$���ݝ�5�CN��~.((t�X�[�)�)��H l^�@-��GN�0�r �����&�:�o�A�� ��� ��(��S�o70��:�X��Xjº�>и�u�o��&㩊|�����ʾ��?�¥k,}�$���Qc�f�Bg����� HS+Y��y�u��m�ފ,Ė�(9T��F��S�6Ɣzs�2�:��v3�}>��5�R�F#�~ Yk�`��l��	�$��g���yН�6��o+�o��O6v���a:��!
��4˄:{X�=�p�=���^��W��k�� �XgQ��v�Y�H��%Tcο�{��g��k�@�_��.֠M|�lW�hh����.��V��q���U�O@#�n#��@FC�{�����] �B�1�O^�' �*�Һ/�z���w1L��j4Gd�-�:�������}��9��ᴡ��̣�-� a
#��M�"��<	
��I�3z���!=�W���u�{wJ���;.V�N(���=�
�
3n��9�Ď{ڕ������p��"d���Q@k�WRUS���~�cS����Lh9|8�R��aY����tqc	=��1�i1��ѽͩm\͔����L��=�NH�(�buݬ>*e��S`��)�h������1���|�%r�[�)K��y�.36!!�k#��#>��	S��U� ,��!2E�A�T�� ���D�l�*uE���JE怙l>혪^{�L�������L������\����{�����#S���?r���J�"�vZ�@{`g����Ȝ���u��B�s<]�ͪm����u,�f9gQA���e�7�C�6�ROF�� nҍE�Q**�C���$�P�$�}Yi�7����z5*�	#Ą���"-�*H(�'� U�q G�:nP�Y�,f��H���_po1Us�A��c���+o��Q4���e,0�b�|�:g�Z��1b\逫U�ϼ��[E{&Ķ�֛��=�g�{�9?�L�L- ��j#��v��c?��7�.E+�-N�-�0�-��&�U0i���#��Eg��;��l*����>7A���w�6���0	�jݳ~�詤l��e��Ԍ�-�|3��>��r�0��km>~]�F�����_E�ٙ�����V.yզ�r����/کT��}/�G��'���Mv�eg۠�����_�'xv��+T�]y����ϲ�;��g�sˎ�h��q�IO�L,1r���V�v]�l4�Y�E����T�]҉���K�p�o���50Y#�bƏz��������<�,�y�������+��~��_�*�d�䏄îEѬ��\o�:&05�u�
P�6�`?��L������ (�K��j|��J	t���k���b���S�|��S��uBF�JK��Ġ����0H
ر�#`
fӐ�m�ka��I���td���md��Ĩ0�{)�HvD*�aD��m ���m����_i������E����
3�B��&R�,SV)��F���t)H`]R��c����VY��	�����4�Ux������C�1�Q�KF�E6O�ϼ'�,b��I��Q)���p��uv�g[&�z��5��NE"sL�ͧ�}�%`ƪ�\@�l���9 �.��jœ��k�����Z���w��}�^/����돊O�����w�T�۶c�~[��*@�nK�=Z�Z�2,?�>q�u�U��*��=	��d�DK+Z�i9�`݅�p "�E�((�rCW�3�Yc�&�!�a1J�ᔞ�������u��K��B��u����i(�G�+�4�[?(=�|�Fs+]eP&6�9��NK�:�_K�H��F� �~�ν�g���'����(y��Q�^��T����*��j*<���8g�6HFӄ��^�R����Ixx�ӵe�H82Z����K�XK]XFܝ@�Qd�|�Ė鼻jK�(%>n�̾�ڹ�Uѵ��um��ٺa�A��J��&�^��v��q['3=L28	�O��~A9)��WH�[}�1s0���*��&��x�Rywpr��[.�������G6ϡ�Vb���uMHC�ysm�f$�RY'�΅�S�0��aG����� M�m�ZD)(]�1�z;��Φ9k��N:�Ν7�vl�hŴ����>�^D����9�<Xj��c�N?�N�<�#�-�K}71!Ye��ў69Z�si�����Hl3@�j�������^ j���x�pQI���1V~Jv	��a$��p�� S Rtv2>;)Jt��~@Wԭn�&S0�@�N�Ȅ����=`�"S<��+��)���Qg��}}��x�0�1�}_j�z�i�+9��H��L|�q������Ƥ�M>u�U�Ri�Q��ǬU9tk���*�F�+"|MpOO����1Tk$�>0�5��%������
��K�o>;��P�i���x֍��Z��w�b=������t<��XQY���i��
ҫ�|�m�)���0Բ@N<��2gv�����-����T��:I�<������Z��mv��0�������9�rS�m�9����V؟�|��+�l� ��+�暣��OI�ՄL����5��v�� �1��* S�	� ��Ed�:V�J6�=��$��5�(7���$��*��o<c��ϟ����b�a���߰�XDɸ4��EU,�[mNZP�~�h9����PP�j&m�4G�L�s6l�� K�)e�h����l6,��.mZ�f)y��3<�����`� �i�� F�s0G� ���8�%������]�������
ˌ������1B;�ھ�j����f�=�T����Xְ�T��F�w:e.��@�5GVEr~\bz�>���+��@�K� Y?�����Ŋ+��|$fEVY���6��F�V�(ާ���ϦUQ2�g
�so��R�|k��_q"J8�&|�:���Am�6va�!�>�'��p�G�,Տ�tƚ��L��n�ܞX��vU�9-ʵf������M�0������-�|o��a��a6��eAH�%����8;������]��@ ww���^�bEZ�EZZJq�C�@HB���$w��]�9'	�@ߖ������Ng2s䑟����kgD�X\�O8zo�4�?���0a���֝7�V ,� P� P���@�4O�P�@X������߾�v �����*�K)9�kM���]�#���������v;k1�P�vz1V����Đ	����Θ�ң�Y^���X���!h&�L�9j^�(`��,���F-��B��Yb��i�����-b�B�_� �V�cv](��wv��@��u\�����+��d���4*�X�R�gCi�і�k(鈤ODC������#:G�P|SGTT-�1����_{�����s;���jh�%���@��jE��M~�}����}����X�#-�#���q�D�tL���it�h�}=<�44l�@�@L���2�L��"��1d�N������u�RF!_{40�������m��>��uO8`���״�[��4��՚%+�H��&e`;�?i����K��:�6����uZɺ��
9VN��Xk+�b�t6^��Cn�L^�>�]�Z��|���v�h*�a0D��"NO�Q,\i�NؕT&r�^H�j��"�6��T	��6��]}�J��4�@.�;E���bg�s��A��$	��)�*H�FU1�I~��g�1�ϵ@���\����Id�nL`S��U#z^�
����&.�EEN���`ZMi�nb�+ҿ�7iE�C�o�4Aj)`u��Ф�V�Y�	B�X-��:=� q��u;)0h��1KK����#b+��P!�ۉ@�2� +�ռ�4F���Y�<<¾XZg���������E&H��R���[���lB�9��.Z�f�'��g�T�&�y��ڣ��{>�l`E��zP$P V�G,U�R�46Od�W��F�Б�F#��wi��d)0|l�Z�XR��c�)	��d9��ο�yr�u��'�Ϯ��R���q�+�K#­u7���4�R	;�ك�ƜW�o'ca�r�����ji����"���M7�o	�����iӰn��L�7�G׉�l0�~$�s�r�4�����;���?C�sjg��M1X�i�}c@�B��
�_�g{��]r�]���s,�` ���z��֛����ߺ���)�����1;yyA7�֯R
XI'*��P�FJ�C���դ����N%�Hfٛ�eD�3��ݤ�����XG�p�u|o�a*�n������[X����V�_�I�Y\�?Ĩ3�� |��g,���6��VUy��Ta򁄒MGw���H�8x`�Zco~��f/�d�ѬN5���sw�[�\
l��k-ˍx��9g�b����l�.eKD�Q��6*ɬ�ѬZ�[�/�ZJ��vP��IV�ρ9vr�v�pJp�Q�
o�����5r_��� L��*)C�'��s���b ��q�~��(=f8�N�k1����%Dyj��l&���ثD-v��}�S���X{�H�8mH��ĆKFb�£[G�sV'ou�U��Ҕb���r������"��P!��]� �NWڎ���I�0k�&�����m��q������
:;#�t�$Bf% �UN-h���
*�lh�W��C�w�x�:�Ck��BI�9&�&M>��:?�N��������]���z%�C$ ���%��H~��/45���_a���t��J����Qh��X�*�SN<�N?r*ɘ���� aET�ea=A٘�]��63I���Cw�k=���i#��ksV�{�Ť�z�N�MQ���cCK����X5��
ʫU�B���E#g�����  ������١��S��(�*w�����rJk�vI���Be�a�Y���{�SѰ���>9��?t��,ŤhRY5g�b��t���0�/�A����)hjF�R�.J�p�8�g�QD�.�zI��g��Q�W=��Z�$C�[�pAĊi��SFY.f�F3A�p��Rq%&��fN�O�*:��E����4���)���'��=�ͧ�*֯�O�t�A�K7tN�8AfO�:)^,â5O�i������B+��K����m0`��T��2�����fݑ��L؜bl+rٸ:aZX����W6+v7�	,Y$Սm����Pk"�M����&��zUR�%r��b��7�уɕ;��S�7Ix�����Љe �-���U3V �)��X��k�����`?q�]s����G��3���|p/�Z)����w��j x��t0�hx%:����#��vU��5:O-�x?U����0�U%dYY5f�����|���� m��y�9�3 �����,���p*����q��X: �&�|��j헿���}�1v�ŷٴߐ�Hj�H�SG�z�[�X�dH��%�����Ӑ �:��-�+�pĒ.��K�2U?�X���5R

[X�ܘwӺ�T$�1.1�$`q��f�#YK�?���Fa�:|��/�	'�Ϳ�����Ux����ov/��H�h2~�:�{-]&�;�m�鄢����:�V�F`��ϳU��}���֭����`��z�� �N:� [	��R��k���b���~�Oe4"~���k��#��$1A�1o_�����D��>ʅ�\C�cQ��� ��)�e_�*K��P5d��
�K`�!�o����ri��Ӵ�{�s軣��5l�� �@���O� #���d����}&Uo�V�1:H��l^��� ����"*
;��z.�)TVZU뀧a�tI�/}X����O	��~�\3'������Wn����	�狍S�&�o���JU��)/����z�lEt�3�Sxm ?��J���څdSa����v�����u���B�8T�f}m�o�ި��{;M�)���}'�ϙ|����e���`�l]m��#���f�p�IGٹ'�cM�[ S��O�+Y���Z���eP~�ˊ쳕k�����O��=3������M9� �����t48����21���F����86�4��q*��Hۋ$6�V6�6�L �L���d�?����4+���ޭt��k�&L�L�
 |���l�������P3��ߧ������Y'��m�>��1�tY�P�ȁ`��(�dahQ�O��JC�l9݃ؾV�ki�X�"4I�����]C���5��;��*�����bI^��0TR��B�@ڜ; ��\cM@E�2�	\������D�)�U�n����7p��X�S\��D̸���uY�ύ ��b�^SB�#]����]/��4.i�V��.�a2\G|�-��}g�R[\��z�i���Zac�M�<�2:�K+1��}���Q�0�YV��VXa��0)m,'��i=��Fz�@NH��R#�^{��ߩ�УZ��Ѭy���6p@?+�'f�k�Q�RL-x ��I6|�����d�1i���G&۴���g%Xj�`[�n��x�#���.�K�:Ϟh��-��Q��
<Ԅ;.��Af8PP��H9y=��Y;��SJ["|��q�@�6t��, H�
��_��A��?�c~��<?|��8�����H�0�?k��//�:O1��]\-;る��hL}�������{���f�I�d���T�1�d�Ц����P��q�ϧ�(�S�AP���%���o|�>AkW���6��5D'�r=F��V��֊��̍-������S���:{�B�v!��#X��x��0��m׉(�a���v6S�V7	�H��?�X�͛�+k���DH�&����s
Ao/�m��[փ�_��b�=��_l��6�o��u�Y �&��Uv�A#�_h���U�]K��:.�U]R/�7=MM�a�dE�����*�@
V,���xWI�������^�a�7eB�r�4_8�="�8���˒29��Z+�'�^<8h��QE���~`.�WO�ewY'�j����������\`\ ���0�Щ8�LΎ����U��6-��+���Z�-mq:j��xR��LC�:7�o���N�@EQ��~�d\/�]�(��X�5�uK�	]�nTm�9
����:�Q�}��h� S�A{�<�"�:�'���پg;\	��!0��9�wK���%A)k���1��i�S|և=��?SI�����|�t��q��	&/V{�>�N>t��k,�`�q��	�'i��T�!�}c��Hک��K�=�փ�e�ͤ��[/���UiG\p=���|�F7�����j��d���"���twl X��p{f��] ��hET��t "�i��@�[E�J�t�P<�_�vj���y�Ǹ@��� Q�)�C*����DQ�v��N�=CʱYO�V���Sh��IƦ(���B0T.�Ya��"���Px�#8��wRq{��G���T1#�����^�n�	���q�Lפ��К��\l�n�G��.���ĥr�W�;���Dt\�DT�-lRM�S�{ �9�G����7�e���A�د��;���H��1-f�A��S��o�������XB����,��Nꨲ��{��[�v
q���bǟ��=��{�����.�!�iVA�0f�P_�N�o���Ы6wC%��:���nE���X�ħ��Z��I����Ԏ�d&����۪Ѧ��l�I�H,�1ֻ���C��9�`]Yh)*ɒ�j_�&
Q��F@�m+�h�D��n%�6�������Mh�ncü�s��;n�_�{�7MW�ni�Ra�t�e��a=��*E�	�$�^O7�>}� ��y�.��)�(p�1&0VCjL)1Y]ӺI@L�R�����Më�t�C�OA��ݡ�~���l�˩����}?���J1Ջ�`>q�v�	Ga1�-X��R�4%�U�
�T��ت�S����mv7� �V]S,�˷:[
��1�}�.�l��x��qj]�EqQ��w 1��-h�C���V��VZ��0��gb,��U�ZM��El����uߘ��/��T��B��>���o�O�}��J�q�뒩X�����YI4ߛ�����uQ!�qT�4ec^�v����-75[&�L�-l�|�4�=s��\�VE�����5��ӇF����Q�ǆ��ޚ��Z����s �<9.	��%��I;����� ��Q�l��?v�@c�&���s
@��A5��Ȝrp#�^ L�$��5���ٟHw���\�D�����v��Y��*:���%?8�BzJn�9�5�9��RW@@��'��m�B�q�|�C���C�0j�)0ӹ�zX�T��%�G��E������=�����U��%��Qu�w���T���C�j]}g�|�r�%��5��iE��f�G<�{۰S2*�C�����T�+�n��)T���ZZВ��O�ܝc_͵l�ߩ��O��.���	�P�5t5����G��$��OeG� �0�4�,ȳ3��h�̲s����
�Q���ʲ�Z���7KW�?����T;���lR!�|P�Y�}�1{��w�ŧ��o��nGwsߓ�R9��E �ˋ��ͬ��.0�HT��G�K!��L�.	�)9�̩*��شm4,Qb���y�HJ�J�C�������\�뀆�4������R����u�ݩة=|Uv�#4��" ������h��hP��1Wڔ��n�����&Ri>~���7�(Q)"w�\OI�8BE��b�@���_�͒Xu�-4Ү��n*Q�*�B%T#����X)8Q��ʣs�e�	T����#a>O���U�$ F����
�����(����	N��A��K#����٥g�aW�w"7���o����M��j9=S�����>��#��¬���M�mI�mX�ۍ�V��ݞ}�>"�,����v)=셗��Ȧ�L�6�?r ښ6��3�=�Ə�Ŗo|��U������E�`CF�������5X~f��<'3�ƌ쇧R����t�L��R�Ÿj����TM��z:����}��	�)��6)bz�?& h{�]ۊ#��?�6K�eV `D�	�� �l[�~�=�����+~a^u��w���z�J��1�TabK�h$�cd���8X5&�+VjhIR����W���Т ��_��V]���+Ŷm4'�A�\�Zг(Jغe̚l*䁨���/A	h��g5b�楍F-w<M�e��_1�i�x���0�}��	��V��?�}���?/������/�������N���`Pl~]虚�[(:��s��#���n|���-�{R�YX�`8�N������
���jS&�k����UmT2�q��y3U���T�2f�E�m��+
 <)�I����a�Q��N�zz�¬��a}��7l3U���`+��U*l��{ڕW^j9U��;i�ݓvoi }������b+����{w�>���Iz�%������Aͱ}��:(��d�}��C�%�uA�����R��l�uv�mw�	'�k7�~����hz�R��2��T"
���=z��%��4�5UDv��K
�cl
Z79���!��k 6]�V!YS0�D��	@����b3�.�y�J[\�I6J�v?����n ����t�Vj���1c�	9흀�����Stf��>����}�Rڭ��)VUBB��Ơ@&4a�y%X���i  �.@�&�;\J�qQ�_<�+@V��/sX{B��o+����n��=���c`}��6Ry:��"�ֻ����MI$��y7M̺n��	��- �b�� �i>�+ÏJA&PCO�y�g�K���*�}����C����Ue�2u��8dx��D��g�i5����?~6s<%���#��@;ڴ����e`('�M��,��*6��,L@�̯8i���{�E�^z�	h�����Ϩ)���i�}`El<]0/�}��؏��m���6��k�pLYE�q�~��'��[�ko��n9y�=��O�|� =�geDS�臔�i�t��`j��I'#UB�W-�;�� T�ٽ2��wJ7����Lg2���^��-<rܧl�����$ų��KV
ҔI(��!��7�&���!͘��5p#H�Jd�({hs�m�ƋQ�Az-�W����N�F$ύ$�i�vA^(٣3u�gC�.�h:R����y���h��҄�r��5��Ԡ��T�Z�h�������٢~j�V���$~��f��.��7�����Ge���0cdFO��6�z�7�w��~YHt�H׹����+ke$J�	�j(���f��g% �D�C>�h9�s>�k��|���N�/��ڪ��!j�1��HJ Q��-������U6�hŅ^��&�[˫�o�K��نb4���˺d>~)�'U���[����;v�O�$�9ز
�یś��s,?��n���X%���:M�R�Xm�3q������Q&p�� ��?ۖRaٙf_�a3N��z	�ȅM��X�w�]po��}�-|��o�-L�#D}Qk[jDh�r�{̳O,����H��3�G�;o����̆"���L)�VRH�p(�S���$�쵰��^P+��
�����S��ν��i�l@��P��Z��UI���7a�"�s<z@�����C}�3��ԽZO�դ��d��-��Q�2D��1']�o �s�Fr��Hx���^#�]���耂�I�Qz�F�ͱj,v�t��*U��h��=�l;�C��_>�ϻ�c��V���sKs���j-�Z�B��w�Ͷ��XXl�k�QvE'z���#���O��~�����瞷���w�I�a�P�<�'���=b�oLl�o}�A����<+�Jg6�3/:���x��[i# ��LK�I�}�p��J� ���=�����xԚj�-;-�z����c���Z��]l�J$%��(�ZH�� "��H*�������s�=��l����v��O��W$����v+�[z�$���&���t��V�\�
t�=RX;X#$ya�P�>Y�� �9s@Ę�w�k�8��@����J�l*�?x��܎�"�)�/~-�T�gw�t��ەFێwS�hP�53$�
��N�T��G�!��Fė�+�Y��l��"�OPH)D��^��1�n��;'�z��'���2���,<WD6�rU�ꝶW��a";D@4�a��u��&��6\�)������gw�W�<���X�BDF��:/�]�8W1x~G�lԎ�^��;���w�1/A�w�5@@:��rU1���.�6�D�.�� VH��[���R�\��bG&n{���a��q��'�cqz,����\&�Oф�`�֤ #f�PƛЦ��:��o�32s��W�jܿ5Pn��F���,"������@��5�^� ��\g{�6ɞ�y����ʊJ�Ѡy��!�n�hк\@�^6;$��z���q+BudQ�M5���66��hϲ��=o����Q;±n���Ȉ���{�S�CFN�^X�� e�^���.\V�J6Rwh`� �S+ ��s{p7o������%$�ӧ�Y����*�hS�Ȩ�[�=	0qj�T�b�'�;Q�m�!��C���!�N��y�D���b ��&: ��HJ����,��-����T8p,&��J��n�
�!K������ϔEI�S��y4�;�&CZ.�Dͪ���m�x��A�x�E\�D����$��ՕXh RS`M��J}��X�bJe��N�1v���ں5��7��&�2�
����(ʧ�@0k`Z��; �6@���p�j�l!�W#��(�3
f/���eU��%`ּ�v�C��&��>y���s}����i���`��U�[d{����Խ���Ooْ�E6u�a���9r�)�%��ll�Dʺ�>xi���x,m)�De2w�YI��"���zwX���r�C�}5s�-]Uh)�0� �55 �.˧	��k�!���'������T������זK�*	�WQY�w�H�(�5ۊ힇�j�^q)�[���lmW�����AwN������=R�U)��5��� �T� ��J�f͠L�F*���l�r��J�V��B E�A�Ƥ�l_|#b�×ȸ8x���JL�e��@ʬV&��Y��Z��c`������:�!=�{�}�i�	����~�?p�&��
 �%	��2H�M�21��B纥�.��<�<����.�㓯Z�!�X+�5��k���'�ҖoW3k��	#l���b������o� ��;ؾ~�c[4�m�d���GL�5��Z�b��z��  i���m��>v����g�gS�a�=�+G�xɕ�Q��ˎ<���H���Dy��Gc�½����{�'M	kM�3o�7��_��%L�o��矵�����s��/;��4,#Ff��y��oK�5[a9~[���G���'OG��	�n�M_��o9�,�F�n���!�zЁvH���v�2����ڱ�b��1�O�Ъ�iA��V��2B��Jk&0&ZXs%��{E���kG�&��� _���mءs���GD�������?��`(�v��XBi�;��=��HX4���4�m�_<�������@'h��!�&�ymE��	੻���,x�zp�=#/J9(8����'�e.���4*Nr�c�NB�S(蒆O)__I���AC� ��� u��PE��R��3R��l���"�K煏[��gh��S�t�V�eKNYT����bl;*%� ,��v���/��pT�6G#ѻ��9�F�L���%J�~����F��M��<[�t�l���~T^,��9s��SO=e�׿��?<%|��C��cH�$���A��v侣����M��
RNx0%��� �����K՚c�0P�0?1l��l�e�$֐�j#��=?F����#H��Y}�^#n�,��͸SY��e�1h͈:�^�q?�7`R��.FV
�l0-,B\IIy�`u^O?>�bZ����S���o>���,�
 VRyCZ5	�Ң�E�(�.������A��R[���	��:�J��Yta3���ꉠ��k L)L` @�|B�W4���k�y����{���w��aWN�[���NV�WZ)�3E�	�����Q#��ᖌ�֍T�Df�:U[��X/N�e'Z���
�x�eÎl^��JL����U4�������"l>vq4x��5����}��ߎ9�x{w�[��Ԓ���y�i�K�1�2m�� }D�lu��Ӹ&���g�q�'�|(����S��uʵ���>�%�5;~"�Z[���'z�؜��e�m���f���_|�ڞ}�}[����'��@�ZB$ނ���)��4X��[`{�s��'�m�ﻏ͙=߾�j>$T:�P��O+�-0���o�z]��K�q��A ��)�\QMJ������*�eP�'U�<,6�1��|�F����a0n�ko����e#=>�Y>�±���L�9r:���c䍣%I��י�P�)0O+q��e���%�"d�]�l�=V���Q�q�s�&IL���ʫh��J�N��\�my��3�g�VR\�d~:ө���*�ՏN��N7��ѥ�?�OMyU\P|���cҦ����L�F-V$%�u9v޹���b_u�����GZz���f+�?�W���J�^e6�o��C�?��������/��C I��-8�0}���;�_�kq�ͥ�Q$:�֙t����]F�Gu� ���lݦ�n��K�������l��іK���S'��o��m�[���&�6�a�f�c�l��������/b���1�l-n�)l'�z���Q�����(�i�˰o��M��A��D���=X�L&H�#�}��׬{��٪�h5ڲ�=Ȯ��:R�(����f|)ʀ�.�6JC�:ӈ�tl/�W�Bx!��F�"��O,[X��C! ��?�B�/m�y6P��kŬ	�8'b�Bp��M{�|�<��S���ڠu?�`ݝ	���?O��3��3W�(s�$�^)Y�(t(Boa;��{�#�б�*w�_���C���
KQ����D�����d��S� �<!�w��p��ٰ��_�k�FJ�)M	���z��_�����K��Svg�<���v��=�`����l��N>�1�V(�8�% PZ}M����Z��=�(�}��t\����=0a�~5S�!v��G��^�n�I[����S�.��
rs)��� �F���N��(�t�$�-�)�Mk�x�^y����c���.�穢��v]�}x5u"�i�:�K��g���Y0 �8r��h���id�*��5T�ы�m4�Q%��eH�*(#ʛHҝ	��F�%Pͤ�	݃HD��w��H縻��J`)d�71yw�_~�%@b�{��b(����V�5J1�t�E�SnI/����
��� e�5����,&�ӧ\�x��y=���t
�L>Vh���TmY�/D*x�gs��V�1ٰ�U�M�#�"�{��E�$I�B�W	0,ڂw��m�\�gͱ}=Ү��f�������f��*�o��O9��n�����%u�oF��Yw��s��t��/i�:tZ,����w_g0�,�CG�wǽ��eX<o�I�߇P����MWr=�a�o����VU�ۻ"�� �LJ��%�hC��@�Zm1)^LR�"�QJ�Q�����iν?%�i�zؒOf�.�\�7�ã��T-����j_�t��k�G!�pW{�&��Wu�6y9�H�D�<GJm���èД�e.��נ�~�bR��3 ������~[2�k�e��+�9���t.qʨ����"��h��5����n�ʸS�d<����\��R�\����M���A����F�J�Q8S�=�~��9���Sr����k/
wV�Vk$/6J����l��������_~"(�S�l��(�w��׻H��: ������?��;�{��WlѼe6z�d�Z�j����4��i�A���}�)��n�ﻻEp>x�u�m��6y�ݐLa�Cbm�:��%߮�e�|M�r?�Q�غ-5��*�J�XnJ>��H���H<��@*{K�S�m��=�ۛ�a��EVV^�}8�a���w<����%]��_�nLm�$�Od�8x(��R�Z��`�ij?�"R�l6�T5�1�9y�M�}"��RU$#0鎍Hw�_�����|�����O�{�y�o�M�<��,'� �d���V��`�Mܯ3fdXlD h��H����18u���f�/��������
g����?:�0a�����́�+ނ�P�,�ҿ��g��|y�P:,��{�| �K����X_H��g(+$7~緂���   IDATX�²5�z���K:j���h�\��,��T���B�c�A�B���k!_Z� �Q��i�8�u��
=�� ,@�)@]��C��Ib�����r�}2��F�/����~�����>� �������W=�lX�.���v�J��}�x������{9�<����#�! �e�^u��w�~��wg�jʕ㉚���qIa�ZA���2{����ыRv����d 0�uK���L\EERJ
Bph���$w��䚍���F��I�&��hl���8Vw��]�Qa�f��$]U��c�����:T*��7wr|
� �v��$-葄�Xlp�|~�l%Hou4�<,�"<]2_~���!�Gz�	 ���U�c�i�V�vo�$�+ؘ�Yh�P�WCc�j�
�sʧ�@BJ�U�&QI�Zς��쇘�zA���w��$Ѿ �[[7R5G���xRC�ҧ�cJ��v��Bo�!��*���}m���s�ҕTGF��j��X%z�N�,@rB,����l���������>oI���]�	��>�����_��Х�xUR��T��~mO����fTЂ��J��dD��7-�{��Lڦg��P�f3�o��^z�I�'�Ͽ�E���s�����ʵz��l���6(�9iAT}�.��?��A7���F��L�t ~c{�m+E��Ҵ	&-�w`��Q]��b��D���U��ƚ~��s�����:�	`/���r�n�r�?���b@5�&� �\;+�4@�2����a���S����i+�Cp��������2~�x/��	����v���!�Z~JO��4����%;����4��B5���Oi���[�����#��U� �*1�Y�+�B [
i��X��U2n��������6㌶��i�JWD����q2��N=��?�p�ڇ����i6�-���kW؞��n���M7 �h4�^�d�e�Eڔ��Q��>��l��}�:��搞�`�و�����\Cʹ��-�j���:i��C��9�FO��v���SL2�qWio����u���_]!m�Π�ז-E��
�������Up�W@~9ck�Y�޽m#�rb�-��c��3=	���2 ��-U��[Y������ݿ��<̘�t�V;���K�ѷ��W"�{E��M.�o��I�5$��#�V,�㽐��AP��0#�!l6���U��^ �v��qT ���V����&����;��[�&Os[�y3z��..\}８�!5F��ϩ�1ab��2I��~���� &�O#.��y�
����ؓ��+
�i��p�Ҁ��U�4bY}��=_!���z��t� 8/�
kBHΏ/\=*��B 򤫦�:sW��]�Q��� a��� S�+"J1B��ӛX�R2�)�/��ޞk�J���G���ak(��҈h��I==��#v�qǡ���&�bϿ��{M7�M"���>|�]zɅ��-�7�M��N;�0��`����W씋/���e}o��`��.�籑)w�J�DJ���!7qw��d�R�)�rsvC�ҍ4j'-o��1լ�G�ЁfI�؍46�v�.*��7�`_5�hd�Y_OS%�7��F%�]Q���*�`,�䴌E�Qy=z�RI�$�
@�>��"�L��.Lw�wEe���Q叮��W=�6��u �<�����R�΅��c�Y����+�
zg"bm�n�����3%�q�
|�ə�b��&י���Ak������V|�ZZ�ȋד*@�3 ��^[,��D\"%L����QeW���b�{��7}
��ą��{$��/�?Ҿ�h�R�$��Ǩg7Z��퉁8G]&}"-�0 ?�E��"�4Y�%� �&e�MA쾶F߯^ݸ��L�+E�� �"��t�.�.:�$6b��5�fm�����dْ�k���ّ�fg�v�؁-�i��X��"�smE琜��H��x+�ll�<v�R����&V����п�{�E���͏��
�$m�̹���-`,���R��H�ǒ63O7��6�R��%�rp���МH�7�>�ǹ���5��F�s�Z�/�����ˮ���L��e�
��.�q�d�L"C�^ᔀV4�D�b�* ��� yҐ�S�q��h&�N�^{M�ԭ]���←X�/�N��mS� )�-=�-�Z��a����}�i�O��J���	vT�)V�Y��ߡA���ӭT ��Vl���%u�*��n�b�{��u�6�����yR,��O�J�����x͹6���3�"u���|�a[<o��!�Hf>�Y2���h\��@_��j�Y�A�����x��{w�q6t�(�r�6qh�=��ߢm�ۆ<���y�^��K3��Egh�̢�����7D�Q��CY�S��7߷5��;�s F�܇V������Y`�,&-��u����()!X�c�#�ZVZe�0�.Aȟ˶���}fi��=k.�K�=���w+)s�(�Gd�D�h+�e����]��D�����Ϣ)F�}4cAA���(� i#�-��S�.E��YP���}!ۅ��Ƿ� ��	���x�@�)'L�
�(�T�j��(���`�5!�| `p��Z#M_3k�@=@�_�=;��A��x������(<�¾T�^ה�|���*��.���v��Y��V����Ե�"�~ fT����;`WH&횣��j��]�BEE��N	 I?�H2��S��:-����CywЯ�4���EJ�*��.<j�\���l��-6�{
����TH���opTٟ(�����O(�7�#��왳l4���.�ȣ�E���EoߩS��L3�{y}�����,�����;s�#��'�(�������=�V��[Նr���C��#
���_p�@ţ������F^L�~,BB��T6��م���|Q��e|����p������[`��
����VZ��� 4��G9o�]s�4T:+�@9qj�J�qX-9T",�U��x�9�x��lHW���3��VڗY�h�n��I�{R'�iw���T���p
 ���"���N"��FF-5�%T�D����6�>SJC*�US;Ou�T\��}]�r�ːU�����"�`P��Z�B��o%���TK	bo�ەuŤ���v��3����hQ�{�D�%X�$�/3Rա�V�绳�"h5䅆����l=�.��Rg���C�R*BEE������*l�#��"�����5��'��.�ʥhyR2�x'�D��ֶV��-�6[[
i���)�g�S`��V
h��D˰�̀}URꞧ�����k����EC�]>��� ��R8"�Kƫ�`�"�����TG����xN~O�k�u�=RE)]y�=��mv��g�/oZ��k��U6b�hRQ��Ln� Ô��M�x���Ys��b�h5���@c8h|�㕎��
*,�ץhg�k�16Ȅ��(�9��F\z`Z��_�4�T����zZ��4�b�k ,����������f�oc�u���⌓h�mX��������v��WZkS�=���v����������w\�<��C�#��Te��.&Ym���םt{)@�E.�����@k�H�z{��C��s���D����ݒβ˯��>��������� �}�&��A�����ÏYҁc�9��f��O�{o�IC��!m 3��c��7_��]w�56��E�>����f̣��x���S�أ�w�lâeU�� ,� ��o�p�J���d�dӅb	M�9���.�|�����B�P���׎8t_���~o�vg�_|,sk&��j�[�l�[9��9Cm ���0d�՚<!��P:J����7w��>+��a[��뭪�Q��5(��DU���%b��� �J\��-�r�B���y
�$ya�k��3��Vv)si����Z�/�o*�����q���0�����V쨚ֻ����g��)В��*���f�z`*#��*�����P�S�����?;]�/�&?��^=~6�wu%׉)Jn�@��9�*��D,KRj�l�q��FX��mD�Iq _�o�j�o���[i���S����O�o��&w��6J �gA*r�ڌ�3azR�}�(��j"'6��}�@+UbN�0�>G�����o��.9-��~���[qn`SQ�9��V����H�`D1��:Tk�Jps4�4���F�*�#��Ѳ���IR�<�0l�J1��� ��f	hl����)}��)�(�>Eܟ�����mM��d�0���R���ȟE���r�B�	 HU22���1,`M�]��F-��bSt0�q�|9.�H�{w,8�j��@���x����BW��I,]c%���,Ha�F�������8�(���I@����T҃1�\��JZ��IzRl* �s��W5��(�aб$əY,��v�����|U�$�}Χ�T|*����X�H���OT�G�ublY�(�a��Z��	og$=�p]�`��C�lj�<�<=+Ƕ ��.Fƪ�'�[p�q�ک��i�Χ
s"M�l}]$`�^���n�<C�0^c֝��	�G٣����~�֔Sø�IX.��-K=�1�m����9����l[:k��o،x�
 @̢�m���x �,��s�kڽ/�Ĕ��[,��b�1��vE�:b�!�8e׃��[�#�EK�F�]&v�T�6o�X�U��A���=zq�<d���V:,�a[)L\<��$rmd�Y+�X@Zƅ��umX�4j�g��ۆ�h2Z�:P�@[vv�3[��Kn/��4"�< ~6)X�P�}�0�U�a=,_%bn/	�^�_�εIj,�J�U}-坦�BA��_:���jA�{���q�����Ҳ��䌖;8�\V+Z�2��]�~�]z�Ev�Yg�E���?�h�s�;ⰳa���E��W�m�?n{�A�g�~��'��2�3�*CX�,
�
77"���}=m�]{�-v�G�j�����UU50��ۉG�킎ڣ�]u�/���7�/���y��W�W0m[7Q��b���������(���d��ۮ���q�Q�ue��ӹ�km�.�ЃURȓh�{��w�1�#���f-�w��9��i��Ͻ�dE-�*	i�<'X�\[�_��1� �m0�Æ!�"=θ_�v���n�	��m�pذ�N8�B����3����bs�'�`]�x)&�]T���w�a0��wj:�����&��khUWU H�ݧ��.Us�y��?~�	{MmgWx��c��;�\ �������n�����o���A�.,`�����>H��\�.Z�9�KX�孋X��M�!��j�'`�9#�o�1�Z�ϙc�0NW`+J�zU`���_��U��0����Y?W}�"WUmC{H����A�h�G[\I�x�J"�W	?<&\ 1$b�-�v�x�K}v�M�K ���|I"�j�g�iA�sc͓��b�XoT�) ���v���A؏�ЂLN��6�h\!�"�R������h�r�#J��/(�F���f����7l�?�9��:�`��#�CF���s3=sf϶��c:�n��F J�-i/��ݪ�+=J>���l���g�a�ʊq�� ��Aϴ������R[UTh�=%���; �۴rv��>T��v#��h�g�{�V.�i}q`Ǘ�V�T�X�\���I�$�����X�\��ٟw��&��E���x����)�D�~��Xf� &�o	���UA�����W��5���\y)�막�G,T�Yl�2�S5a�]^[[�%{C*k�.��Y��`�+#Q`T���
�31�{s�T��Ӌ>��-!U��*;ژ����<w��1 �L�u�>C�5j 1���%J ��3����q6�FRL��S�J�Rw��r�'��F����I�SN��ڲ�By*e7��s��q�X�]��v > Yu�%���' �]�s�,��m����@-F�����	���;krB��ى'L���;��,��`M;�s����{f�ή��2\� �w�����Y�8�f��h�P��:�V�{��R�:�	7�E�oX��wr�]�14#�m�lX*4�ܺSNZzHC	�@�B'���l�� �ۺy@��9V؞ҫ�S�1 6�|a�f��W��l�Z�$�3������m<'��4I��Vֱ�us���"���+/8�.�������6�
�����8F�2�U1^Z�ҏs���x��*vI�{c�*���ߕ*�"�Qw!)l�k21x:V-��>ȹ�����h<��*j�$�~������e
��J!H(P�vA�@4��$ � 𯂯��x���&� �z<���z�+U�
t^t�yv҉��F�T͟�&؄E��/1��M [XҾyv�E'�C��^~�i;0u6����u�HE���v�����qDbA�|Q��u�����'αSI�o]5���M�@��Ɵ'�|����l���0��՜�T#N��s�/~q6&�I6�9�֛o��{{ t���8]j��~�����ً/��n��V;��������`��{�A���ۧ4g��0;㴓 d�9d"�R,杋��}SK�J5q��(a�}�$���27������c������S�b�/��B��m�,<Z��U�V۰��s�U�f�"��*����P�V�g�3'e��-�����[�hM�V(������_z��F�?�~��~�u������ ��`D��r'�@��F�;���ܝ��C����Lqe�-V|'�A���!MW-ǡ���k5@���O��su>��Kړx�|iJq���y:Ful�9�202��������"�U՛E����Q���H"1�z~B�챢��B�m�գ��#���!}��K��?矎�"��Pp� ���)�]�(���n�����N6���y����RE�Fz��R�������e#��x�鏓��w�e�{����O?c�Oڍ	�PQo�G���;�t-9 ������O�/�pz�#����n7�d:ή��r럓FZ���l�}:s����R�X�Z�P]��Y ��V��h*�K~�Q�ͽ�p�8�*ۖ �J��0��(���ݩ�C��S�PzQ����T�Q�j6W�f�2	�8C�~������Ӹ��D�F𞍔�Ǩ3�W�F�i%`U�!}O̔6��$��Q�%��L@+��T"���:Rz��6���*�df`ݑ�&�m b*���:��M�@�����۫��A��=^
grR�Y�9�_��,+�j��^+�W#T��fC�<���H:Q E�#v*�hT���t���Ha��&�L�_#�Y*`Jn��ԨwK�N�2��ƭ�#t�� 6mQ��4���J|ź2�@D��Սx,5��Z4FEI����D�U:�J57H e��9o<���?��1������=�Q���Kk��F�B��2���w�w?z�.]AZ����9�v�d����ԥ�)D�&Y�_:'i��}�)ۆW\~�UR	��H�yC]�@	�� ���h7��
���t* �`5�f�����@��i��z�$� }��=%�۹��0N	8�W��[�D�'?�@c~i��5_/\i�Ͽl�]w6�ۯ�ז-�o#�!@�' &�/����x_�Q�w�r+��Ums�Kᾉ�3^Le�V��&`$#H����&m����T` �M��&��LGv0�X�D���Yb|�٩�w���C�i��<���vUFI��\r�a�$�1���=?\�4��m�T8ӱ��^�>�����SN����e�w�=���"��Fuplnﰅ��'p�g��׸�a.����]�v�G7Zhq��`>��M����+���#��<Ś�*�sΤCl$?	��]�EO�0��BK���=�0�t���Zc9�5�qŒ���Ѓ��c�*TSy,�}��b[J�ihu�?��K�wI�SO>GлҮ��
�8��-��f#G�X�F�Tl݈��`���I'S�ƶ�R���:�2l�:ú�͜jdl�]\k�6�h�Ԫ��vԑٻ�~�J��HP_E�����R��@ME���c���֒�Kp���k�V�����͏���>��8�Z�>VjiĞ�]é��	�|�N@lg���̏���֥��"��u��'e�`9�2��	�N��őm���-���^��A��4W�9-��洞묻�>� gTT�Z��gM��ތ���qe�:�u���L2	y.�Aw݆�f7`�
��/�{�C��!�;��!x<A��c���a�b�6wJG�π��
�4z�޸�z�F�^K�{>B���B
"����T���'�VL�� ؅i�v�1G8A�ģ�{���O��/9�SU�� lƔs.����|��~���j�5W�Xj������v�
{����Mǁ�c'��9�g_����Ğ05 �H���ފ������.=�`��Y'-�st�H�6�q'h��~/8܌ߎ��ҪM�2��d�Ȕƍ�@U PEc<V���b�� ��j��[fT�I�.�VUU1�_C��y�|�F��mDF:8!���$A~x/+�*1�G?y����2tm��w�RD�z9��NGi�#�M(�DT-!�R�l�0<
��A���43�b�x���c4U��'Ę������iT��s��̝�Z��a�k�3iSH�H�YZ�Y-!��d�ov�18n���'��A'`�9�R9atTs%p^ѼNf}	��(-F��峕�8�o('�G�εS���i�t���O=�}�ŧ6��w��O�&��~�[�H���	�j���[o��ۙ���e�}���5�X�	�XG�/�5m����Վ�D�:�YQ<R���*\`Yq(�b�KS��.6;��H]���*����	�H'�s�j���r�Hr i X��TC5bZ��^�niQ��gC�V�(MD* J��f��0������;��o��~y�v�ͷ#�^��6�,�u�V�=|�Uz�c���	K#]�ʗXU�A�'u_���ǨX0����ΥO_-�7�d�,*�ziʼ�VHL��S������3�\F�r�V��S��a�k�����z���nU��oW,�k����엷�a���:�{���k�)�h,_c��=ns%�(���z�i�%Xl���2���|+�b��qV4}9����\y�Y���?B�QO=��Cn	3���MXG̷��T�"����t�O߂���/�;H$�p�	�yk���X������Kv�-7��)S������/����UI{�}<}�]w����ޞ|�
������U��H�4<����I���y}��_aR`|{��J�VðVV�ڵ7\o'�x</���/�ܦ��}1s6F���?��F�n��8��:�Yo�A��e\�Qb�i��u���\*U;l�`\�HIg��IA��)8#bd|���;����폲a��wȍ���j����6!�U*8l#�^ �/?v����{i�0������PIRD֨�LǑA3e}|�)�����K�Q�����ƃ�p����j�K[܉��~/�"�uXֻŰY5읅�0>tI*�͏D���
��	Tj�혂k�Ԛ�IV��n��.xOd���D$��`�5a�:�н

p�}�v�\�	�;@�vb噿zRWՂ��W��ڤA���S���,��B*$�0ͬ(ڀ֧������F�6D�3gη^z���1v&�1	�?�PE�U-i�ar�y�� �9�F��\9f4f��3&.�t��T �b�n���@m*'�iO?�[[�f��}�iv�A�/o~�`�Kd"//�e�j X :�X4�K}�Z(�T�2O�T��)@iE��j0Kpj#�L7��4+�vE����HM�@�543h��a�,����5�^-��<�kb�R����D��h��6S���D�Z�$��E�P�Ţ5�ZNn�k���PmG���b(aX�d�X�l;)i���4�HE}f���1`��`��}��r�Riป97�a��ɛ�s	�	jA�x���%����{�*O���G�$��tX6�e�/�2�h����|(`�B :N�L(fa6P����o�ㄇ,-�	�X�BRO����[��e��GM�m��u��Q_�|���7-�E�G���cW��"� ��Z����}�t�r+iO�������"����lO|��L��O>bmD �H���_i�b��Gp/k �ju�0���$�'pa^m(��M�I�C��4�R�.V����`��ķc��X�2�r '���P�?]��ZL&�����5:h��{3@S��0� �H��tF���$n��ɹ��2Sa���F4#t�Lζ�W����]��{n�_�q/����iVzZ2I>o��#Q�u�]��I�Eh�a��ꤧ$��@�
����4����[cMi�&�-�:(5/*�4%���6-Ji�����G[������x���=��u��>Wv�$7�G4�l�ҕv�5Wځ�^`����r2읏����k����j���Cl ��c�ؑA(�����f�=��oN��{귶�!��6ɐ��߿f^��ؙ�_�v.z�%�[�{ˎ�z����g�׸�6x�AVEE��J6��٫ʹ�o��S����=l����_��]w�MV��ڷj�T`�1���Ek���o���N��`��!cwE�mG{�-��bQm�,\jGy3>�_�������n=st>z���Q{���������a��x��%|����s�T8eڤ�����ٳfyۣE��Q�o�=��kT�b՟4�VfITeJ#YmK�["�_�T���|U!y�V1
��g�d  �N��s��v�=��L���-��OI�tu��[�Iͬ5\�nS�T
A���|hN��~R���<��$!:Ԭ݁O�}��$=���^Z����J#&]i�4�h3%�W�����H����,S��+Ū5G-��I;J'ُ4oL*�� ��K���X�����5�>� }�b*cXi�%�g)��K���$��#�,f�C�><�Ćz294�� az��`���Z�C�/]�D����c�]t�x6��6��e'�k�~��x+�E��A�N�f_��9�9݈�ζ'֞z���� 1lP�^>A���_�JJ��-.1�KL������~`�V	Cv�%�8(��1��o �r���Z�������s���O��3��Drӈ̸I�De|>Ͼ��=_JT
�����PA �F��S�=�=�:�WT�F����J,���6�@ЬF�64/�z�����%ߺ@u�I.f�V�dO>�:�6��4a7������|�@�KX�nGs������~�h.���?`??q��	�5�[B��]�ì|�jgI��8D��y� ��9D%K/�3�޽{�$�*|�Wn�E,�����>�{��lsW��4�V5V5�|���rC�u�V�!�Ԯ�D�*ؐ��XG)w�)�S`{M�Ֆ,\f�P�ɦ�mو�cx�6w���Y d��������`gx�Ԝ�\�D�f5[���n�J�T$}S�|��lPcF�f�AQK�v�QC%���[
��d�2W~X��5��fc��bt���G�@���Ӟ��'n���sϱ#��H�6��I�EǞ��ާԪ�l$����@�#�g@��I�Q��>ClZ��6� ��i�d�yC���Z��:Z�D*��+�����,�l�)U���_&���k����&�gK�Th��N�Sa������6�R���B�Ű�.��V��^,I�3}���,��:{��������k*�6z��N�>�@�����Z cW�"[}{s��Ti���u�s%��ƨ����2zj�S��t�KJĒ�TPYGjC_��ņH���3D�b"ܪ�t����F�F��������l؅���JLu7�M7_g{���t�i�l���(��.'����v����o��0�k쐃���K����5����������+n����p�?Ӗ/�;mۖ�g'�r����=���ŵ��ggq����Ξx�M;�R�j@�w*���du��14 ݃�(��A��kٯ�k�(��Tzs1nm��|���ѐEڕw=c{�9���f����S���T	׵���ޞA��F����i����H���)Ě�p�m&UK��.��)��x�^���N`ml%X\�zp������ʿ�~{��W�f�|4ґ�l������h��r��2
I")dj�/#��o�X%�
 Jc�H	C��>@��@@\���."�7_��s��G˴[U�J�0��^2���l�	�V,"�����_g]Y�	��@�~4�����K/�H�+�FZ�F���W}��ib��3��rCs.x� �h�PvHY���vR��>H�!�>?7/Q�	����)-�/%\U&<�ݦf��6!�TLI$�o�s!��k���i\�B���2���L?���;h��(�BkrbR?+��#��r��K���tTl����s��dЕ���,�}��#��k�=��{�%떗j��;����_m֧Ӭ'�Q�]tB��ҟ�Ąδӎ?���?��CO��Jp�"<��m��a���䒥Kp�.��=�Fуl��Ŷq�R+�
M�i�ī�4܋^�ۨ`{���m��	�w�MT�I�˦�tf��/�'�)JX��@yQ��@�4Rhju��&!�/->QxըѶ�w��6OL7]�q5� oUe���L��c{{�1�����m6h�ۍ�h�M�l0m�.��rO��s�Qh��l{���
e ��`�h"=jxwOS���g#���aC�+k�:н�"���S�/g/���&Y<Z>1�`���0�T�A�4n�}��bm�Î��M!}���l��Mv��'�K��Ӯ��dа� ���o���Lg��tR��B�gQ��D6��6l>R�F��1����c��A���?�����(5�'��C쮻�1x��3Iq"��ޝ6�JZJp/���L��(MT���$�{�Ek{�
� �0'��"l� �%��M���Y�*����,RdlPQ|���ۤI��w���.8�D��P������}4�-��4�k*U`���]y�E0�%�+��m��/��f�L�R9�F�o1��4wF�E�k{��"����~/�(�g��)P�%�&J4���@U�m�ɩ������P����R#e1Ҳ�P�Qcc-�&) �<�+I�*�~����q#.A ���2�7�-T٥��)@�T�Aq\*�o0F������\iד���6�u�m ��ͅ��KC��>C�P_)D`�[*szy����ʼQ��Ӻ�5b�b�0�Q��|����t`)�6g�*���G�1m�`��`̵��rR)�Z
#�(�S$b��1��VvN�(���{G�o��6�vyE��a�մ�����3β�>�fu��|��T}��⅋m5��X��# 4/��!��w8g�J~>�L�K!ȇ_�&5MJ���|��?�ƍo��E4oc�Ap 8����]��Ƿ��̽6�����񬕖�)n��⒍���a�>�R�6�sO��OZo��{�Iv����Wh�ҩ.�F��+��'0�jI�Ŭ�x�-,��^�
��y����k�ϼ��-�@��{єC #��a��&��H�yM�2�>��3X��v���>���ll�:����[��+���Z,Z2s�]��e[���d;������lX�d�_�/j�R���AQ�V��c�E���dj�W�w�W�&VZI	ī`o�up�yH����b�~�:�'q�$H���xV��g� $�4�1���Ӥ9����t�xHϤ5P��`�K�^���:o @�'z~�s����p�d�/	��lT ԡ��4y ��x� �Uב$�N1�bK#��8�,���;���*gօh]3�`���b5,���޵B�z�
{���ޚ��*��:���R?*�j��������&�%Y��h"L�����s����8��S�лa�K~6�@/�#63���.B�.R$6Q�|�i)�1�ʏ#�J)����5�m�9v�1�Z!�ۯ`7\~��Y��~�;��W_m�;�*2N���_}e�@������tXՓ�T96��N:�h;�ʡ�_z�V-\b=qI^^���m���L��v���n����4�]�t���x@�7T��&���dӚ��m����lkM������]v����2E�����(>)g�b,:ތ4���kۈ�7�L�U
sO�9�VȽ�T[�|�H��Pb��L*�d� k�A�*+I������[}�
�g�vM��Ƞ1�8"�1���ڝ�~�\;ɢ>ƒ�n���h԰OX��f}��]�����%��UT>��\dǝr���,�) �dK�D��UقN'�XMno �5ڋ�����ťv���m�E��g��w�!ف�-��^�����(�ED|�=;���[OsblkQ�h�ꑇ�6(�8��S�^D��u�zwV����@VI�6;��cm��U�g�O��w�nD�G������KP����H�%���ߵ�]
 B�J���֩L�`��U]����nE�@� =���Y����G�ib= Z�޲!��+Ɠ���Ƶ{���)�ȷ�$���{5�ZqU��q�IS�b�7Z >&}$�ht��!�B	m�*J�b��gM,���)
ۍ�:�ͳ�^L�6m,  �x����J%(R�$:�Ġs�F�-�0F�C.���!pwY���X�t�I�'0>շ��tl]#Z���ؔb w��Ϻd�J��L|�I��K���p:�֮T ����ٰĮ����+N����n��6X�6x���l��lu �V@p<��]̃&�������-���`�![��-0Ǥ�i����h�54��I�.[����>�vcs:s��r5��ֆ�CUE���GQK)Z�ml�Z��9g�S�P�8����}�B˩�A,�1�p!���x$�-W`��R2�f�J�`��
}�7���S%x����;_Z_�N�;�>~g��~�͜[@�b	�PA��2�t�-�{)�*{�_1�s �q6�
��$�4vw�����~��F�ʙN�sU�w��F�MrW*
7Pp"��d��Ё�3�i޺a#��
P�E��yO��^k�^|A� [�%P5��
�~5%౹��J���.f��0�,�I����
�C��f��Hw�-6Y�,m���0�4o�'���lj�-��Ӄu��r�;��9&�6��R�S`��q�N���V�	6ʮ{� ��ֳ�]T�n�ֆ�$P] ��t=���=(���NBZ3����|D���2�`��=�N
���(8Lb=�v�?��!���a�z������?��k�v �� ��d��84�1�e���f�N�S�7^5)���	ĈM�#J�3jl�S�x�-AT��z;����"9zF椌£	��d��\�A���:�fUr@v$=�a�����-��؆�a߷�Q����kՖL�R�BR��\� �7�[q|�����W\�k��%'�D1�$�~B����;+�Yj����#Z�M���3�j|�ۀtὢ��1ѝ��£9��/�l�k�	D�kIe\�����L�I�j�/���f�^;���m5��@�-��W]�~:�Ǎ�,�ܾ��];`MT_���Y�˘M�}>S��i6t�A��A
��}�����o�IG��Q�}�Aእ����h�'�Qf'�v�M?�����-$�5g�3F}����ju1e�[鵶���6D�����ޤ�u0 o,V����`�J{�JX�x��a0j�>��CB�6OUC���ƅߵe"]w�F�7p4�	a!���j�1�;a["��>^en�����4��OCw��i�M�mw�h�RH%���>h�\t�y��G���/.V�l%e����[ia�}���v�a~��fX	�8��cc���,��?�nd�.v�n�n��{f��M���e���u˗b��M9�k�o�����E�g	�G�Rc���_���=�7��{s]'R�چn�7�F>=��F��t6f��a ��BP��S�*N�0��ާG�L[���>~�M?f��t�n�7k�|X�"ۊ�d����3�}��PDQ�(��n+6��L�f�ڵ�ˀOы@�b�F���1㕏��T	�k��ױ����F&�����3{�o�>X� ?�毨�	�X�a��"E�q�Z{��o�GMj��M�E�#,4��=�>��ٶ�_/B#i
=��T�f[!��D�j�S7�.�O^j�rq�Qlk��dSQ���Z����*H�Hma�أT�9����%p�"ש�3F�Xu-J�H7�EU�B#�ɠ��
ғѰj`�����7D�Jg�ôH�����j�F5��X�����W���O�خ��*R�k���YJ
;�2�E�߿&�,�$�,Ҳ� #@(�/W�k!Ut)FK:K�3Ԇ�Lb)L�
: XU�bS��(�١���#�)�����#Lw�	x�7��@��.X
���Jk�֦��镡�wJ��sk�*���K����&:\\{�6��ÓN?���_aç`k�p]c4�-!��y��8���o�笊&���;�'��I�s���yl#��@����͜5�VG�X!3Z_�y���Jo�����~u��̛�����L�׺Q��=?��T�
���kbNn�DQ����k�TU���;�u�{@&�-���x��3��/�H�[��ecñ�y��uآ��X+l+slނ�6��v4L�FZ��5�O��&�a��5h��!�.C"��g�I�o����k��]�f����tL��@�$i�ҕ6��i�ZN�|��is�.�9U��DK�z�1��*|bS�w��So��j���;9���o��<�15����c�$�U�%&�C,�Xr���q����R��n &Io��Wxn�5/��&�A؎���s�< �ҿJ(�|j	��a;�Q�4�	��X���{P���醄����s�_@����cpv�;���,���EV�?Q)H�����9����죣���s��/����~-�o�b��a���=�9x�����(N-��G��a�C��kcq���E��'bvƵ���-/�r����W�d������*�w>�N:���z�����N�%˖�GT�2i�I�Ԍ���X(��iY����g&BL���YH�~�0�o��D���5�`�s���`�}&ᚼ�a�1��S��y#�fˣ2�&`%��ʚ����B#���Қk؀Ri��v���=�p���jy�x�D�˘���q�D����# Ry��ɠ|R�Yԧ�m���2�c���H�t��kl���$6$�Gr.�P�	�D�֍�Q��tfm\\�e�@��믳�=�~��K�{,;���d}HՖoJ���S:!	���T l�����&�u���x�m�Բ��͔ɷ�1?`�}8w�Iz�A��V���}lS�&�@Ñ@j��l3�y@_��������rrY>Ҷ�^�a!T)��5,����d!�mdҕ�fS'�?E D=���M���C5�r*�5�ˁ��l��z{��:��b���_���i��b߮f�)����ɉ�{�E(�/�	{���p�'@"&D� bT�n��y�WU� �����|�z�ȵ�m���jM���ʆ�'��� ���y�˘e��0��z38;�~� �\,>���M ��I��8^El4�&%Czۺ�3��	���oEs];E�K�̢��'!���t�J˩Pé{E�P���TS�(U�V�_hT��k� ���@�S4GzZV'-,��?�H� ӓM۬v��Jt�1�J=�5��I�>��7���δ{����[��a��m���+��F�JxA��X�$�r��I~>V���Q�Z�	S�:�.�I)�x�7�R�L@c�d��ޠ{�0$�	�T�$0&��D݁6h���wf!ܰ��~����JŨ% _LP�� U�Izl#i�s�>��<�p{�����A���R: lM�}�L�m��`!���[7P��Fl0@�&�!`�7�"*��Fs�h�9~� ,��&���zp�(�PldՖ�=�.�~%61�H�)e�7���s<��Oe� ��٣���UT!��V�u�J��fb�(}��u�	�A�J��LQD���*�{;s*���q�h�jr�e�R��6g��T%�:�!6Rl0c��I�m�Jk�!�/��lZ��`�6mX�ܢ[	��r@M'�5�-g�gX���m���N�����SU5LK"�kbZ7�h�����GTS�ܳG:L,��Ҏ��
ir�V���~�S���G�9�W>B+�@��)_ނ5��Z� \^��VC"R���Ä�!K���"V���h��s���*�E70�F��
��KC')��� Sҧ	��N�
)%g����Xt�� ���/C9"�{��)wD�3�/=�{(Y������@�0���;����A�59}m��*�[����e�@�?�����K�ѹ��h#���Li,�2�_���۽�e%��PM6�N>�p��"Ӏ�v��c1�,-ނ(��}������/�i_/�3N: &�Ke����6��u��|9w..�=mظq���_|f_t��1j�-�l������s�`X������9������u�������~y�S��{؈ѷP���=��S6d�X���+O�-���� 2;�<Hc ��� JZ$��Ĩ�:ЅD�s���&΍i%"�T�"�(R|��h�0ll���B4�ܯ｝�[�pz��CT��_ �L���އ߽�vloD���~�oh�r۴t�%�*
`G��Q�ؤ*H�a��wᒥV\^����'�ıCmԐ+AT�n�2�;�t���K�ٜa���k2�X��|�I)��/N�k����T0�ƽ��4�\��?�	�a7�L *F�R���&�-[}�Q�Oڷ��Qi	C7��TR	�5�;d�8z6�v{���Ï�ɓv�{���P���k�؜��{c����[K(R�b�����R���-��E&�~-�K���D ҩ�ѽi�t�E��9�F�b�d$-�R�IA{l�w��v��{xQH#��)�,,d
WR���
�V��2J��o�jL��9 �QQ'�)ZHHZ���/M��*>c��Ú 1�O������]�(~8��bH�I�w�1�`S�o�Mǵ�^�p�2�b�\E��b�3\Ţ��ǛD���ac`/ [H�F#HMGs���F��,�˒ e-j��L'��z�F���C�������������4]n�'0_R�V��YpU��H��z;�K y7)���%�v�m��#�$Ԍ70�kQ����ۿ?�b�ך�JJ�xf�K$ *#�<@>[��p%�w-%~���T��.��Pz!���1��rr������g�5�_�I��v믟������n<3�V-Y�UV2	mh6P��t�B�����B�dSJ#ş��K��"�ZvmX�z�����v�k[8?�|��b���ǎ�u
א���Bc<�������~�؏��8�k��s�a�Q�_+���H`���)��z��
b��=�x�=���C�3��OQ��5��a�F��ǁ�U���.���2�B�u"��6ƛ*�a��Gs=~bٌ�ރ�`�=��GE�s�����VJ�M��lKo%`�~��!k��cmf<%qb��Ȃ�M
�nk�I�1�kU��\��";#0��t`\�� (Z��?�+l�W?>���K���O(q`pм�bR
�e
/\G;�0�
��v_��.B��&^|)%�uFsG�_zh�!�|W��B����7���Joh0�ס!K\��G�������ދqt�(\Y9��@�<�Ą����
��?�_�P�:l���ZE �bC�z�a�����D��UD��AX��RR�,�j+P�|�İ��P�?�y�]u-,VΣ�ثv�ٗ��Q�\�~��^`=q��M��p�)�U%䀫��/i[��^����Kβ�����>���|��T�nGy,�0��>#͘j'{��MUe^6}�^z�yؤ|=�p��|��N����Ge�t��>��ݿyQ/@�.T!���@����;�S'�m7d���ؗ ���4F-��O\L�,d��-����ֺ��H��46m��Z�ۘ��!����ʣ
l"Z{��8_x�@�&�`�Ja*۶ō<ǐ&햎��E�̓O�t{���{9���>hd�'�"B�$83��s�>H׮_���^l黖��c�v�@ϣ�f%� 1��� ���'�'�mMұ~h�f_~���K�D5��y9V,�j��:�v�u�7�]��Ҿ�����⡉���c��3����M��=,"�ؔ�1�Kgq��R��ʆ�]����W_�%�����O=�;���Z��!n_4����3�,�5kI}u�2�b�SP�t-�*�CiK��ZZ4�T�Zc%Bw)�B�G�V3��`�T��� 5���RI��0B-��[�nF��;�6`p8��1�0ɲE���v`�K��"�QŌg�]i
�a���#�鰀�;�Z���Ͷ�XՀ�y4-Ja��M�2�� ��ds��]�'�D�+��8�^�#ِ�ɛ�j1+��o�.[��`m�Đ��͐k>f�l�s�R�P����T����[I=ʛ.��V��4:ITq퓲��(�`7R9��;/�[�������a���qM�HC'#o̩��zҮE�J�#L L����Ѣ�`���"�L��e! ��Fsy��\��K���F�(X~v2�)�5�a�׆+�=� ������.��~	�����betK�� �E�z�y��#�;�.��.{m�7֫�p�f��I���gut�Ʃ�T/�2���%�����fs���"˨�V�h�3V���-E� �D?��Ӱ]�W�m�s��D��7UPd
e��x��
Vo� ��!_�d�O'bC�!]��xEY��t��n��k�K�S �r}ԎJ^�jE�`��<zE^���X�QE	�j����*���:l���b�`���r܃G�}!�!�h��rR�d�iʠ0���$)�(�*�:գaL�M�	,m�H_�iV�p�F��:I0�k�p6���}�#�8@F=�BNT7��2ΊI�j܄��%��v:$��myG��Gv���wbK����Q�_&��� 8c+^������[���P������/&ȨXI)�pu��
����A@)v]��|�]R���ސ<��1�앋��%�s0i���w���h��/%t
�)��uZ�ΎAg�˥sT ��� ��T�_��W��F�9x��;�g!�K,��%�1�&��q���Qϗ����&���tw%QQ�D��|�+��'�D��je�=��-�|9����� �������n]��ҺѼ���v(͘*������H�$t�� �ڻ％�R9Me���;	��v��l����z����쐾�?�3J��4#N"$�Z�����l��q��#;�d<�~m�<���\��.Z� �4?To%�.�ZY�jZ{$��ś�3���1���L2S�'��yʨZZl��j �����	s=��*�ECT�ŀ;���lO�����!9r6!�)�':'� dZn�^�w����Pr�H;A�� �QC�[�K/t6!O'S,0 	R
'�tl��\-�D<��9z��s�(f����}�^��f�/����@�e�GJ�Ϡ\�p�٤����C��4�޻���;��Yw��M����7q�?����3^�B@�zhQѢ>�b-bYd�ISճp�!v )߾����IJ��ݎ:�  �qnP��o�,������.����4��������o��0��uQ�W�����x����G�FqCVj�M q'׍�a��*��O���	�UAZ�b�ʦ֧�`�?o�}E5nLӴ��l��]������1p9��f>/F��uZ�&��0�y�u�z�7�BvY���x6�t*T�6�%�S�n��=U��h1^<�~W:����TYԦ�Ř�� ���Į)��H2�R����r�br�' �hbĘ�G���&��D/1V�x�	%ȝZ3Qs��z؉��I���EHGL
��
���*��x<]q������w��~u�=�e�rR_I�I�:*�}�c�´J$�"��$��zgR�)��R!H3�+�O���X#�a4�i�B*�*���3��t�ο���c:�3lgC L��H0� ��N���
X�ft����v�9�څW�^x۲v�@ss�&��0�I�λ��U�gb>+�����V�w���V��ؖ-^c9��'7s�I����_y����"��DZO��dK'���Q��7i�b��o5�sb;\�;*-\��ݷ߲լ�Ih�:Y�eP9�J�QTZvI�- �y֣�k�Gab)??M�>'�����۴�H���%R�O�h%3y�گ��]mMH)��#b05��8�/��a��.�uXAB���\ˣ4o�U�\�H�m�
+�)/rBz��?F�h+م6�-��-	߼H��&λ�����J�[���zJz���_� �^��˖,�
b���%��ߩC���@��	`
��?��߃|Z�BvT�n�Z|B���)`��TZAVk ��P���	&;�o0ag�+��l��@^�<v��}�=�#*p��_ Ek�]�� C��%��-2�U1]��\� h��~�.e4�^�jF�K�X빧-}�E����?k珜��T��/�f-X�ws���O��B�pRd+���B��a>l���pvư���� ��O"yRSMT�]��;v����᧥ػ��M���͚0�M�E�����zC�d-�T���ƹ���D6��(�B.Y��q��{�a�-U>I9}�4L�u���ϐq�«�8��<�^�E�ae��\G�}�ֵ�V����dL_{�	��7��)S�k�JN�u8��-]��N��f��qv�u��K�~���8�� D�W����^QmͤM�.�Rr��w�\vIKyE���a2D��+�l)�
��b�P�� "]�l+���M��lК �QJ%5�i�f5gՅ>�&\�{ JOC�0l�`�E�o�7sl��],DMl�F�å�'��ISM	dm��^��D�^MF���E��I{�7��}���v�m�}��W֕�P�L�m[��V���j�f���ئu��B['mO�������Fr��C?iq��[< ��	���0� ���!}����\��>��k6P�<�t��JkQw�a��^VD�Y��3ٔz���=?���JVx+"EDi*%�	�v��ꢒu;�c���)��	s%�3���),�A���ːF�j	��V��Ru� �#=�vՋ�1�R�����9)R!̂J���%>�b� �ӡ��F�t�hL�I�C�:�ש4�W�a(��)k�� =ќ�v=Kh<���G�Ot��<�}�\���" d.T���X6٢�=�![��D�P1����`]���8"�f�Rfi�aj �*_��J����҉A��V,������6����{��k.9�n��z{��g3m��V,�4�CU�~�5�jZ*]�����H���$��h]e�@b�J�j�&e�e�ݿY �]�Oh.�R
S`������c2}����g��X�+�S1!����Pb Be����N�{��b�dv[p?�+�ĳO��a{��Y��]D0[V'��
�$��^e3��<U�Y ���z�E���������/s洆tp#��=�6���J���1	��RR;(��j
+js	J������P��[�f+(��6L)�X��4�w��B�#��**���J_�*c�hX��c�(�.][m�K�O��7~<����5�&�� �x�G��
��S�X�(��Gr�߻ OUV7J���LK�V��2Jd` ����j��(��)�����u�_�l�<�l�J=�Rf(�_WcL�jf]�gF�h�5�k��lf�Ic�~�?�\�f��?��t�܉���T�i<�s�
:�I㫲^>|.���|���{�^���YA1�z����� �0��ф�����b\�\���h�;��{Jj�S`��wJ���\c]E�9���gX,��l5���ź�c�&�uN����&�~Ҵ������A�7�� ];"ؤGv��|���*�¹a\��z�='���0�U���"��R^6���I��D��P��,H�#pN�\l����':���^�f�cV"�\8_�2��)��=��C���~9�& ��K��8;���H���\ĝxs?qW{�wm��%T3��o����)���c�P!D#�����Z��H/������O��=�^Ɨg$��W^{9��f��(�����g�Fd�j��N���>�s-�"�R66�|Lc���|'�������b�
UI�	y"�z+rVC�V�(��B���'���b����7�>�c��{�n�,�֬Z�q� �G�ȨQ�h\�����0sgϲl4���>�)[�+��+Ɩ��(}�w�Wy��Ḅ6�_[�}Gme't�(k �5�&���>��+{�/�T*��2��ƍe�`����H�"��|��U�5�w g��T^��q�Dn���v�u��s VMZOTqײ���.����5�M�]K�Hs��8�lP�-,�T��%U\�Dj���<pb��7 ����l_�M�C/#�n8d���|B�YJI5�8%�[6C�+�`��C3��q�D�=�lHD`$zfQ��������m�L[��\[�?������T�l���HϦR��@T����N�J��R�i,x�� %����z����v-"�b	 �_0���^�,�=��{��wi�r�j��E�{��f���&#�������s��,&%�eY �
��VXs��Pׂ��D�fZ:��**͢C�RE
D�$��l�Ǥ@@jJ�u���Ѧ��۟�[�;�n��z�㶻l1�|C���԰,&�	����
Ed��OzY:/�e�v!�5� ���t5*��B+�G�Fx�e#��*,�%�=�D��OY�M��`º]�pJ*�����B� ^5s/ W�3�ڋI�U�Xct�M��^jǞxkN���'�o�� � \��oZAw����*�>%@�&�Ɔ�x�b��� �y�DC�>��ͤ!��I�ɰ��`|��;(��q�"���Q|N���g�{�H�bPOe�U��D�NUt�s�'R�jeV	`�����#�D���)�Ny�q�2�Z�{ռ�:�j�rc�3��d2bY��g�����i��R\Ws��[h��J�8�1_��S�s�����=�gB|h�+ %�XR/�6*/��"��*Q^�*Y C=!c�F�E):�2��s:[�(aċ�3RY�;X;�#-�r��
�5e��^����_�`�ʹڼ�I�Qx�ipO{���0��B���?/�ґ�h�c��ĕd�jHck|gQa/`�/���@b�B:�p�O��8UA�5��V����gIB��ּP��� �к�@Y�s>�K�M^�n�Jv��q�94�i�8F���b�>�w��]P������7LN��4N��� ��9��a=�
|��W��b��%x��y�)M���\�ycL>�A(ݝ?�q��t�u��W�yT��meYm	ٖ9j/{�F�}~�]y�h;`m6Xn:�+t3�b�x"�T��
�#Y�.c���Hդ�9-�\*}�`��c,�o��=��TT�!cX@@�YV�9��v�A�l�C�/q�~��S�^�iĳN=Q����' 0�m<�N!��^v��{̳�:�'�aӦ�%J�`��y��c����{�.��R[�|�ec����d*��6��^CG[i�@I؜��I�I��J5I�\�`k�uK�$���»�{�Et�sۍJE5�^Cۥ�>+Dt��?p����]l���>H-Z�F��j�[T�ewؼ�i�F������E45�&�S���#FGwi�W"���f*1Ȥ�P�@����N�l��w�8���h�Sw�c�՗cp�&�z�T��ʷB&S<��D�|��RS=v�^�Z��7ifMZ�أ��g��$
 MSTN	G-��zVzPa�x�\+ް܎>�8��1����9W�&��_IrIV'��6��5�@kV����,�9|!-�F�qjV��&!��Zn-�^>��k0�l����I�#�Ah{�b4���o�Z����*{%���C����-�+=���@�B��^~�֐�UJ�3���f��p��h��7F�f�P4�z�56C�NLr�	�n,G�|�"9�H̍T�X�B �.���WgQC�w"�c;(����`�g�RlE��6����$c���b���~�'�i��d�=��I���8� ��YT�f��dPņs=��d�Y���mlj�t�P!J%�u�jRF7T;�е��~��������}v�w�*,N����*�V�@��]ڎ��D��ס�R���d�/�Ռ+��i��9P���MC<l)'���`���� ��g
UI����)����cz�3�bh�jäjY-��l %�U�_y��C�[�/��g��s �3 M��tti�b6ł���J�Ƀ�H�k��}��S�/&B�bc�M0�c�n�L��z4�!y�c��a�;���IG��Z�=��f��Jf�ɐS�ҳ����6i�4�^*�t^�8z����5�8�f��U�I������M�)��:l��G��T�NHl�t��hx���mހ),iJz��ȬWv#�l���f�� hS%��{M%�Ĉ�����d�s߻d���jRұ���pȼ�H}NL$�1@1�`R�K���p� �f�>�ϖ��;/B�ݳ�K:4��Q ��y���&�S@ꟁ�����)���zߟ`;�H?����v�S���i��$-��:P<��
z$�ٙ��9 �y��κ�����@�<$(n	4�M��� �ʖL����a�*�����|I�#���?��&�R�<�v�HT��k� ��[}}��Ȧ9f�^��X��tI]�p�5��wp�:��Np�,{�5�W�=̐y�}P��L\�\:��P	j{��T���g��@+!��v��	�%�Sd_�.,:UƔZ꽟}�h���fG�3��O�����6u��6h�.V]�N%6VH��#��	��{LOr�{{�؏��I�����|�^}��<�ʢ/ˈz�|�|0�D�r�ޖޫ��������k�����b/����y�=�B�*5���A��֫m�^���״	�{X�_�x#�7=�R��n��fZ	�i�+�̳�d�]y�	V�V��w>�o+�1�}�����7��׭Xe�,P)� �djNc��f�Ă,a8�����T� )mۓn Z�caw���*J�a�X<s��3(�a���H0pW`�)�O�yvRo����{UW�����B�x�4�^�r6e�һ����7*!�^�a��Ɛj����Dw+��hyH1y�H1��'"@^�b�m"�_W��'�� �����偤����x$�'o��0c�a�ʩ����^O�Ro�� ��I�0T�[���)��@�uk=E}���[p=&��h�:��*�,ޮS���̊��2hf�A����p_f1���
��F���Z�3`b�N��Z1��{ɮ��h����e�qJDyo�3��pޝ��T"���a�|��/>��*.Mpti\[�dױ��Q��L���У; "l0�\_�9�! L?¼G�}�t*H�\M�@`���~��4���C�S����pgp�O>b�%6��Q���<� �f�J��[o*��%-�.�/�BZ9�6����XcqjՎ��R�nm�5�Ẁ�$U�d�{��m7�e��v���;lźU6��Km���sT�l�HJ��`)$5����,��& �O�Ո�Iz�l�`� _�
�eU��ґ�	x���ᒯUѵ#� _a�KxS	_��D�|�@�v������J���|����:��D��}o[G����o!6� )�W,2
�� �}�Gv(=R�`��z��^�S���X�V�a��n��q��2����(M%}��D-�Z濫��Gk�*&��$�&`���*�Pu-c��LvE���� �E}����'��Ŵq��YӇ�ڤ�=lԀL���JZ�|��kQ-������o�\QD`�И�+��4�kK�z"��E�)�@��ӎ#�K �:��ȠP{	
��a̼v�V����(Z}a����� �Xq�%RUh���!k)Zdd�AɄf6���4�~&i`�����L�0!�"0�\3����N�*~���t䏾N�����=��9^#�)h��K2s�0�;u�i�|vP~�w�^� ����w�T��U�҇���sk�����.X.������_�L/ml�T5d � '"f�7Xw>k1��H���8PQ1����^��Ќ���������y��K�+�O��������A�TP��;�����;�!a�����A� �[�������O:6�HE���D�����{�G-��D�M�5�	�͟m�歵C����
g�"��h��8h_� �Z[l&R�ܱ��N�٨6\���b_�]n�/[k]Dኵ6�k0^BP&�s�Nc��a��ڍw\eil�ň�_y�C���-��`��+o�"��8R��e+�X�u*�Τ
�=B����O"`O� �h7a���7٤=�e�N��܋|yd�"l�,ҕ�F�H���?f6D~�ܱ���>�H��"@Wı��'��J�>r�͡?^7N���4��I�*����NϗF'����ق%�hX ��#-�f˙� ���T��&!��]��!�����s ���ټ��$�J���)�"� -�k3d�`ҋ�����7�F�5h�XP{���QM�h- f�7�����h,d�P�P�i�oj&��fV���PMc!��-��w�,�QR�kc,��ú�����=����7aWl2j9�t+�&`t0�'��2��7�4c%�U�U PUI��6z����ʎ��f|蚹�)	h�rO�\�Y(Z JQf�g�S�k[�p�6z� ��o�|��G
��p��q��������{��S��h�� �jb���f��Z	�������'����[9��*�G8�6X�xBe�ZfT��E �X�e<}3UeqlΩ�W[( �8j���O47ر��A[�������F@%��RBQ�A_��B��c*�*
����HY`�	W`�NLȲU�ev˽O�7��Ե��ch0����"J:3E��q51�?\'5��$�)�L)�u]g%�1�����$nL��4"'���i�&��a���S�;��w����4U� �4Z��Xi�/��&M�j���y�J�޻L�O+\u�h&����t33��&���U�t�H��0C���x�KS)�����_>6��a����K�'VM�ҽ_�]D��r�*��>��Q�01�Ƒʸ߈�_����./�X s)���� C��&����zR��lP���R,׷0���ֆ$�=c���׫��iA�W�hd���%��+�"�'5���1��0�V�) �^D���ͣ=�lK����z����6`��J*��1�q1d��w�4&��N�'���-�
�>tN����S:�_�%�W���ccԿ�hh̸~bK�}S���.������c�p�P1�? (5��`M�5�*���ꫨ�zҒ�@��sOQ��0��L�t�2i�~��a������\2T�{�nOJ/&�ƿ�Z?ǀ�
��g�?���r�.|;Z�is�~�3do�T(�<���5�����l �"�]h,�w-�q�o/����[9�*��>C�����a�`�ʡ��`P�����es�-+�<lb�7.��&dw�S5��z��#.>_��E�
n�9��0��8�6i��ؘ�|�/�_᧳��@,! �?�KR� �=�:��-���|�1Hn�w��J߲gqsoZ���6� @���73�����Y�-n����{$�v�I,bf��q��|������L��_��J˖��[з,Y�ή��&@� �2u����������=�һ�-J5�9��Cg�v)�\�_o�}6�―4�C��TE��n��t7�{Y�a��,�14�nbsL"�	��/"	�Ŗm���&��]b���K��|��W�<in"�.��2ٰa 
Yk$at�6L�'�}m#w�ŎD�R�.��Z@G���W�H����Zk���嶀VF��M������6=�	�O����%��N{zV��a/$:��+�����̕rI�U����St�h�R��f�5����e�-/%Fܞ�<K�k}e�-�uN	�4*��Y췒j�0�6N)�IW�Ϫ��+J�(Y5���}���-��,gт�����ˣ�=���ZV�����l�&)��b؈�l:8Tm8��ӎ��
�2-�VP��.���i3 қm
ƶ�k[�}���.��<}��Z��X��Di0]�DX��v6\���IrOD���#;�Lh��hw�C
j��:��Yn���(�s
=�I��@�팫|p�8>�W	�U����M1�~u�}蚚�x��ZSB{���˭/�L5�sa�D�7M����B�1j�}R[�ٰ�U�/J@�KE#l���շ=a�}�]u�Mv��Qd�͙	mj!��6滊V��J?֠QKL�nf	�,��X�� ��g��P����'ҏ�nC -�9���,R��b'P�%	^凖F1�&,I���j:zh�������{�diD�:`+�wk�f��F�GE0��q���37�Hn�z� �h��ьF���#��FU�t+��yf�>L�hX߁̿�6o�,<x(�Lw�-GG���F6	��a��~��z,eT�"#�
%I��$VJz�J�,�0���˪-�ڿt��D��j�Q����9yY����Q�Db�-�R��~1-��!Yd����@��,��a��	R��f�nF��m��?��;e����PґT&s=r{��U�+oB���X��.;"ٖL��Q��Y����j�+�G�6n�)o���Ԇ6d�����s�)n���uC)Y1��W�9��y�����S)ǟÄ���;1�?t�a��- �4Y�y
�'1=�
Ϗ�3aߑC|����K~�	X[��u�?-0��U�"�����|�
Ҩ���[3�y�].��
�gh��k[
_;�V�><��	�׋��袠[�m�J=���پF�_Q9T�V�j+ �i�k�䀠b�rE6���+B���� ^|U�%&�?� �������6Q^*[�Fd��������T�̆f�����m{��s-ʚ%ߐ�i��� <e����z�j�H��חI�����E��ځEK�y�!�6j�'��CN:î��t���߳�,H�l�9yVA��L�STVU����s�	TThw�S�q*�
�'g���j���k��H����_ig�~�M�̼�(m������x�A�z5��?��v"����xW�r�}�H�Z��������?��}6sBZZq�>cw�߲f�-��Km,���1slj$*�bBi�����>{�nF��0�;"�J��4� U�}�����}oހ_�z9��)�֭Wo47�>� � �q�I���K%�t%l|o��*�i��i@8�C=�cذ�X�����G�]p���ǞT� �s���2<f�vJ*��075x�I���f��r��v��C���물��~���XR�֢�jƜ�z+Z��[��l��M̵�0g�V�aU�YjЛ�eL$����$e٨���^�% ʩ{�mCG�����V�n8h7�����J�sB=i�:� H�9��+pj��4�(U��C~lmm0��}dÕ�M=:�^�#��t)�]~����yV+�-�VH��aG�k����ii�"ZN- !<���(�qCd���PAz��cq�D�l�G��H6�X��a%�`��>�|�`�\(�ݖFLm��yG�+���f�QD��#�I��u���׭��^**��9�P���ئ�e�h��季�TГk��r�J؋*ˣIw�QNj�m�At˼oPWy�H9���Օo�ـ5����ї���Π'����wQ��ѣK�[,�O�ҔjST*Cǯ�[�H�T�)VOZ*��_k�@��Dy�iQ�8]X����p�xx�k_�C�~�+#�bRk�;�x���;&�7������tK�I�ł����Z�o.� �)�c>����7������c{�o���ߺ�Qc�z���N��1�Kf7̋��Jߘ���J�1 ��T�̱�>���F��hZ�mdo�C9��w�̙�n]a�鱺��د�'�����&0XPj�q��铚�eM��Z(��'0v�Ž?i��6 9�6R��6xp@��m�E.¨�͏��M�|��������z�6�8ښ�R��Y�b1��ބ��b/>���t���1s�|�c�4�j:]��XZ��%*���d)I��0��%�KF�2d�c�i�Z�Y41"՝� q-R��X�����@�"I���:�5I�5l@g�"�o�W�9?P�]���G��7����i(�=j��-����k�X*Ă�!��ii^|?U����'T�����;&Y��q(��^���{� ,���Yj��0������*��!���:!ĝ�[���-M@����
R���*��E࣓��֎ ��_3Zu�)�#@���ZҐ��Rڪ�*A�qq�l��*9�&>;w�+���01�A�#&�C����z���RA��	i�楖�^d�����3�����'�𲁺��S8d���C�����N�}�!���ir6���[�o��
D���4�;~����[��۹v�䡶��ݬ��{�#����P�(�08�D&��!�1��t�Ki���;���_����{�7��;�k/�]F���~�
�f?~������ʛ_�~�l����n��<�&���GI	������:���=t���ۊ�ܤa[6��1 �es?�g��+���tVo{���l�=v�ތ�x�ew�ʄ|=�V	ME�����A���1�h�	l�!���Qo,Q����y���o�>��4]�>4��ȣ�ƥ�ƺC�p~\)��2sS�|���b��k���TF��Qv�5WY��X-E�0S�uD���j0�E�!�2��{
���T֥c1��?b!T�&҄����S�'bЀ�5�ZD�N����=�n�痶x�R <��&l)�d5���c�"��ơ���	�(�0!�.�bx�o�3�.@'��(iE�uT�%�cI�U�i-���J�O�]Dܝ���{;���.&�����*j���Ϥ,֬����'����{��Q��0Ho��9���_�c�Hw-S+౞�Q���v�%�H�%
���kqv-�	� ��?��ѻ�yPޭcS��u9XB��1jJw�i__D!�����|��������28�X6�}���6!��a�n6{�R� �s=Ө!�9# �R��j9�T�r�J�uơ���C�:�G���s�k���PHO��&����W�#O����d����٧�lK-�	�	`�v}�R�ҝEa�GUH^b�C��W-|�;��)�5�E�� _���_�`sGˊ��O�q��ZL5v$���*�v���Ka���koy�^~�#��3���K  �H@��������ԓel �s�Ƣ��Yg��8�I�*��o���3�S:w'H�rFҾ$@�0�+I�`f���ʣWiE5!_�r��Ժ�5�'�ˊ����tb�ǌ�=�CSG�YUT��� 7.r
.���_RL�"���Zh�r�ZU1F`�EeC�dӨ�\A�z\��y�ɒՈ��_w5u�N�|>�ҁD�XEm�~����`�b`�Z��F"���&h��>% n%�g��A�щ,�6&��Y0sD���h�?$���
����I�(�XYL+U"���Ys��@:��O��V@I [
UK�(�~B��wq����鬿�Y�]�=Hp�AH���P`�x�'/pa�z�tH��q�%UGz�Q��S}����KG}��b^`Bg��@3��ץ �_��Y�QsP��
Y��`\���l�8<�j)�J�� !kal+�_�:��և��Q,�� �3h�Y�J;g֨&v��e�41
��WF�	�@����=m{W2ۖ_a�z����.�1im��1�Z��il���1��l-b�8��h)w<~>�n�w�7'���5"2M.Q�x�6	��6����l4������{/<e��Vڱt*�9���|���T�D�~��gK��!�C�,4��W.�=&��e�m��NL�^��գ�M˞����)b;�Ͽ���C#�ؼ��,��+����-��Gٞ�s0c�`�.x��>�`;zj{�yv�	��>{����~��`�K��MD|�������������f�/g�o��1�:���o��y�����H=$�c��N>-�.��H��ڨ3�Rs�t�����>��<@'%��zO���>k��ؤ�w	����JE�����1� ���I@n��6$&��n�\g3VV=�A������D�0��R�lBp�&:$b������Z1U��l���
-�#1a�}�m�UE�t�G��U��o���E����F!21�U/���� ��J��j@���n��]cI=�?��D�O�L*J`���h-���i��Jɤ�2R�@��\��B:�JE24�B+U��	��9��/Ҟ{g�}��BkO��V�GQ����H�l�"� �nm���_*<@dV�ߣ�H��$�#��^0��!��еZ \=���,L�,���oO=�9����Z�}6g*�~G�y6E	��S`y1ڔJ�8E �
�M�ߖ��q(�T�7�og#4V�G��V	�f��p`���<��4�-Q���|�Ȉ]��(���7��e��1���&�\�}VO��~�}�'
�X�O�0O/��m�z����m�&�.��~�!�tkw�s�H��4��y���~�Ѓ���k��tF&E_ F*�B��:�4������a2�D۠�,,`(c��,$\��_���N�s���~}ÝV�]K�$*��@���V��%ݘ*� O ��Cۊq�(3��k�u	�k�*/-�F#���C3��T��	�AFr�a��ip]Cq�6�$ LE"b�;��igW�rs�]*[�{?�&
�X��| �|4�d�$�Ct�o}�vpt_{����矴�Cy��$榘J�e���Ef�d R`�gT��H�Nf�&u�\Wڲ��mv��)O�@��훜��0>]�e���+F�I���FV<ǕŚ��C�3�"y2)��L�ax}+���0ȚOQH�X������W��߷1�չ�1�8�g�nk�C60=VC�W�]_��A��T�h+��0P��-��a���׮�r{��=	�Rlڵ����ɾ�f�:�_s��B"���*�[k7�.�`	O��h�d�Y�bY��8�L�)��Uz��6�|)|`NU�}Q!D���6����k��-}w���g9H�)C~|�:1�}y�x�##U�G���{9Z
=A K� �����!Q��cѿ���.U`	�O�Y��>���[�9;�a4F�`^0��C���������f�Z�.|,�i�A��@��EP���k'j�����O�D�TUUp#� �pF��+�*@�}��Fukྲ��ށY�TPp�a��!�-p�� hz����sȎ�����iO1r�4"`�z1�;��'�L�D}z�b�5��J�ڢ��g��e"��m$h�}�2R���A�.|\GkKw4V%�DH�Q��X�:��,.�OƎ�����f�;�؉6���2߫�ZA�ɦLi_���N>�r��j%57�ƌԁ+:�[�L�tS�F^~�][�f�]~��,����O�a�)�9|/�m�j���"�:�8��ic���"r�C�:�O/�_߯�ƍd�O��T�9�٧3��lg\z��b�Q�f2�O�U��=�;���mo�߻{.�N��۽w]o/��K[��ڦ�]i����f}5W��VУ�������g�r�}9{@o��|i��l����}�TX��2-�"8�ã��/&�4+�k�Y]��U��h?�.q�Y��� 荂�\Ah)
`�e��ifR�д��e��R�w�)�/'~d�����'�B1cMB��Jf㯣�#�J2��A�U��7���bS�#�Q�Nx%�L;KG��h�ӑ`��[�m>p�F�b[щ��J=�~t�.���bHMĲ�ʼ2N��ǭTw�Qx��+��F����
[�l�ǚ޳��Ea��H3i���4ah��6���M���R�J�bTAQiE�|�y��hy!��G7�;�6m^�M���ƫؽ����ER̀�]S�FO{��ZFpj�[F�`YC�E�Rؐ�"Ҝ9�%s�M<;ČiQ����+&6�aLU�@o����6	����>O���m���%��p���B���Ia[�n�
O�H,4:`���9�
p�o�%����:j����,R]��1{�����'���C�VZm�ʲ���~#�s%3QyM�"B��:0 ��_�\�r<���r+ڥ_��G��h��̝wY񦕞�,6��A���h����ˤ��Q;@�7�{��Q�b��)��	���/¡�u��.�UM'&GkE5)�&�s��z��H����;�C��9�-Xl}F��iO���7�V#-ʹ{b��6����fϴ�;�Tw�=��3v�yg�J�@e��y�	V�:���lV�;�#��^�>~�	�)<������~	��t��;`<��n���⌯X�"��j���qEs�Z[%���vQ���n�@[��SD�ܑik�AU�9r�o��e	g̈�#�H6"��Ͻ'b�C�ƽ\�K�>�={C���Z��z@��W��t|�dڻr�B��%�X{���Ø�qjaj�����-��#J�а�n��M���7	�� |ME6��\���M6�Y	]�X�)i(g}�~�qM�`�x�[@;���i����Q� �>�n/n�=(�h���'�J3~@,�x�l��#߄H~� �[k���x隳w;��>­��-�� l����O�z��G���> 1��Jx�u���C�F��;H	���7���Cpv;b0���؃�N9t�d>��o��o��I�y"R0Ç�"A�l�SF H̶��a_�B�A!�%���
�]o���Tx��5z��#�i�*���t��C���8�
iԂT�4i3���pw�U�L8#|��[k����T��Y�~^�����w?���:��/����ȱ8�M�=�
"���{X-_���Ci��@��tS!�D�*�`�.��'�|j��7͝C���N<�K�?����}���f�����n�U*�=k,��`�v�swİ��@��)3poԦ
�M�7}k��}&����o�y�;w�����b���E�ޏ�b���SC?��]z�r�/f,�����z��ا϶�^�N;�`�b#z�O���}���Ǌ���%F�7pRkl2��J��9��yӐ|>U��O��, $]�b0��&F��6�X(/E��J�x�F,	�F�D�o�By�.�S�=|Z�8�(�fh2pԠq�Vm^Xq� ��V��,��k�H!ί)�n ��Y�e���KQ%�r^\����^w�~�Q�QJ��9D���wL�e���z3^����X �@`L��(�H�$"�`Z�\�{��hz5��)�u�*jk�1j��U�05����h<�Z�0�aN�Y��wVGi~���K9����7r�[�I=p��ͤ���M�M��i�իR��>%�
��Dz��ƨ�\;��;."�.�'����3fZI��w�	��[m��"���+�jMZ�T����A��R��Bt�Y�+�꿶J�9`+<S:t�]\�3sD�Z�>Y���)e "��h�Rbא���S�3�B���Pj�T|�o�^�0��m���ב>�f�dH��V���
%�e�~��³O��M*IN	|�~{M����FK����'�e����jW_{�Eѷ��WZ�ѻq��\*��3�T˩�Wi����5k�zx*սӔ`{��7�S���n����k�]ZH�v >��0UF���"'��m�_�v�w��m`�+�,�4Ե�x" Z&`�g�S�� �λ�	S��3���f�B�=i64�"D��'e;ה���zN��dt�Z+����?	@�-�50��֧gw��|dGSI��q>�0�
@�ާ�\6��'@��fB�hf7R�3���6F}:P�49�+��K��6���_��HWI��QZu#�Q�%��%��L���% ��j�~����{L<PbX�;d�d}��1�IG�x�9��&`�.]�jl�a������i��9S�O�I��S�� F�C�����D��[�'[��YU��B������������j�?���h�|H�}�}�G&/X���L � Hd]@�4�������l��z�1B�SB�����?������z�g;�
�붠Wƈe�������0������j m~h��~���8��T鵎^B�)���)=� J����g�T��ӡ*]��=Sr*�mH���S�)��r�&�E�8�T�K���C�5���-� Ga����:��<s��|�ߗ���� �x����u�#�,����_p]t�`/��ӞݎD' �`�QU�a���5�3�F_<�?��Cw\�U�D��	�1y;L�{���6X�ډTҳ�#�ޔ\G���Z����a��l��Q޾���+/��N:�D{ᵿ��3��G�-�7V����'�F��`g��$��G��%. Փ��F��W�6�#��M5|�]��6�ʠo���ve��/�7��&�6�cC t`����b+@�1�j�h�q��ľ��=�MEe���ι�~���v�%�ك��֮~鷶��S�VY��G��"�4��G�|�ar�4�-��#�U����6�MZUsj��Nd�c��ZN�W�	�;��4&�&��N-��A�Q�Wy�Y��v�4�&�ƦO5�r�.�e���̷��&�jiD�l*�l���O��#��a�0o��wP����� ������-�fF��fKn0��z�@B��{H#j轚f�1�ƽ˖�{�Q�~��#��S��x�����\���h��>g���^{-�+[<~A1���T�_2�|~��o9��ӊ	Boo�3�!�)�j�� ���-{����\�6�_��ɽ��v�J4	],� }$�CT�]#h�ժ�����kc�T��̒��2J�HM8:H����GV���G*�2�B8�j�$�D#�A�k�$Y9����	/&�fU�wXn�";�݊]�V��Jj�x�:ѕ"���ēH��A�$���#Ӂ11:�{'���p��*B�SUa;6�@����0�=��_���T�X�Z�0h�8�ܫ㎹�b��Z�Һ f��X,:�+�0�;�N<~�ɀ=����d�//�����.<o���8�Fl��}�l��U�����2tضX���)�~�R;\��_}�+�$�)�v�p:�T%�VD[���5V��;�Cm�!�X�
3i7�X=Sz|�u���펟�����_ZY�^���B?�t.�Q]���.)�6Z?�w�9��������w�D��3�
�="{$})��=���˻m�QK�oŕ�#�w΅�w�KNb��]��U��#�%,ٹ�|�׀�q�$Gg�s&��m���lѴڀX���A+E�Wb>L�䉂�i����	G���9�
%/�K�g}����i�!���%� ����������/��MZ��4�켄h�>;JQ �2��ZY?��Fl�$:l��5V�u� M� ����qNQ��F-bb��b9� �r4�.�,�?�������#��z��k���L��[��#=��� ��B/��kO���y�R{��w��6$�.���8�I��ߍ���:z�Q�(Z	�I��8��p�:�1v�Ԙ�'GIi��%v��^"2&3v���_}h*Ы��/�w�{q�����k���qG��c,���I����E����;�~\�O�v������<$�k���^WE����n �R���u�!��U�d�ӯ��^k���-7���A�����}/1f�u>���	�z�I�O�d+�l�������i���3{���S��Z�L��8y���$���n'��h+��ß��$L�ۭM��P���	�v
b�$��@����(�>ظ����E�!�o �m�����a��?�k���ꋙ�l�{�r�e��Us�_�=���~��K��㐝��t�V���@����r;A�gΤ��AA�!Ep�iG��ۮ�j��wY*���xf[���c�k�cm_:]�k�z|�+"y���l������&B�G`�r�=�y y�	Sg� �'�أ�y�V{I��N��+o��B���G~������c���N�a��(��pGI,�#=�wh��T��Љ�,��K����]�M�2
��`��얙~L�]�>�1q�j�^����GP����q�h7F�>4v6�p��v���Ěd��k���[���F$" �0�8g�8[�=T�	W_u�8�`*ɣZ:4}��1ϵ�0�� qr-)ɻ����8�յVAh�"��-�ȸ���0�AZ��G{��^;9�� b�X�O 1��'*�0��P���\�>�$�c5)X��^[���h@���ɉFH��h��7��.�s
�ѽ�f�H���=��{���Wo9�ٳ>l�uݴ!����B;-���E��S�����FKe]�^;�Ƴ�
q�_���&�����`~������#��tq�� �����g��On<�f�'�e�GӠgs2B����fa_��R+�Ck+5h��61����Mv�%w�>��K��%?�X��6�������gބ����i��p�mC���g^���mq%�(&
P����v���@�#v��Z!�{Ӛ���{��ƥ];��� .<���x�Aw��_?d߿�b���'?��z8b�؟]�]��33y7��5�{�)A������v�$g���Z7
�|y��]v�M7ۉK���n��m^�Ͳ�>$a�f�An���S���}<ɔ���A[����bE$'��L�?N>q��?�e-��M�$i��~��>�@�r�S\^(g"ɦ�D�d��sϹ��+��ҩ��2*D�k�� �G u�;;;i���%\,�k:�"AO�>�%p��t��요��5Ilu����;)%Bj39$/n�D�nf [Ô,�!�۹3z(]�YCi�E耴���[u55N��Py�C��i��Hd}{,�U���u�G�I��6n\*f�(����pA�E�?�J���n��Sx�V{�g��Y��A�Eb��-���!��A��
h��@����V<$�X+�;��)2�I�>�\��ڂ��H�����~0��)	\�y
��|x�F�F�|����V�|e���.����O�TE>�{,Y�g5����ߴ�=FqQ�rƝ"�����{�����C�e�+�oG�g��%R�~BI�F�(�B�ƒ�1E�����>��0��'L=�ញ>����DL�aދ�es��~#�;&U����^W��ڕ�'iۍ�]�VL��Ԧu"��q��k#q�-o���T��Wy㟹�k憐hExH�I#QȐ�G{{�����a��v�y�ك��ɍ3��h;�����^~m�]��,i�q �h��w����]�я-�Z����F���o~�-�R�k$(���r-|��\`g@��12�.R�y����MD���;+��)������H~;Š !~,
��[���,.�|�����*�㊥�����~���ڊ��m2m�g_z՞x����~��_y�U�[�{��Ha���ަ̙o/���62p0s���p ^�E}?��)���!I��G�V����6��/	
jq�E ��[��fU�<����Ն�B�������}�.g"�͡��4��R��.��
5��X�kG{�٤���׶؇�߷	s�٬�s���A&A��㽯�@ݍnQ.*�'��j�����$�(�� �e���s+��M�G�A�Gm�=�%����J�	�j���y��EC��@��9p�tp
�#9d��I��n��� ��B;�X�nS��>�|�$r�H�����������!��H�CҐ���L�~�����v ��:��3�+_8Ͳ�ɏ~�(���h�7J[%i��e��D��i.,���ƌi!\|=����f�ޞ
o/�`�@!�+��³��j���J)&�9 ���{x~ζ���u��5zꙧ�CO<�LG�M�������M��/� ��?��h\a��n��|�m߳�������?��W��Kl��2'�{�5�Y�ܼk�bگ��y��(g�4m<Ӵ��y��rW��ţp���`X ���A��z4�����m��_�.&6�	�'���i߹���?�����ط���W%�A�j�@�v�X������Q�����4}.	�Z�@`bOS�W_{��s�yv��h�}��
ӊ��bj>n�H��2� )8�P���(
,�h�=	D7�Bph{"�N3�f���=: ��Q��e׎V�(I�$g�A��Ga*k��e��	��ު���#��И�P��kbWG��nBK#��]���@��k{��q�p,tS��+�����t���$Z� �G��qc�t��8<Lk��J`��}��6�8�W{ấcR�پ˰M�}�N̸˙�N�_��uA
��g�:�g\@����{:��KT�uhy�%P��N��bIqa����D
�a�[ډ	��Uq�N_������a�JB��,dP�>�^2��O��r�~�%N�z������Fn��\?����k�i{�iP��K8lME�[g^��L��t/+�i�k�;�\��_}�!Xch����E#ɗ�@�rק�|���b}����֘��+��%�!
�x�>��LKg������=D�T��B�ĵ���[�cI������	hp<���ӝ/���z��0^��H�h��<�'���	��ϻ=&-���*�>��Ϲ$�3����9Pɾ��`� K�?>s�ˋu��q�x�N�a ��t��Q�n�B�y�|�=������|�^~�)[��Z�*�C{p�]}�V��P'��;�dS�ZJ�5��_��%W\�F�q�����U,�@وm�9����&8;!T�gٱG·�@��J[$n��:a��~�q�J��ͯY+�〉��N_���(�^�|��}u#�"��9�A� �;�����߰/_~�}��?q�	�x1fỶp�����5WO��n���#
K��ig�e��c���[H���1�$��r
���yXd���!�AF����]u�����"�*9tU��k>�*�Ie��S��S��*|%m��a @H���&a� �l8B\chPU�L�d�yY����oٮwW�:F���5���kk�� ��R�A���/�d���ٞ{�yZT�1� ?]��Z�S�3j�HC*�j�0�hC<G!�J���T��1⁸Ju"'I�$����N׀]�k������I�{���,�Q�d�c<�W�e��G+r|#�!aH���J�'da�-�N&3묦Sd���W\��Q���HzcI4��#hj��7��߅�^d�)�IU��Oɐ�@��L���	IG�v'?��ِ�g��a,2q�P��}3��4��	N"�s���p&�"C�?dlޕ��m�{�[A��^a�,�r�_���vl~�m��
{��͐�[���ZF���omݞf�AKq֜���O�s/��C�����D�&a`O��������¥6��Xi�8�ڹ��0p�I^j���9�Ղ���xF�<KL�����;�&�����C�5��Ʈz��?���_w6�����C!۵u��/��X,�	�:^���	%�_|���Uaº���(��<6C��V�ޮ��&[vх���<`�п���ډMm9����v�����u����w����;�����{��L�)������K �������X^=��R�N���NL�Y�a�2�}�u!m� �M�Z�=���Yđ�$�r P��
��I�OOqm�=�s@L�/&���"��dq?-L�ǢS&N��e���|>}�U%�pp�$&5��b�z���x�u�P��^Wa�1!;|���n��l�g;���B/pܸ"Ct�������iӝՓ������'�|R���^D(yb�bP�aQ$Fp��J"��K/��A��gt�p=10�X�d�P�&'a�ƺ��E��� �����LGZ�E0Ռ㇤7�)�b4�A��'����δ�%b�T��'��%B(������P�!ڀ'	�9�8������ �ȫ�o� *��1~���c����?-�O%bM/�CN`4��yv��-��'����'%����8��Ե�_�0G�w	��ߒrpʏ���A$Au��B����{?n��FHh��<�ui��1�Kh4}8&ઉN��<$l��~�C�>ሹ��%���	l���P�O{�~�5�;�Ƥ��{��������z��կC��{ŁAˬ�ׁ���?>sƦq�b*z��\����5��}x��d�*c_8=�����v�Y��m���G��)@�s8|��7���������P�1)7
a� ����Q)J�T
�"����a����F�K�a�R�lb�w�G4��~xNŨ���P�G99�@���w��>!�96���0�H:� /���;�������s�dL;�O���:g�Ǟ��
;d͇g����l��d�)3����bHT��wLv1�L�u�:�di"�*Q��^���'�
��<���M� (0�ᬄ�A�|�'���"V���T���`k�d֕��������ZFY 9����`m�M�4��;�4'���;��D-��&�iEQ��"۵m�=&S��8\��ٷ7X� ��i�53-9@U��0�!�� iK����-#�$n�NG(��t<(}�OmW!�e�[K�O��$Qt_Tq�rH����W2�)wkoĿY	)&OΏ���F���=` �f���Q*����4�K��e�4Hg���,��� �U�X�1�sՠ>����w~�h/�g����Qa{��@R��)�[���-�J�Ip|L�ŒǂbĒ���+g�45獞{�F�����k#]��$���N~��3.��u;d�qB�A�?r�/@�(b2�r�(�o����IL��۳oU���,/���@�C[g�P����=���ۿh鈤L����]{��ݶbS9�� #���8���.F�ke 
�����5��|Nb��'�E���JD���$1�{E�!��_���y�}�b��=t�8�S�Y:c$Ҋ��ۑcy��P{M���֖�Y�R	�j�K����PI��|�v��/�[���=��w�I�,S 	�eO�"�P���tE|x����*Bȵ%�j�L|��HD3m��f��o��e_Ą��.�4p�9I�V�Ƒt��?!J1���D�C���`f4I�DD[�Gd�{iw*�ҿu��Q+_ȏv���6P���s]��%(>���7o>{���I�OE����2U���i�k��?c�<\�\��m����-��j(߃v\���)��i��~꜉n fH�+&�D��� jB�W�rN�p����F|6����r0"�eߓ��X�������=�>a�}�:�R�����l��΢(F��`#Ϗ���a&ڙ��P@�C�@��w�R�r����Aі�Ď\4>������!^k�K����u�Q��=�D����D�������Zwh�rM��wȿ�O����x�*���UzM��k[
1ҩ�"�����C`"���z�Ccّ����Jp\۝�qCYN��+V=!Q�g��GӔzO�v��hD��F����k��.���v��������f���K��%��O�)B��<Y�/�/�3p	2/�=��\��������ӈ��"Ib�o�}���ı4���1M�1��{�k^rG��9��zL�Z�ZJ1��&�P�\�*Ҡ�����`�0 @�M�d�?}|�$�E�[JJ];2���3&��#́:�X�hC�#�̬���ѳ�v�� �0��g�ȝ6˚�>5��I�zA�R���$�F��J^h[a~!j�T�l�*�Fi��WY`-���ny bc��VN"�^c�4笕Qx�m�I��oGk��[sfZ�F{i$�qE�f33f#��l���}r�]~�;���?v��_o�m8d�����p�����aO>��5P1��\M�����[�q?�@������S.�&���a����z*��P$�1�ѳ���j�6����giM919�P����6��S�#����f]R��O�S=[�h��/���9�����x�U0�Z�EO a���_��s�ˇ_t��i{��_|�i�͓����$G�T�q�D��\?-��4��D4��d�6H@�n�=�@qttAb��u�%TD��_�}�U�Z%Տhgѻi�x� ~^7�v���D)�1x6u*���$*h6ؒ��킳�D��5��g^�%2jW���H����/����]z�+<)�Bm�v�_�΁ӊ8,$�)3l��u$���fqm�҃�D���%����GK=��8]������Y��1֨(	�D����H�.s�0�c�q|B�\������pm-��X�ms���'ؗ�\b�HȜ�A>�9��'���p���s���m&��f����]�LH�=���[o!��]m7^y�U�=��$���=x��VK��֐���k��;䁺в����ny�+�7GAIf�B#BP�H�cX�}�RSxN}`�F2�^��r�����=�m�^l��ٯ���1��˲��A�釛��^�X�71��B&CIǧ+�O�jO�QDa�i�5�7 �]yݍv�y�����-[�y�M���|�[�Q�] AR��g��S�L�~o
ϥ
�4�7Y(Րl�<��f(}I���!�8�Ԃ�X���C6�#�nw�
�$!�$�Ȅ3��/��@��{Bn�h�rF��+Z�~#ע���%e��{�ٲ3�v���*pp�u�p�z�s��ԉ�W�5��![	��"~7�ƠPY��%��:H"Lr���E�x���k܁T<1��8�)�]��$z�S"5�x@�*q��HJ:��$��"K14�J�0C<��|�͈�1<���y���m\�?��˝z��h�����}Ca���kw+<3��4�<]�L�As����0f�fD�`���ŽC�MmX�O�Q��{�C��#�v�$"x�9D��� �ٱ6�[��+~�u<�ub�5qǹ��ļ�`,��֫��p�=xq|���z��O}*����R���o�z7K�3 Y��y|.q#���F��Ջ$T����{���X>�����]E'wg�LE^�݋ȽU��h�ڑ����{�%��H{Szg.�+�:��$g�{� 9���^D�C����5�E��{��6��R�폹����
��ٚ�x�:7B׵~��A��gv�j��@�w�!_w��X��$L�n"~ãXv���ԾE�V@֣������=�QY55��`��I�9$^"k��448伢 'ʓ�ܭ1��7��KSu|��U���L^f��ϩj[C��J?��x��8�l뉲�kw�xLň4N�4��C=���CY�2�gtƤ�M�Dˆ�#*ߑWVZ~��6k�\��7���K]����ۆ���~_��;�-����x{���l��Iэotۼ����c��lB-.��Q�Tc��.Q�B�J�O-&o�hɫ�rS+������r�B�1>uAF��ƑX<�#`Ӫ��h�1I&g"�;�.��=�0��k_�2q�|6;��i�$ZjƸ�w���?�ZN�[n��ŬQ^���Q^�.�@��@���*v�U��.�k�)�H|qP/���� �8�P�NU�* %m��C�|��� ��q�%*3_M{���6�Vk��N%�!Y���j�7��6o��x�+;mU�&�˄ g�UYu�_����;�_��i��$���u2��M@�fa�A����.~Bhd1�螇9	�0}�g�/S��� /�$`4�y���ܚ��k����˴�@4��a�#�۵��h�Q��~!?�7�+���C[�A�aJ�+�^d��e�I��O�ן|�dXk$!R5�fʒ@�ղ�rk��_�xpzv�3��������l:
����zu�U�k��8��|���j3�ZFc�	�vE�pS����:�sP�I�R�B���,����&� �]�=c�X��@����=k_��R��w�O~�{7�3��hَ�����K���%�$�ݣ5&Ę;Ł/_I;H�l��h y�2hۅ�_h�~����S�ՏX��n�53\�ܮ	R$2z@�z����E����;��^$Bb���H���(,��H�FI���]&���B� 	ē�T��qȦ$���i�J��d�X�R����k��8�1{&�Mj;�sJ>jEX���lUW#z������+;K�;�	������(U�!.��e�Y�q;��h��gEŀ㗯m��D�8�u�Mע�t2�5���_����@.b#�*~����� ��U򤉸L����j���o��׉�Ƌg΀JN�8+.�n�5�_���J���@�G��������TY� .d�?�	x�V�0V\��^�`��!��$��W�+�׆|Qbq�F	X<<	�x��U��N��,�������3�Զ�06��C��.�.5��"�����(ʴ��8b�+��;Ƥ-<*�>�:"����>/`A�Z�Y�[���y�VcV;���ؔ���t^(IK������C���3�tCP����^���,E� ����Eg�KA��|\�D�3c{е�\,�RIX���cPɘ�T��s�����O�R�Z��r���^�..-���b�R�O�я�$>F���k$��$�t�e�����ya��u�<���yGp$���5�}�s�Hׂ�UZ:�a�����<��S[��#�	�M�&R����0��`[/�u�'	�=�1�!q{b	�Ⴊ��h� T���O����g	�a�O�*eż�2�0��nT��s�y���Z<��D��^��1�l8Yjd#6X��߼9��혀�4[���VC�eh�Y�R�z4D[���$�4� ��AZ�AMc�������d�]p�}��߳������Y�l��I��Ԍ"'�Y�����:t�bPc2N���B�-�X�!	nb|�2��:x#�1Z n_��s|����{���U_Z�ë�Mn�y�������pan#T�B)h+�h�����*�Ǖ�n1�Iu:{�lۄȬ�1<� �O��o�<h��Z�E��������m)��H��$�A|�{��{�^�3���/OyX_p�|$	p��Z�o�xL5bU�x#�3�Z�2Ya�4�T#'�:Z���E�L�1�	4�E|��5��]�I2RA�|6��Cd&�	�H2�6kn;l.-�x$F�z 
�9�B+�]%P ���G�3x�$e���F����l�f<;]��B8�A��gY�>�F����֠�M���Ah��1���=q�5k�{)vh�f�`��6a�\��U�|4����^wٱ��hלs��uGَ�v��-��+y�uҹe��D+���]_��z��{��<̻���K�!&՞G;/�p���2(�t)5��D�>l��}ʹ♜�O"�ы[5� ���C�w;�ݲ3���_m��,p
[iW��ޗ�����v��~bM|�D�%*�n�>�sS���P��"c���S�D蓌��u����_���y�2��+?��}�
���	��5��<� b���(�V�k�O���a��(�%�I&��<�h�A���_I���H�;I��y��\k��ϙ�
ې�PA/�G.��b�j���="��O'�H!~R���O�|$�eN�I������)�lO=����������3$2�Y�n�8`B�����U-�X%�!&���5��%�w�5k� '�������;-?�="��M",�a��۷|B��v(�i����	S� nYo/����>���xx�>۷{7zih��(��*(�f�0�K�B�b��
ϓ����La�!'ݱ�ᮂ̀�i���}=�_�I����ؓU[_
Ir��s�YP�>��D&m�@*.�V$�S���5x���>4��gú�w�E���6�X�]��#��>�7�,�$������^��㡍�,c�=0��2޽��h��A\H<mQO�J/�4�\����t�S\�%N���{r�ڸ��e`*�q�t��Mz�OZ}��3���I�ѵq�Iw^�]�n��Y��%��{�s5�+J��f��۝��>����=r�w�� 1!���iEP�O"�����Kp��X֩$9��~��Ʈy��>~���^��~0���}�>轹{�u	AV2�=���_���k���c���'a�����Xp����g�#T�Nm�J+|pUއ]�t������45�7��Ta�<���;P��X$qS���3$Z0ILYj�[I
R��~�^�*�T4���dt�Ƚn�Nۀ�������K���u:��"t U
~����~Dm9�A��S���q���m������v�����aR7b�0ɕ$B��!�ݺ��h�$Y^v<H�=-Ֆ
����㏞�пts���EҒr����q/\�T���)��s�Xd9�l�X�x���uB�$�q�܉�-�1_B�0���} �M��19==9���^~~�-g�p|f2����|�z���P�@�����K��~��2.ۚ�w[d�<{�g�����6~� �l�D<�Us�|��`�1�ˣP���l쿄u)�f�5x J�Fܚs[�mՔ�jIK���p�����K��s�s�?y��J'ػo�B���z�-v�qg�Yn#A���OO'aCNd�)�u;S���YO�Ęp��"��F�D��m�n��v�~�5��`�(���}ᰁ ?�3s��	 e1�D� �k����� ��G��2���~W,
�(P�����٩6Y�ʃUv��WXlz�����Y3��,�b7_}.����_��*چ�+߻�vq»��|	m�z~�� E��๳�Hd�>��[V�goa��;�;��m0H0y�2fg��ɧ��c�5���}��>�b&��S�+���A�Qc�����{wY4��o}�h���#AC�_�q�9i����O��o��~~�������*g�8���5IP� ㈍б�*9��$,T��Y<�����ϝjW\�[��� ������}*�6�4��k:SB�~�����'A��h��h<�T}��+'�$8V���h�}q��cU,PL��6r_�t#�;QS[��X�RX�\�h��h�\�P}���+.M�
�ޢ�@���N�J�W�G�]��v��2�-�C�DT��1^�J�XEg�C1HY�XG��}�3p��	��@Bŋ�$�/��u��:�yɟ�/�Hp�{f�
	]���Y��#��d��>������U�2�A�˚�-��NR� 2	��Ia�;;���^�D;n�8��uV��t(מ'�'�vΔ��ֺ�>�$6����0�V`�����P�Wd�*�8Uk$�p	�s���,�K���-�Z)(�^�R�WR0���=;��1��q��3��4�B��Ǻ�&�ֲ�aJ�4L�XH�E^������1+�H�t�j>�a�5�Uu�47��#އ7I?�X}��x_w���{������D�����8��[�))�{�to�F�Oں�W������^��I���ñA�D������Xp�ם���Zlc���{,��׿��u�9/1sR�7�-tNH�W8םh�0'U�U�Y�U��2k��I��H[��y���{��zD?�Z4A�ИF�c���oQ��v�V� �
�0E��&�h��S�j#�uL�h��1������P�Y�} (�s
f�<M�pt��S��`�=��6o?`��7y�Q�\���� 61�Axl��V�!2kJLV/zv���+���+��l0.��U2���I lpV"{QWS�0�\;��Oϔ^��g$�����uAf*�� f�����ER��?�M�������5i�D�n������P��<�~`�A.J�5��Bׂw�(N�_I�G�u�&��/�nZ���]e��r�$b���x4�4Q'���5{l��G[3e&$�0՚~O�h
S�u�Ѹ�{������x���qg��G"�1>���Xn
��%��靹�����#�~l�i`�s�!c�w=�>^S?���_����w�:��,�y�ᓳ2l��,9�a�JY-�+v-�V:n
{ܫyg�UW1���ڦ-Sqy��
21J>XOK+#�&L���@�N�)n(V�Zڠ�!�ho?(.�V<�?�w�F��\��0}_��eB��ց<���Sd�H7ߡU�I���MG�k��Rx��Vv��yEM��O��Sh�j@z�֯���0�W�As�j �7��XO���mc�5�Ӿ�
{�����)�dJ:A ��[,#�֌mR'�_C&���~�g�"�ީ�&�s�&E���T�>
U�������\�?�j����p%��ᐍM��	�vzt���O�7o:�~���o~��O�,�R%&
��iz��I��C�cpȶS�����w"N{�-=��W:�[��k��OB�ݍ͙�`�&l�t@�x}�H�C z��9��ń`IgJZ
CB��3Q,�v&$�I1�� �N��H,Nd]�q��!n��C����W*䑩x��y2�a~�g6Lb#�.��p�i�B�0s�,��i?hH��W����s�)��[?��*�ʡĝhbn�/�����L�qB<�^���gOgp��>�a���p5q/JڴeepI��=�T�kwB	h��aZH9^�\!]��w�_e���l��"d'�I�!bks�V!�b%g�����c]���_^ã�=Q�����WW�d��g�l瞵�ϳKcb�բ���p�S�0��t��֖�Y��V��4��u
�)��Y41Q��X���(%A��t�Bsm4Q=��I�q.�E2,�L)yV[X��Z���<�:���)ܫ,�#!���U8�I���8�(z�d�H\u�I�H�3މ���.Εg��hB�(F\�ġM�kʘ>Vɮ>܈ko�cU�z0 ��{�-y��&�#~^���t�!FD��n���I�xh���1�MI�ӛ�ڄԎ�"��s-T���C���鯍^�N��5	��$�]7��1�i=~|������&�s�ŝ��S�.*V�ɚR{5�/������2�{���3'aJ�x� `_������0M8�5�Hl�yp	�A���{�T�!�C�a���Њ$3)3H���{�7�s�{��N#��WH�4q*��|/R�_t\2-FAM�A����L/d[�oW5H����

#��"���� �]EDac����� ��A��0(�ZbT���ջ��QJ�Hg�����Qj*2R��z?���MH�{��{�k�=��s�������	ˎ5B��b�#[ IGD��Ȧ��B:�x[ڂ`ֆU��=
b����$�n����)�j�C��hm>q @݄�e���:��@aܻ��|�î9�$��C��-����$������<\�� |W\�9ˉDؕV�V��%���󸃖E^�eX�O�wN;�5�`x-HW�(�;�U���e|�I^"թ>9���Lݏ�M��T%�o'w����xr>>��PF�Rr%뭥� ��W��Y�:����<�C�V%U�����Țo���h���/��m���<�k�'�#�����IPGF��q�d���<�FI�1��{��߆a�#aڱ��MS���|�B��TE��isE	��V�&��w��D�+�=��z���5�G[��W�x�F�N��?����rS�Hh x��v�E����q�&m�c����:j��5g��9i��r�ME�n��c�	��|��̼ۆH��e��_r��?Ta�|T������$�
��uP�H�C�Z���R2���T��0�7�#��R�@zZ�l|V�U�j��7�	p�R� �]���EAn�x���?�G_��n������އwg�C�\�d�k�}2M�W�;@&�I�N�;o������_���jKF�lH^�$��HA*#!�6��zA{��}OGL�?+@��#�l��o��[e��ͬ�|Z|�3��-C3o����Y�Pa?'s�)p���-���t* �w�M1k��Ɖ���F�4�P�>�xE�L���ߨ,�$���H�AH^�|Z���8�P&�e肈/��8���Jd'4�I
PL�D��?��àSCi<?&%u@QRX8���Q.Yl��"?���ܱ�N�ĘAۊS��-��HwO�z.^�
'[%\Lh���n��?#_Є���f-�|Fгh����z@�h5���ʀ�7g�{w;� ��a��\���\�"c�����&[`%��V^�d����'"��� ��qw��dzM	�������Ι���-�~f�8�r��+�P��8]ιD�1�#�wMxK$T�*����c-�@FU;�'�ՙe���ƭ��v	$�B�up+!��x���#��d��(�)4W&B�W�B�&Clw�E
����8���X� ��= �*ɣ	�3�սNg��bs ���3�%|<ޗ(@"����� G,h_4��q�X_������a$Db�G��EQ�BYCu�p��x�����=U�PY]�}��}�u�}�@���Wf�8(އKu��S��Z��P�W�o� a�??�E^��嵉���H�*���2?�	S&롗�w�3�.��0��J$����g}Ց��$�S��?>s�Y0�'������8�0<�!�h�bQ+#��[̓��"K�������A��������2Z�d�"�*��E�8ԆyP�$�<�)�^�1FV(�5���bse"]�E'_�$4��:�8ce���k���94Y(�Ӧ�C%�W�U<3J�)6 MPK��Q�I�_Y$Ap�\�%ɈH�2^�UK5��;��#� ���L8#[6m��[�a�q�mL{\8d	j/����{��3@�h�p�D\0����|��1�I-�0��P�ƪ�f�0�����n'=�u�H��s�L,�pZi�L20����c:��O���IlD���4Z�~M�ɳO��Iq6%�^=��M=����"r�bW�%`;5@�2�Ct�DZ�nG$�Q���52�C�%t��ߑ�������������HYZ���Ǘ�}5�B:�!FR:���(�����FU�*�
q�D��d��5��Ã{�lJIZE=�r�*�������'��yO�g��� ��	���=����.>�tk�����ی��ئ��l��cl��Vq`7�|��\�"1�G3����NZ�=�L⒋��Eu�v���Q1��*P���Ll�ʉ�����|#�:����K��8�����!�a�	v�.G��=�O,q���%)��'^@�s�]v��p�F�K����j7�r?s�}�K߱���v��'ۜR�;vS»����l��lnϼ��V�1��s�5`��`[w�d�K1�����7�V;--'����1��~,�d�Qs�!��i��Y`x4�f�[���A)�Hg��2u��JZ�r�0S�w����;��[��~�]L��0�l��N����b�?8\�.h���n�t��vڙgۍ���^^��%����;~��5��u5���q�?E�+*@�2H���(F�(�{�L�Km��Y��6ڧ��qK�aj��~���s�3CǊ".ͪNZ�B����T��)��k�� ��8� �)���3Q="�T�ҷsmu�f�:`�(ٕ]O<�F��	�GM*��-Q��e��H�j�ܟ�x�G�zAb��]��3I�5b�#n��4%����Aý��g_�d�s�֮�y������h����>~&$�5t�>K��!��^Z��L� <�^�{��k+�q���Y,5���s"1��B4��L4�y��`u�K��ڊ��9��A�4�=HL��1����
�X6�c���%r)Ι��n!����AR<���,LM��vc%@�|Q;�}ˮ�Q��@)�K�ůe])n��
��>�s�
�>UKJR^����,}��w��s$�&�8+���H�,Ԏd�v��@���Jq���� A\H>{:@ I�!Oz�G��l0���~ك�[@G������``C��=�<��3��j_�h�$m��.�҇;[59ʿ����a�Ĥ?��*��J{N�ɢ�iѹĒ�S���\����Y���tP�8�]qC�@�q���N:O��%�+�)T�gM���05��78ґ(ep��\�GD?GP �y�V�&���1�D?q��́Z|���Q�*���3�dx�����M�J�R�F�� ����k��S"�1@ɷ1�62���g��5��K�V��Ϝ��[��}_BO�N��]��6��5J�#�'n���(�"�ҕbzMZB~8+Lr��A�F�A�.������t���n<{��)�3'{zL�7�rl�g���~���Ν��P;�24,k-s�\K�BƏ=�n�CyB*�^Q#�Q�u��[�o4�7��+�C} t)�t$!��Њ(X�9�Đ�'��{0B������n3u���[��}�1�u�+B����d���M[�S���4�~���u i�#@��Ght#��^@�ШK i[�(o��X� �����ol��9v�Ys���m_���D��֫�ڴ���>��oێx����S�(j�.�1F���Wl��dL�PA�<qE�l2�Tϒ ���}�uۖ�xm��<F�L%��~�h��=�AH$��9|����U���%I�`c�+��ΠM�JC��M6�! *�`��p�ؠ���D�B��D𑭒 %MzFQ���1�
A�T�����|��x�l;���f_�����UI´���k�w��O��0��1kAÇh�~�cR��XiI�sϷ�q��^�/�����P����&��r퉶x'�^|���$��^������/Z��E����}�=�ά3| �~d0��(n�R����@�8�z�}�C��n�#�g�1͞y�O�{�G��{�h�]zα"�f�@��Qh�|n�#�h��mv
6_'=�V7ڴ�4۰y����q��m�����O�L�ZM�
��#��C��Sb��'Y>�0͇j���x9�E��~���	LJ83D���\|:U���N�`�h�+o�С++ĺ˚~�e0u:�ׁ��>��2� G�ӵq3�TH��{�|����e��_�ľ��o�>Zar�裍�Pv�y$c��>"o7���]n�]p��|�]��+��3Ϸ��
�:��Ic��y�YG���)�&��6�|:�T|���xڈ7�x��w�bk`b����:��,��g���%W��x�FG�"�b?���@��1Ŵ���~G�?��#�`"���B�D��{瓊4��t���{������ne�%OD2�A9i����g���vn<��l��)`G(`c%�}C�����AɃ�)M�G��AӇ�P�6���&p��W�}��8ژ�DW1��h��~k�!	��Ni��7��}�H�Y��N���B~cRa���׶u�ZH6����&&���0O7���k��es~�<#��j�k�u~a6���Abh� 4��B�*d����cӽi�6m�<�`T`��t�Ė�H�b@�(�z�J�Iq��F��F�I��l�:�F� f����X�;�|�Gk��2%��-4G�݁
���"�Z��NI�ǽ���_h?S�>��"ǳQ�B|I��A5c��<�r;�����)�{�f^����XI<P�k�Q�Q��{�{2��{hz��N+��nqH�LB���^����I���)�A(1�X����"4$��TmV���y�M�Y���z��ư��[����4�*�qqU��{�Hʣ��h�F��KRT���e2�1��8��'�x}��Ւ��Qce��,��a�@K\|��o����3��#8��J���5MP<��`�z�##��g�ZH��>�>����%p�SH��<���kt4b���C��[䅩y�Yƾ8����Ō=���AE;N�7"ܷ>��H��w��MGG��ߘ����B��W�0��!�O�:��h=j�N��`R���� (\�l-0��N��Ejr����d&�ܸ��a�	A?���i�MCu;����zG�_"�OX��3�����O����E	~%SO3��gKN<�*���6ةG���h,o���l
�O�C��Z���0/���eP� �����SeI�MJesx��XE�~�xl 9��'��i����_g�{v0���hIJ��.�f2l����~EE�B�gQ�d%2�Z'LK"�����5��t�'c�����9(3��}�~�;;ߦb��8��&�eZ�$�s8o�,p|�3'50�A,�gՋh�/.d��6oXKBoɍ3x��'��z3ցI�(j����(���L��6Bn��7�_U�(h�c�R}�1���Ri1
��k��� Z2UU��D8P���qr ���x{2��a��"���B�#!�Z�f�p�(wA09�):В4��u��":��!��ۯ�/���B�q��GX���w ����V��	�/q#�?\��y���]sՙ��t{�^NE����4ڃ9;�*k /v��%��?�+�_�F��ݿ�N$�l��EE;�~�g�q2^Av-�%�u.��3��8R�D8P�$���4A��t���k*��>ξ�N���-�6k�	���כJ��S�����6�G �cp�,�i&O���<��0�S�UPK���4��z�� ���Aޯ��D�v���J�"�>��%�	�K�`�=���E!D����҆����{[=-F�sI<��ƤH��f��x�0	{J�D�S��~pϓ����dw11��_��� �'���p5!�^���z�����%����o����$���|R$�H|�u�m���o���\ƴu��۴�~��{:yՕW��0_q��s��ш���?�C�江�X��MH�C�G����i���#����'�5��5q�,��՗�$�r}c��	I!1jB�5��6m�4ĭ5�ʴ4�e{w���'��⌋��6
/J��>�DدC$&"A�A�\[�g�V��w�癅a>�w����J�A?�a�*P�$�{>b�1<��i�*Ti�>�|��AT�R�x-�����	h��A��c��j�n�P �ӵhF�M�A����i��%zk#��ɵ��Hv���à�i5tS��l��$�$b���<�4��q�(-��o����s w��츥Ki-�َ][i�k.ϴ%f��Hx�!�p��
{(�>5��s�I� Z��D{�����r��h�Iz�M$ej)
R�P�2OX�3�u�ʏ�T��h8��Z|������e���e<��5���s�m�g����jח��X聢�Ǵ-Eo'�wS�����L�"�
U]e���S�yl^c��{��
l�k��s�t^�q	 4�
$��ɻP:=�n�-B�8$z�D�AE���K��Y�h����~�xHpG�ѵR0��	�!�Y@�:.8��I��݆��	�IR����[tJ�;m�i����VѢ}��{_T�h��HB{<�)1ѽ�Q�N�%JG�`)��P��\��ɇ�.!^`�(��i �	��ÿ����o��4�]1���K�G��N�����)N)�Iz�C-��w'n�a��?>3&]S'�4G�s��z箧���I�	8���VUV-�JF�բ���"Ҩ���%W��5Du=�t�_�I��T�M���E ]q$�3wB���qQ0�Ѓ�Աk��\Dɍ>��g�#�� n-	�ZK����ԃR�(�E�^A:�
Z�1T�cM�s��@<,1�J�/�
�	j��9�{���@Iܣ.Zw!*�r�+öu~)e�B:5�,����0�M�NPS�r��@�lIJPka�>�(�4�C�Gű���s�v۷� ��lϮ�v��)6eR���&!���&�I����`�G����������	�	T2'q�}���a;���D2�>���� F�,@u���d�1�yӅG����*�#��kMC9���^�j�"��8��x��|@�\���H�d�&�|�%Җ���0ϖ���sN�m�|a۪2������Φr'8юyq�:���; �Hr�����i@��Z2�S���Nf>��V�d4�9D�\iմ��u�������2� �k�c����>o9�� ����=�=Z`7�r�3I�A���v���䆊>��TQg���X͟�?�w2R�f��
ˤD&
H�/߶E�zk;�<���K7��G"��P��d5���icO�)�Mn��O� ����2b'�x��xq��ڰ�B2ٶ�}?{$Q-����1�8���m��I������f󧣞_���N.tzkk������ȴ�W�zdٞmH+4������nъU�S�`F'���oP�0BS��W ��A�k��`J���W 7�ME1?m�U7�ؽ|�uٷèƫ�,e5�ܰ�8Rⵀ�6�$|A�o}�j��Ͼo���O��j?��Y V�`L>L���ƫH®��|����3�ٜ����믶��W��=C;��y�2�Ӿt���[o`°2w��u����cuh\��2��sl?��|�Q���م�Kr#9i�!�Aң�G����1G/���wY�}����z:i	MR	E��L%�e�T$Q^��,ʟz3��g9l<:_�đR�'�T=���J�6�&b�K�@�@p4�M"�'މ�*ޫ�uث5/�B\��$"�;uq��C�p��yh�1=��OX(I� m�(��$�$a�XB�k���: �'P�T�C�Ձzdء�~��/���GD:��X�SG���g$^�~�%k'�v���,������Z|�QbP
�EI_og�[���;=���x�q$�����h-����m��("��E�����Y"�A����k�eSl��������c�$X��(�i�)q��\���W�hp&WndR���Z�u���ފ%�,��|1�V��2n�]6lJ���CN:H��8!�X�N���I�CR�W�SS�!�9�H���iϽ��f�q#Ӱ�a���_!H�7A��~K�:��nD������w�惶���$�[V�P4� �5�n�0�Z'��3�'1$��f����L'd�A=%`��U�Tn�R��x�-��#�[��f�+SՐ�pd��Y�q���/
%%���;%��Y�_NhY���:&<K��ؖ`|ʁ`b�������pB���҇ڏz"c�t�9�EHT�D�e�����4.a	�"��B�S<�L�*"��`�9j����؋w��ZL�O�ݟ~��9	S���=<O� �&��}�{p�˴U>l�, U��k��W���8�Еn.ML�x���H#��\{I���Ңh�j<x�{p�U���B��
�������](�����a������#n���$I�J��AM{�ݪU%��o`b<��J�gRM11�t��
i��+�|�FT�i�&`�k�ZhR/���ܐ�CV���_�	=�s�4��_UF �))�+�e_{g�m�S����񑄆@bA�r �������q"��"��+m�����qGkk>�`	#�v�BZ��" ��W_��g�aGϞf+V�Y��u<�3�#��5�����٧ϰW_^K���ɴ�����ك���S�N�F���6˒�O�kkW|`�v]4w��r�;��3UM�MH�����~�� M���/�TsJ����D[�2��� �LS�ϱ�[��Z;Ქ�1�ڛ[޷�y6w�bF�3��d�,�6�k�.	S;����ښ���T��<�z�RT5�Y��X6��G��i�P�nY	���1E��7�� �7i s�x5��-_������S�ȵŹYvŉg�s��n$�y��:��ZfJ@�r��HA��Ҍi�� ?��i!o�d;��9���US��L��h5G�n�����N���;�=QzxV�T�+@�w�V��GY_o����W/	5qI��V�Joj @���d­�֬/��[v��0��K�̵,\v��.8�����`0�*{�Y�;�<�xZ̈́q����V�!S��A�*Z>�C��8����v���]kK�Tr) ى$�CC(�w��˚ Fp�>ķ���vV/:�h��j���"��df	�ّ�����r�����~�s�"M$7����n��NZv���w��;�o,ho9���=l� `�ҋz���޲��z�������ڸI������t3r+sp&(BU~݊��-8�ln`H#�y�n�%�hš�#��Y:H=��ZiA�)2X�;>�a�&�s�jy��d���%�Ok��>`���?�k�0h�m�.]b��j��� )��pPk��5A���m��n0H��<Ad�>��1�CM�"'���ԓOо-���x��{ޅ����A�rPT��M�f�.UKnx�D�8��Oki�Ա�Fڇp�tHw@�b-b��I�ȥ���ȴ���޻f��$�(�>᷶�T�%�Sqz�S���?JB���`V_����D~n<����6�&���� O$��
�d���l�mG�����I¹s����m�E+7=���h�T<���W���|��7�H��4Rp�f�c�����D���ߊP����!&g$a��4�e+�����J'���x_��״
�T��ò�QZ��"���&Dh�a�O��9���l|�St�~sr/q ����<wY��,@�/����S��|q����'l<��vb�d�������f$!S+qljӵME�"�|���"��$��:V�O��,rŒ�3���v�ڿ�+�/!���>Z�PV��ʙ88D�")�	�wP�%Ʀ�F�&��4���<��@���C(���>��j>�!���K�ʵW�_��>^��(&QK���{��u���� �e5����k����~�$�M|0�Mx+�MDr����N�� ʜ�!v��"�މ$��>J�ťHB���������Ap"�!�w��Ǝeסš����Vӄ�3�%!K�:6�LL%�c��T����e����9� �J�\h
|Yia���؇�l:$��%���%����<���6PvȺ�C�B&��0,#����/;���d%�����30|�-!�sd=�TS&Zm�k$�AԉJn��XMX�h`�u4����d �7P�o�TaGqӉ�p��s�|`\p�\�2b�p�!�=~�v
P}
m�m5�-��H������`���4I2�c�m�-�d�z�3�H�gN��X=uQQ+���߁/�6g
\!6q_W��e���q�VՎ�!	��K����5H�7*;� 䇤�%Cj�-�#����~��,��w��v�������i��^aO=�O�I��#1M�H��*�:�V�_&�fwkO�������'�[�>�qx|�u���c�>�e,�+����%��N�����/��LG �;�{��S�"�yе~�[�����.�k�-���COZ!��$H<a�K+�'��9�=u�x��3���H�8�$�E�>��F��G�2
��ߒ�`�+A�QH��=W΀�H�F9��𫠃�@�|T��Y���}��Xd�D�T��"AN�1��]xıV2y��]�C����*�Zc7��Y�飏lɒ�m}Y���_����l^�me�Ӊ�óy�%ۀ���8�u�'�K�8��/H��p�5�D:e�.t@�^0>�J'k?۵<��L��	b��OVZ�A=CzO��B��Nd�� Ʉ���L�m��_Xa߼�*��߳?��G�k�&��/f�T�}���Θ�N��~:��'N���O;���o��������/����`_��ϭ`\�UU�رp�J���aQPUSšI��{�er�
ۙ�@!.7SJ�N�FM,j�GVh�܋Tl�RH�c�Tl��ѥP{
BV	|��3�:��)ڂs�x��Pܽs���CU>��^�U�	���$.؍B��Ʌ+6���r<��C6焹��ͺu�N;�3�H^=OR���6hEw��Ƣ~��#���`t���0��\�&\B~uߋ�bK�e�������J�iǝl߼�s��d���\�Yo�����i+τ��>X�Ӟ�=�-��Ч,�#����G�M�ċD���8_T�MҨ*I@"�ٹE����G-��l�Ѳ���@u9���	�Hƪ,�81�X��o+�;�   IDAT_Y����� ��⋱2ir����ψ�
����*��)F[�l�� %&���d�H����C��:Evg���3rP�≨�1C%���i�Gc���O1��e���?M��eG/b�"�o���Or�iɔ�fA��N�'��w�sF%R(�?��ǚgI�?�_�en�ߧ�hL�_��Kv��A7 'G�x�ui����J�)��c�b��w�ڵ=��%欻�v���?�*׎�H�����Nb5�W���kʈ��g2EL��_M��O���ו��o�Sk��ǶҎ�E���d+W�G��E���.�>��J�B�k�f��m���Ϝ�i��� f(�Wo�k�ll$$��x� ��Ree��d��W�M6H��q���� Qn""�Z1�A%1�W��AiS��T��\ٿ�S���v�W�y�))S�O�](�p�=J��F�H�2,N�@�a!��M��_�Y�T|��t��>Xk}���~�d[��"H��$�HaÆi��W��!�j������;$�l�>?��z�j�r-�@��T���4�i�T�dRK��pкh���{A�� ���@��#�fA*��M��5�����,���v��_�A�*��.��|6w�=��˴�y6�t�q�i�v{�� 2�ߏ�!�=3\i��B�=��{煕v&U�T�DV,_��3�]���>8R��q��I*w�߄�<ȕj�f��ڔq~{���C�-���đ�� �xHӗ�q��7:
��+�JF�A:I4��S}�|2f ���PJִtYV����E31�	 ��!�{�<c^�Z��&�<3�n�����ϴˡ�݃v��ۄ�Ejqp�F�2�ILR흷Vآ9s�ۿ���g���=vܒ%�bCv���ZAI����kv���v�9'!�8�&_�0����=�#�k�\{�)p�ZF�[��Ƅ>�d����Է��!��c�< {Z�J$5�'M �����㜲'�P9P�!��.��8~G��UŤ_����-ꔛE+�%5a�;=1qz���P�h��1�g_=��E0N��7?�kb���e�f�d�6�4�vF����o�N=�"�������R&c#D�.1PU�j	���T�ń��WQ�#uy�����"�o� �F 6��L �j@���䘡��$]c�<SO!�Tjd�q4Y��i$��?��~p�v����^�і���N��Z�q,5d#dp= ��B}mׯ�q��2+�˱?��O9�GO8�����^{����
���[b��5mٱq�4��<K�hJ�k�VZt�C eUu�ւ�Hs:|�)���/dC9CܜÇ�ĳ�
Z�鈆J��Ok�t�����l����A�H (�|����qF��-��ڻk�ɧ���A�z�!F���!3��a��z<>�x�}���=Bq�ʫ���A�t�6���2�$������L�>��vtV�S����~��;a���X�?�D���n+�E!L�5igS����=����5����_I0���K��w2�{����n���sHj��ԉxO��.�mi�Zf�ٞf��Z��>k�;h��\���B��8�~�P������9��Ω6c��x� c N	LR�Ç|��eMeY��~΅�,xo�Z���9�!W�!O��!W����3�ӡ��������9�1=�5(��u7��}^��M�e#?��J��-{%?�a8^*�9�%���j8�O?�"q��NY���<�m�ʙ������}�'�}ݞ{�C��dq��ou�Eh*7 j�,~�:3C�q���3M�cn���XJ:��3Xz��l���x�P/9�S����K5��Q�0��$T�œ�PR��h�@7LQ�ʳ֐��!�ߒRRGb⒠<Ə������F1.gB�������&�@?j�}՛����_~��$a$.��t�H��\\�:B�w�f���N�T��j���	� �O24��|b�x�Е��cQ"t��δ�WN�MU��R�NU\\��V¥M >�������"�9n_Ui5�.������B8��z��Í�%@%9]Q�Gё�i�J֘(i�� ����$��n�� ��t�G3��ZnA���Nh��a���D�;���VMgo�<�7H�ǔ�?��=T&-p��̠� Q���O9��\8�2��A����
�y�@;L�sɢ�{�`L��}��_���qLO^r	�2�<}6�B��E�(=2U��~6� �/�N;0`G"N�KY{`S���!r���������m3��m{v����P�U�l`��41N���ηm�����-hV���mUC� �!䅼1�@�W�'p׎~��`��]R������@j�$@h���sf-Bn�����ߙKYMup��C#��,>BΗZ�
v<$�1���>��wn��Y\߽$��+��p��=�-^v$������7�5Z�w�;hwf�N���+J�1�u(��|��W-=6�I�T�' ���s��'�# �j�	�X�{w����Q��IIG$���>�Y<P?�R�b�Nn� A2ğ8
�^��f�$ZL���\Ϻm�RҊ��/k+*�z"��Z�h�-�[˭�t�����,����M�h��@s�=������e��#��oW,����0�/���i�Vډ���O�:xEl`�|I�Q�� ����"��K�$0��*��b��C��������aD�w�� #�J���$L�/H&3�OKS��D�A�{�d����͟�ow�z�͘�f_��O���áUm$�<�4�ƾ�{�7z^_S���WVi�v�8@�x���n�b]���#=e[h�^z�ivϽ�[Ai�-��}�?���ʦL�bI���PHv�ؤ�_�h�����/an��\Ŋ ��|	['U���
Z�LL�_�&��@v@��u8�I�ቆ*A�u����ڸ$:!C�� :�9GI\՞J�K0Ğ�k��uvΪ��R�DW�jJlb�p���<���r�A���r�4%'������2� i�&�@ZEh	���n�H�(�z�4�Eb� '���*H�s�^1��s�`_K�[RD!
�N����;�S�<`��3�<��8�4K�p�F�cO������z�G��J��ְߺ�T^�Dob�t[z<��$��� va|�Os�����v��g���L�h��g[� �����΃HWdMc� յ c
�c��]?Hf s��>@���ɾY$��q�ϐ�B	��Fg��qHJFC�'��֍�^;2�$g��� 1O^C�n�~���u~�b��	�����n����������uklǙ'��'C��!Ξ���Sϼƚ��^l��_&��ݳ{�e��6���LW��*qo�]{/@�%��S@��_N	H�ӡVj[ꓑ$Nɗ�q��]�Z�r aF,�ƄV=;�\�g�K_r�������C7/�J���B�X���#�ő��`@B� ��GD��e��J�nRG��g~�Ϝ�	�S�u$>4��.�E$hY	��a�T��;���)S�R�Z
�-51�!��n8����K�&�h��Dݔ�)�RKr˖-��Y@�
�x7��oQmȲ@A���0	ǚ����^p�Y��%'�F�$�������� ��Z���(�ǵ�8��,Z������lm��R� !�����i%��֧��V	�[
�Aн���?���	���K&�7������b�q�eM��b�w�I��,kF�� ;[S}Gۢ�ٖ �{��j'VX���(��b��&Ő�T��bEiqN�]$H�r
8p8,2R�'��~��(�KI�Q�m��w�0V�eg.]L�v�(�;%/FMcM�BM���x�i���ԓ��>��An��o
0��rk��P��)����j�$0��xdf�_
؞�CI�2��e�ѽ�!��c&�O�K����?�ǴX;�n�=e�)��h�8���� W"O�Z �L�&�2��Q��s�$}��3їB[������۾���m)ZC����kf�˗K.��.��ZkmF� >����6����cbrd�[�t�����u���o���xf�5ġӡ���"�P{8xā��d�[��� hJgg6�C���@�$��)�bQ|����q�{�5�t���K�f�˖��� ��pp�8�{��T���n�+18��| nc��Λe[∣�.��"yO%D�C��{~b��}��?�6}��r[8����L��a����C���{[I��+��qc�j�5"τ���9����4�`�%y�� ������j��`Є�&������M�#.���Ӡ`�nG�w5�vS�%ۜ�GXkm��0Ywσ���%b�m�!&}��*܇���HiL�&ڏ~�;��Vn�_�췼?O<-;�v&�b�m�<��%�澹j�}�_��{�^�M��cm��yX�h{��r�Ƞ��O�����YB��.��wZ8k�M,���XO��	�갭۰���wJ�8�L|�:�&�HxA�I��@�}��a�ҝ�+(H�XH�����~�q�u�i�{��7{��4ā��9$'�F��b�s@�T��ZZ��sm]���y�i�H��Y�+.����żp/(}|�.x��d�S0 �����-H�4X0�xB�l�cG�Ź�;�v�*���l�؄�#�҂�A+��V�_z�%g\?�d����wY!�+��uL��6�cL˵˜���o�K!�CAS�L��4V��"���������S��4<��+�&��V�����O�dK����&��b�~+��t?r*]�G�-#yt��련��|-�!���;~�fф��:��@i"U�t���G8R2,��tO���������adڤ��BU"�*�x��ܻ��:�,��̶��� zS�a��:8�=����]H���dx���1���o2�6�y!�0�O�Gi�9@�7ty��?��S��|�e�àɩx�~�[�֊��W�u�$�1)/�}�M�ho�R�5�J�k��j�J�ml<g |�pb��%������Mb����o��07QI�{���[����£ZQj�� 	RE��@ ���d+�#�< M�t�B����^��r�~���t))_&�n|��3Xݪ5)��1X�$���ʔ��G>���ipͺ��!�R�3������ Q���Hu[_Qi��'@̶��c�*��'�11���D�� �OZC�|�� fΚ�A����@�!���?��.)x����M����)E�}

��N���ߟ�0*��$�z���\�Y7��&��RO⭧^��|��[���ͫX� �'ܿ� 
�v�ыq��G;��ᲝT�$�X��d�qu�d������e�g����i���4LR��ۿ�	n��2M*�)B~z_)�:��B�����O�f�m���y@���۲K��҅���iI�T���{R�|O9	H=/E��A���_4GҤ���CNI����(;�S=�R9������iw�Z=zg�1�B3GC
��I[	K���;��B�Hf�7_�[#g���Rwms��R�k�LZ6�H�����B ��JSG�Py��w;0�C��rZ�"p�6���}NH�q�N�N�I7���V�o���0S�	����j%�Vq����H�>Dh�ȪA��T"% o���[m>��qn�h�����s��%��QN�\|<���_^����SH��Xm=w���[��\tƦNV��b����$�x�u;Tq��� B��A;��x���;��������r��>Fy�ت88���}8���^d$A�u������ ȧ
�!��nDR�x5�ǁT�q���T��`l��?�O��~�%jum�{�$�id$Ij�i���Ɓ�44TYVj�!�� =�dG�x��u6s�<�km���$�h����ܝ�V�R
 Q���E|F�@`O=q�]H2��~�Bf'U�>-,q��x߸op�t2��_�I���Y�5�6	Q���{$�L$�D/fb2��:B0��EK�������䇻��(hŤyGYn�D�PP�eå$u�"(�g9ʁ���N p�ɄyC�O�Μ��Ө�S�4�Ȩ��L�F��t�'�<�u�i�'�oK��:���MȄ='NQh|Y5�Ӳ��Aˉۣ�\Ѡ�I���g��$�x(�!���(I�xk�&��D_>���ҋ��{lΑHlW���S��&�B��H˴�h����#����'�Gڇ{3w��Xl�1��m�\s�a"ޓ���D|���hwh鄻(&Y��'�\Ob �����L,NsS��p�q�w'���r}�#�M�chZʲ�Q�q�Dl��9�L��L�Zm��:���x^�$6���B�b�l��MZ_*Z��ȶPr&�� �#�8�s=�DP�>�8G��5�΅F��G�ˉȒ<�r~Jwq _[�E�tPF��!��;���@	��Q��
�I]�]u}4eʽ�T�b��&_�@�B#��(��o�K�*$L�)���b�׉��K��H_(8��4� W��p.��ז�N�������6ʤ��wD��W%�v�%�OB�5���>>s�]�?�s��Ѧ��5�CM�a���
�&դh������-��&Q,�e�uu��=XP�$-W�x0�鰟8q�{}�nܸ�>��Ƒ�l�22j�  ۃ<�V����4I$>DP��*BU"K���T���Y@9L���<���C��֛pf�l������G���%�:>5�ߑ�k�4� 7ۉ�u�?GΤډ�Pr�F�069˺�At WFť[qMU ��7V��}Q����#���d1Li�k!고���Gp�V�JYh��I<9 45Ѐ��̒B�K�G
0����� �O��vj�v5w٬IS��������VB�`:�jr}�]��2�?��4��Y6�#�E��2��H1jǛP���/��)3t��6e{�/�x?�9�V��h�`<x<�^�@�L�MD��zT��A�:��5��3���
�ZI�[1X�ao��GT�M�!6>?�Yk5��xBm��L�y$�L�����'*e���f�xD%�l܄\����}ݶ�z��1}�ʰG5���ҷ��:�9����4";�;w1Mv�������s�;�I��| �t����T+������lX�1 $�$���Rѡ��|�����:x�� ��i���f�4"���R�
lݖJ��x����@�0kZ�|al�������4d���#����f�]x��~�<{��lR~��r�{g��Z�� ������?�.-�|�N�Ҵ��}�D��u!'�v����홷?�볋�?�V=�(	�u\���t�����5��u�0��u�D�<\�%b��C%�Dѧv��Duś��X�m�A�M���� {�������* UH�t��Jp@h�L���3f:٢q%�^�)�9�����v�:%ɲw/$}v���H��-;�>�2�{�-�7�Cpľ{�o����I6s�|�:�]���g.�K�_��yH��/��VZ�Y _�Hـ�H�a߮�.	+ �)���Cb? *�"�1��;x?	�%�� \�,E���'���磭~�Y	�bH~ˬB�E�E��8�!�d���T��C����Xh�^��x�n>�+�>����U%�a����7jgJ*� Z�8|ﳶd�>}r	��\$5|Ļ(�X�pNG@�S�6��+��Do&9C�2o&ɂ���p���pg�����{7h��l�A^�Y/�͵��>���(���wVZ�����G��'�9�a��ܻݎf�������o��d-~��+`���=L�$+3(K��)��A�㭊]E������d�!nD����3�Ol�]��k�D)Dݙ ���5uS�<g%*,ܴ��G��%{D�6��	5��W[RNq���@Zcj���I]>At����XHێ��k��e�)�9��s�ͽ�Z��+�Oڣ������܌!nʒ]	�G�΢]��ʻ�Q^\T4	[�$�H�5" ��W�5%/�L�֊Θ$�~'煺B�TL�{�!�H�P�.q����r�����f�胋�h{��N��
���3���ɹ������I ���_�}�$̑���DB��B��;�!K;�{�ӣ�u`�4R�)��QU���o$�*7k��8͐�Sh�,Z���Nd�3�p퇶m�6�	[ii�BF>p��K�Ƹ`jOJ8M	XA*)�dϙ�z�le���q� �ɱ[A�iq��,�#ȿ��aU�-�^b�$�ߌI�z=���&��v�~�]$�'U��k�wTׁ�5�	��fZ4(�f3׊W]Ǯ2G�θ��L.��ǡ��u-	���R�,h���'��w!"�Y� [?�'T�Gɕ��Sش	H�Ѿ��!d��PUɾ)�ꦎ{[�7^Xb:��e�	T
袏 �&�֣O8���Ԋ�py�I�HO���g��cd�a�BK.���@ⱏ�l7�f�2م�6r?�~A�qA�G$B�I]=hD)�c�<��U|z���w��$��gy:��R��ePA�5���Ҩ� K �.o<��m �j�� ~����	��p�b �j��*q�	��7^�9׊�E!|=I�ڍ�!8�^Ͼ�R� P4䓙p�I�n�G�7}�	6���\���/�j+W� �D̑ba�^�"��
I`-$��#�9k^��ܟ*ZO��д����9��='^���EaB�סr��HD��JQ����)�sϔPb����d����]�4��p��[ "��E3.˝��LMwm�0�� {u�qG�>�E8��rf�Z5���es�L��h��#gP�����ꏿo��Y`�@F�4�=sEr1�J��Z1��#���Q`�*���� �d�Ѣ�2��v�*�e񢹶s�Vǣ�Rk.=@P��N8Ϳ= ���o�����$�S'Mv�Z{@��y�jZW9 �A�jJV.��Λ9Ӿ���'_�[o8�}���	F3-z����$/S�K/D�Aܦ>�3�ء7=�"�^:�����f8z�<;k�I$Z�X�zoԈ�v�Z�,������z�A���A����n����z{��lʄ�ٳ��l�hq�0��+$����x.h�mX5mز���nָINB��}�!����6�]+��đG, I�2�Λhq�1��]��C���쨣�q��F������	���_�ٜf��v��������w����]�� -J�}n��8��ZiSHv���HLG��!#�A��V��h��b�hY*������(��;����&ٛ�d��x���%�����'�S�[7c�T��7����u$����??�d#�&�0�xH�+t.��O��x�͚?�gI�����Ȥ�;�g|�ڨ��_#������c�PH@;�(|%�#ޗ�s���e@�萰0�Y	�@%�eZ��Z`?�!�'a�%H*��l"rD�>�;:Ľ%	��xx	9�BRs�4�Ys��N�rn@���p��
�5y����$�u7#����v4�3��S��%r=aMbAt%)�0�����b�QC	J�5)+"?I����t'4��D,��R�&�v�i��-5�η2acIe�2��٬{F��k���ɑP/g'g5:�#J��C�~:�
��I>��!1��I��M�tKR-��Vu���>�wq�h+��;�S�&8�����C ���D[��Ybh\o��*J�A	�^���P­� NK+l*��v�Z�S�LqIY�j��E�E�=ɴP4��ϡ)8���$����,)�A��������N�w��G�J x��ܜ9�gI�Z���N�}ږ��
��X)�>{h��@x���3Hb�O� (QF$zP�oD�5T��`%�&�'	�o�~���H�i��b����O�S�x�����@�5�ײz^�'�ĔW�v��Z!`� ۦ����`�u��Y%����߉�-?H��丨`��J�&�Yk@9��
���q\�*�0��ס���i��	�Bd����E	��e�,�_)�w�����@���!6Z'�D~I�]x�ٶ{;�6;�Pڷ#��foJ��؇/�	L��}��<�z7	��r��=l�y�����p�@�H��#;P�*=L��<k�d*� ��.4��'��w�
8Q'.=Ֆ��29�F9<���K��Zu�ǲ�!ɔVۅg�D�@�;�䰑j���2�,ɏ����Wp�x85S�fҠH�l��Xsi�(�S��p ���o��p<d���a�{�ea�B�C����#l���!�M�w�8��w �������{�+ahE�Ν_��w�0*_��t�V��n{IVڞ�Z}VX*\r��m�]n{wbI�c?R�ў|��{���Ht�-�#'K1���-�8��.ީ!y����&�#�ڈ�7XGn�Jed�RҎ��4"OT�iI���4�7�~��tY��,�2�^8>}���!�f��OB��x����$���X�s/`mg��j� ���%�f�:���m��8�o���o�p�s|�,ڰhɑ�ȇq�K	��	%v��9��`��\v��y���_�i���Tx�g��N%QL��������y�\���5H���.�z�X�$Z�p���{AY�h�����cj<�}k���"���yr=��!8�IP"��Q����[Wk�}��ƹ�W�/�B̲>����Wf��/�c�_���\i+�Q�Ő��t���Yo*��,9��l���Mk(|�sp�j�T~xgN��v\��5mV�'���A�Tx��nF��~��hZ�jewpͽ|�8���9~��j�n�5�'�78�k���v ��P�^�Gtt*-��d��c�����نL^�٘�wso{Ɍ$��$>�<<�j��bq�v�� ���n��v{�6�D��YT~����vĜ٬m�Bħ�[�0�p0'#�k��S�������V�/�d�����Wޏx��L�<!M$Sq$^����p�3~�~�!i�u؇��������O%��Q����P|%0L�d;�c�5�$��ʸ\��^H�(ݒ?��8k1�0(�pihl����͒6�`��)ֺ�=+Yo�xQ"�ɤ0"�HHAi��{͕�t
 xt��D��d���(T�ѽ�^e����"��ю" �V$r%#��)�0�����8��XKw�P0�������~�o%a�A7%��_N�u^��udE�9$�� U�RsN�<�	�~�-��KP9�E�a� �Ru-r}
d?R%a�(**�^�ƉAjJG���M���� 0�����Y*����8b�h���fz�V�2�0pj4�A�8��G�����Ak���߱b��e�,�3U�|.e�0*�{���qL�e�#������x���$b�T��K�Ӫ��-1U	�rRX�l_h�2����y�,6Z��(�9j�� �[c�j�!��A*�^"�#4�'=��krw�%QŎО�P���C��a���U���&�	�$R�es�Z�����C@9��7�V#�?���{�I�zH�;� �'Y6��5-MmN���UF��$n!�6����D oC|Vk#{z<	�V��Fk�.G6r��}\�x0T��E%���O!VF묁0U|4�@�*�@���[
�[��QT�C@2-�$ ��j�l�e�B&�t��#;ӻB;���3^��`�5ef��x�T&ӏ�$C��I�f#K�?f^Nq&	�&�>&�B�U%Me..X^A�͈$"=$�5�N)���n���^��"�l����?���X���(�wu�4�,�����{�o���{ ��XL�����w�Y�����ۊ��ݸy;���v��oe_d���c�MŝJ+���c�""�J���5�<ی�Y$����#/�{�N���ESH���_XC�}��T�.BG���!��_�53���!E���#J&�<Yqa&�������H9���gZigM*���@�ƥ��ڱ�i�j' �g���Ja1w�xح��xT���:n�!�@A5�_C�8��G^�t�9�ٟ�{��;��Ym�d%2�����T�=��c�u�]s�yvԢ���c��W_�	$�� E_��;�����W�'�z�d0މ�^p��v�W;��W���DN���2x�Y��v��u�ھ�2�:y��'2p�	_��%'e7�t��"I[�z�����N
Vh� �c��Ҷ߉�"4�Þ�.I�a��5�^l���_��b���=<��SP�/��pC
)�TO<���e]��_�Ч�L�0��E��-�gz0w"R>�VB=��(>��A�\�R�"���&y��kSZi�'�V�P3gu�z�),u�K�F����\�īR��J,�xN��5p�b97��e����:8t�̖�s������R��ː��R��EmZ�G�E8�
Ζ>t�6nz����\,�๶R��v�Cƿ�� �Y�ƐW��[~�x:�JL�(ޛ
�1�!�5�g"�W�����)^��G�0�@���~4F\+���a�b]ɫ�@�����{i��#�;%κ��\�Q�m.���hf`*�g��5E�уPR�V��e�f$�%�*l�̋�P���3oH��IfpV�^�(��!,�D���#��EIqIW2��*��p�ԕ �-�����6sR�=���Ş{�9�Q:�ߨb ��3�%�=tQ��͡�?�d���HO	�Bo��D��r�Ã���{�F�`�HJ��/!�7����ٓ0W
k+���@�bR�2�'G�"djA�"�	֍��:N����K���`�Skic���V�F�`D��45�~^��v˂t]wD-��ӧ;=�ʦ08��:#���K�$t�6�*�?��$.$��l�dJ!ξ��ZO�>��e��5�O ���j	���>д�	A�\&M�M*��F���{l�]�oLU��w�d��Z@sd�!zAUe&����A�M-�(6i@�-���@_��ȤMF+���jU=߃�[��t�Q�DB�h�BJ>H�/�~���!4q<cxH�c<^Q^ћ�N�^Fԩ� w�W^yb�f�6~�D�l��iT�5�����rؽ��m[��jP��$�|h'�FJ��L��^� �n6�(�\*-�(��N�!�V�5 �I"Fی�YbqPH˝��T�I��D��H�9�D�����A(A��%����������C>�$�9�*�$���a�NRS,�@����p��j���!�S���`���]:�h��e⬍uJ��]J�֣�P�)�ǰn�֞8�d	�:�ZU��o%E"�k-�76�u����C�H�f��S��ÑAhm?�g
�C�,�@�����x���
��14qٹ'ڣ��믹��(l��#�w�_��0v˭W�?��zW#�1��m�n'�|<\�j;܀���K�Sq���f<$eL���q�
�`�q?�l��j��sH;0L���(��
sH��/o��%b.n�5><L�hd�$�����<�t��(ܦZY�C���Pe�qʼ�ū�(�|�w�O���}����V�k�=��'����h��8�N?}!1b�x��_|��8~�-=z�m��l_����].���*��
��C�o�� �OF��<۸u��Z��g�Ȥ^6ω��Qk=�w\=NDx�M�TD��d7]w���d���[��Xy�36�.i(�碫��e��d\t5G_d�bbI=(l��i��S�`n"v�ů��XQD�&y�2�����!��^~t���D�F|�T�NMc2�&�W[�a�Y�^�+�y�I��&Q�6�~�B}���e� A��a�-d�Q��O��&�	�/$q����A�+�BV-sQI�1�+�}e�S���V������4y��uW�"EznB��X�#����t7��۪��A���ؕ�T5�Ā���)�wB[�,C��YS����hMs��E��60A�і=�B։�Q�
M�'%�jѱ���"��u��_�tK�3���-�G�"Npf���	̔�	��3/;�н7��li�T�r>� I-�uu�ܟ(��ޫ�1M�zz���|) @����"vIM<�׹OB�IPā�)���$k^m�(�*���.��[p��P8��"Ʌ"�X�����H
tDu֠_	]!'1l�~�b?J'���E�����k��^B��~��	E�g���X����ធP �T�w0�I\9/�"c-5��I:��0Y�(/�����Պ���t�Q�i�AJ��t�)�!�	8�$��@�/5�� �k.�yքRQ����P{G��8 ��ϏϜ���F��q�a:M����?�/���u��+�r>\Q�@N�ElgG��b��w���^U�����ϟO�,����gҢ��MEj@c�$m@��F6�NN��u�&�m�
w���!c��r����H��a*�ޘ���Nq�g"g�Q_C`�ER�k�/�U�bJ&`U�c7>d�� -�`��7Ӓ"cc�`�½�x‍�GZ_ڸ⧥��k`�HI��.��L�66F/�$ץ�t2}�j���.�c��1�$��#�PدŮ>Gn
�V�&U]����3��i[p�r!'#QAkW������>�H6Hl�8�IX�$����'�B������'�r_�w��C����5І!1��$Tv8�u��ڱ��r���F�D�M~o	$i��N�4���dsҐ�z�,� �D���;��!/k� ^E��Rx����\���xO���J����M�-��Σ� q�C�����%��>�dX-�TxE�֬&�53M�UG����-�=��=����Gչ&x׭_o~�� M�F"�!�U{��NI��/�}�BzhB��@J���$Z�� �Of�Umn��}��GP_���y���I����B%�a !�Đ�y]-;	��Zk�HI�3X3�������h�w|ˎ�l>�zf�D��)�뮽
2p����?&��f�$�oF&p;�9�wl0�p`�Ar3�Pk�n��*H�%�Q�k�,�R���Ï��u�Y�N3|,	��R𵗛�aI�������(��0�&��m���-��7�B�j�L-ͰV8U>�W�xͮ��;f�D;j
����m;��t������el?2}�Mǂ�W�3)������a��a���ļ��m^I���Yn�<�G�n��p��3o�1�ώB�8���xh���[m	��G.�����!�I����V`����}���C��1�aP��e�����T\r4��������C���]�&kS�f9s�`*HZ��V�T���P"�6�\i*�#)�ڊczR��A���J��$�.H��G��} �*�rA����`Ӈ��$�	�?��M��W(=%��n���R
�h��r�˻S�#�V�RA�섞�gPA�a	�����	��z��4MB#k�A��!
�h�*J]ڤa�Hʆ��͔7�A�_C H�u���P�Z��_�!ΆaP�x�L�_ݕ�p�6M�����u�1�a?��E{g�VZ��t�� �����#����zAv�I �l5Ԅ�'�l/#7��>��t)���WW��{�cx(��7��n�F��ix�<KǏ?$��	mf�ƒ���X��#�f^l�x�"�K�����u����}���S��./d?���@ܦ�JE�g�h���<q�񠴋��'��D{�D�%�K���>�e��8c���7g;�m��yƵ-�)
��.�ջῦ�M�9͹�!��N�"ٗ�IA/;�6���
Q]+�(}7�:@r��y-�l'5źp�Q�����2���ѤMp�����u!fY8�#����tw5F%����w���[NF*T~�$L�T &
�J�8D����(����� u����T9���P�3t���� ?7�5(�:WѠH�W�!���i���5]"�z��^{�3���ׄ���%!����ດ�c���6s:$�6С�lj�y�y���)�G�p�L�SXx�d�0�-D�$D	���G�I�N�Dpt���@ӭv�Y<}�e�pW��C
�jʆ��O�k������ �ý�d��]!L�P���,4:HJ;Dd��&�  �L�E�I5��ʚZK��m�!%�P��~��OeU����.qXT1
�顚F!�E�
�!��`��hb	1���A�8�h�N�h�`mI!h�"'H�s���I)�n*>l��8:�Ls��b�K⷟{��&'��	��]jy�k��,=�vn7�LU���TZ������1����@=$�Q�!8O�� R�`9%��N����7����^*ɂ�>�SM���,�K�.�p`t� i�l��C@일?�c4"`z,���I$�Ꞑ$7#3�E"�L�I���'��p>�;ja%�P��ē�� Sc��{�Ȋ�)�S�q@���§ɫx|[ݚ�񯴚���pR������ ������ �0�i��ݐ��d�T�Jt챭ͥmX�P��5u��N%�X��+�ٲ%�~�:�Q�����3+��ނ+�˲g_��>w�<;�s+ӑ{쬋?o��M�z����Q��C<���D�*~>�nXf�H��� 9#�%�nYT+!G_1I��Y|��������F��rH!���Q#��iD>���Ñ�ig)f�
4�Vڇ﮵9$���fT�Vܻ���g�  �ܱu�n�b���-�95�~v�r���n��$\"ZH��s3�.ؐe8D2�B�sO�����mv×�i_��Wm)�#�N<�(�X,���d���{ږ�z�-;�(����Z��a�_��Mνb ��XxTBL�+��h�rI�roز�^��KV�C�ڻ�V�3w��^��.�FxJ�$� 7�Lr�}�v|-�w/ڂ1���A~�
#6���H�h��b�]y�nP����t�	L&2��Bav �������^b�x[ �F�h/Y%a�lD_CH�H�d��Zt��rЦ�z4ÓS1�Ѳ��iDsKr6�	N$$YXTu�eS�Ǥ;�zX��"�tڎq$M���D�b�bT_��Y�d#+q���L��_{�~��?���<bǟt�m)GN�>�
!9N(��8I�71���Ja�N2���r&s݄���2��W�}��!T ��E��Ȑ�u?Z��\��u_��m#�N���J���$LI[47?��"����G���� q[r�$c~bC
��}���Օ�fE]�nb�����ø��Z��I�=���V�o7��Ϯ����y �pL�m<-��c���d� pK�����X�aϗO��<�z��^]����B�q��Ï")H.2�p_S�q>����0�v �p!�		V�����%�T>N�$
P�!Z�:�A&H�g�����@�>�8o:�սꡃ ��8��d�}m�, k�C��lE#o og
VZ��h.1���տ��gN�#1p��h1�*p��c�E��"�;s#� ߐB�J-������eHAD$�F���A�����x� ����m:"�"7��G@g,E�$4~"��@�mBÄjI�>?���Sed��@����9̊' �G;q'��"'�^�/F��@D���/��8�_C�$�X�OY^VA�l�aЮ>P�Dd�����Տ���"�Ʃ��A�G����aA(�����M��Uo���J�4�\/S]� #�Lq����َm��[����X'2���|?��MN�F~���I$� ����is� �Z����������:�޸{�&jc2T�.�6*�_O	�|�Z��UB����IK8Xr3C R� 2L�qَ�i��II~
�6'B��5ժ�-M�{yI7�p� ��w �w�U=�"Ue%*~PSF2���QM�Vc�&�֭]��+��&�F/��0(� ��̅[H4OZr,�S�µ���Z­�csB�Bh��0Ԓ���W��}O�k��"X�O0o"�U�Br%i o��;��h����U0?R�C$��<���R&r���`������.�yO�U!�v��à?�ϳaM�wo��TmY݃V ���g{�M��0f����OZ9�,&��+ʬ %�^~�;�n��G�o����|-�A&�`��R������K��O1�����x3�0�\��٫iO=��r˄����$�A��SK�T�T����6^tR\�8Z�ѽ��i኏����1�z�e���������.T&Ol� ���h
&���[�B�o���-�d�}���nd"�@����������,{�B���⸗:���ynK�KAǄ��I��BI��zޙG#f;�t����� X%��0!;��)�4���z�����Y��dPf!�;���n������!��y�X���D�0:sX�#ڨ�.��Y����BX���	��Ҏ��"���q��&�K���B�T��|�=be��ީv���*�z��5;�[.�4Ci!�E���n��t��9�9]��O|�+v�(%C��ζ����S�;$x�	���pQ��^�F"�'S0��y�~H����C��#��,�]��JO�X���Q�L����������{۰a=�nk��>ں�f͝M�I�WW��{[�Q���m���'[�)��U�ߝ�p�.Ć
��[����o-�<�����3mrA�M���CR��Ԣ8�tӶ7�4�����*������}}��T�p:~��¼�O���߉��>���J�cH�D�q2�Z�$S	tC�)�ƍ� ҇t�����j��Z��diO�3/�<��,%��G+1V�/����3BE&!:ݵ0Vmݭ��᪷���y"��}�2&�/��z���r�'ik��Z_q Q�ԃ$�������3DߐȞk}�F.�5�� @7�� ��G�3�K=Y7�[5(I��b��9�bA8IB�����C�^R�VW�9ZD����~��4�|�#Y��{~|�$�ӊ�N9_qV��.�����xa:8E����o��g�A�
iL=@U'�|I�WWb�h>��G/8��Q�W�]�n=���N<�D�IU�uS���k�B�Lpk�X�r=b��+D.����nE��#X�~H���QE !s��c�3�i�fz�,�$��d�����Ck�u�|
��IsF�� �TQT�P(����)NX�� �fQae�DzOF*B
�C��v &�X�q6��*)*����Q����|�(w}�6 �Fi,��8�8D� �J�ju5�@�����Z��m��s��+�������V�o�h8S_��vDӸ�N�N��&�J���߼��H���B�T��p_�$���:h�����l洙�֘�����f�� ��-�Z@Z��	�ڔ&T<��TH�)p
Z�����H��c��;JR�F�W�3I����}o�TSP�S�JT�z=H�a@��m$%�hHm�p,�s/8��+�j��K,�U�3�q��6���4�2��P+;P�{Hwv8��G���ui�tDzJ�� Ϝ=R6��Y,�b�ÿ�C4�*���0�em]����;р��iCm�8�b����x���𾫵�[���' ?��EG3|�q�^IG�4($���9��v�xG5{���Y����V��x��� k��P�l;�S�y�c�J�
�̏����q��~��<�|I� 7�)�F��8 _{w�����^��QQ�Cu��q$}��/���5�/��JԮtԎ����Qk< 2*�9�/4�
3���p�0��
�J�p�:�N;�RHeU]���z=6Ms�����x�͞S��2)��ar5��*��� 4Bm4�)]���x�j&���-9��eu��z�-/��m�9�fL.������M��؋�<�[�Q�ʺ�],~�z׭�Y��M�9�i�4|?�X��bl�L�Y�$�*t$�0*--�hr���q����p��2A���D�,	R~@�����P�q�q�8�Y�~�&����*��>R�������e�Iy�iW�����H�A�أip���g/�2M"֥�M�~�y�^։$Z�o��M�Vq{��s��@Zȇ�m��70���6s-����T����"��[�����#g�}��P�� 콴)5-�@i"a(E׮��L�۵�U%�Х��Ƌ/����qH�3T���S��[����U�0� �K���S"6������k��M������a�>��%����^̜4�.8l��F�� T��#Q�l���Ci����V��$Qg�+��ti�+)��	�t�3���l��9�����I1���c���lUĀc�[l'w�sMx�ѿ�a�(b������m��t���V� o�(�.	�_S��qt�b�(�}���+��^sb�t4���Q&͘n�}��$`���kk�bqd�)���P{H��:e���#��7l��fI��z����łg/StQ+$�����?a�-��i#�h�2��%i��qO�H@�i�W��@��%��u�ۓ��L���� T�)�X����?�S�����!����x�E�ԡP,�Vqg�;�d�[�,N�L�z��VȗA&TR!��=�M��7����_H����h�fW��V�P�%��Z��M�Bm4�ȟL�hEpdD�a���#djҸ	�˜�f�H)���׏U�/S�$�(e\K�U��/_es&0�
V(�?��~���T������D�la�}6�#D�11ZZhm�<��뮸��e��+�xr_f͛ko��ܚ��(L��Wo�N�|��a4�NC?9	��C2B�I$��D� �'@���g��D;�@j�"z��X��iS���j����Z9�j������l����������~p0���w.�S�BS/���
�C�!�c���-����פhm4�yS!�/��Զ��@[9��ԡ �N�wSy� )dI�!�M>�1w���ЮI�x����8�WI�lt��{#�j����Yk��'O����Z2kl�Ν��>�G�?�d�PI	��˫�B���'[>�]��d�݊�e	��/�r3஡����*oA�n���v�}r�>�����4I,RSN��d(� ��P�cZYrP�Ub��5=�#@'s �����hWi� �餢q)���[l$������U���@�*@VV��d)h�$88�0����Ӓ�a�>Xg���{�A{�DƏ�pϑǟlg�}����a ���Rz
c(��䱎�~�)�)F���V�6NdH��^��Xa� ^�i��[_
�>����Z��t�&��#�\�oD�xP�kCc��"*c�| "vV1�e�0H~x�m�}-��hj1���{��K��O=�)Ǘl�4��|�ٷ�W7�V�B�u��x�-[3��Z�.����8<ѾCJd�g��OY'�ɾ�����A'6m�i�����/����G�Sm����$_�=�ȓ ݽ�e��U�ԤC��d��T�Քd:��!"�u��B��խ(��u��������;��d���>�����d�n]o�-pB�i�u�l(��;�\hm$�)R:�6�h
�+�bVO{-h.�~$�i�B�_��;+��U�LM7�u�ԅy.���s��%'�(?����H�lM��̵��z���SUm*��۰^:g������0�9��M���K�\�>��[���=mT�N'��y�n���E�ژ�.f�~01"���k� ������yB��$��g�r��?�����?BZ�V'�Ok����֏P�ZP�m��)t�8+�ae$������()"�Q��t����>�@΅�5�Ȑ����y�%��Q�ES�O�<��=�4x�M�'�6}e�UU"��sJ�@3�P����^�{�n�&[��;���84��0��سs����=}�U����O?�Y�M%.�3Q��{�Z�m7Qxl����->ǹ�2sqc�;k�M{v� ��I���co��k��土8���mg�����$�Yv��D{SCh�\o
�ѐ&+%�bP�v�{q�*$�HȆ(�b8cE�I$qa�G[~rZ���Sm3�����Da6c��1[����$,��9�H��>�w�����Q��Y��� [/�*`�\)H�g@Z0ln!0���c5��FLW�oO�2��S]�l�޽v3Xi���Ƈ�������w���IL��;�)�^*��[?r�!��Πɶ=����=�Xx�&9�zl#�Y(�$	�9.��Jj�˙�H��8�=��SU:��&n��!�(�q�z!���="�aI���ß�m�l��Ɠ��^��Z!�^u��������ކ�,�Wr3-�������t{����܄�{��>���h�;�ڮ���0�dF�t-�ô|�#h�h$�k����Z�����_[<���n��p]�3��#aɅ���N�{�{��IrT_�׺�,��b	zzm%y=�h-I��_	R9��s�d�خ�R=�8d>����%BАN�D���;�pe���˽$X�\�,~pH�Ҕb7r}:�5F-q�!�U���T�!u{\�g�E6��dIM�p��s@HwNvgG�n���a)�o��}~��g9DD��"��b����ZH��X_6mr&�a7��*p�	:f��f �*��4֨��w<�/����p�����SkڹGp=q��J��N�i�l�8yZt�V�p>�m�L,�2H���$�8d�A��A)�B�8��)<�����W������)BM>�=䬶Y�^P��3�D&�$���^�G��p�Zkԛ���<��h�(�gP�ԁh��9�~S9�H"�G8%�J�|��ߢpQpD��A�vV4�)Y�謂K"��vH`��J���E;��������}Ś���h�4�M᝷V��s,s�\Z|u��?>����㤤��c�,�*�z}��X͕/$�=�fL�2��
X��&Aj���g�|�D�Q�k����V�A��s
	�Ё���.8�4
�z��ǿ�3:ŎX<�>d�cρr�㮟Yɤ	�s�^�y��W�3Ek�������'�&�h�!����D<8w�ip�hт�lܸŞ~�������=$��Y�r�

�We�,� iU5�%?�C��!�_�H�ۑ}�ĮD0�Bw��u<D�UCV��8�UAdpv����A� KX[~�A�_4Y�i�z�ڴ#Nr� �'Q��ĸN���xbng� �׵��Σ����e�����hh���?������W�
TP�]�؉���X-2�hі]�u?�x�m޶�n��&;��(��c����1"Zi_�d�p�"�q
#�h�|E?E)���t���j8)�^'\���C�6� �j�= �m�Q!���)����Mb�ޝ�}@(���C�Iy�ݚ�R,oECKQ$1N:Sz�*4�z%�d��Y�zi�79��������S�JA.�N��Ѩ;�_1	��W݅�W��G�}�ŇP� ��S.{
Co͈��@rD^�A���dr#NYzI)o�����+k-���	�4��]<s��bust!$���B�E�t�	��Y��s�{Ь��ư���roz9#dc�&.9Ӊ��倱N�� 3��C�#^Ϗ�/��[(�3'a�wK�[�]�!�5��Wj' �ի���>H+"��(1<�)l 9�����~���Q��6MW	��?�����X{�駙\� �T��%k����t�,ȿJI�T�KJ&;h�ݷ��N����^��˱���˒�tK�|U2�$G���:����tM�up(,� �K�\�*DO:1�d�k�vS'ծ�-�1����K?	���th'��oCWKb��/=�V#���s/�5_�j�s��w�qx�!Hk��N�����k��f:�47��^e)xFS��t�N��C�P�����4*�7V�&i�o�w���"b����bI�h=��Z�!N�,x/uܣLA�#� �Ŝm����M�>G��IV�Ij�H�q��1���X���0��D�'Mb�����z������#@�:ހ�p*Ux
I�!S����+YY#��� >��u3���u�.i���6�'�����޵sο�Y�TSE�6�8@�`��A�,���hG�)
��tPMV>���Y�� a��<{:Ӓ��64��U�-�e���<}�����N�G�sNsM�7( ɀ�Ɗ�}�>�DY4A����_��"4Kx��/��i���ZFԐ*�7��џ���x�F�u#9�ׄ�|�|T�����$�⤦�����$Y2�?��%�x��3��˺|�����0��N�3�%�Fx���
��(j����c��I�0������"�__�+)j�NF� NP ���~�Q;� �%��A�{'h���dt�B��9�p��P��#9p��p �dN�mM����R�!٢���L�&��6�e=z.���P{sp �K:�!1��[o?��د�g[=��pz�C�ҋR�$���rj�������3)˵�{�!��c(�cSu��_�,��~����pE�B��k�����ԅ�S&Z1�JmĨI�{�P�"�Z[���{��(��01�O��$b��={H�CNX�z?/���@�t�H�|P&��:���H(`�8R�.|pj�K.(�!ŗ��[����r�e��]�h_{#U</��}=2VuJ�9�At�K����}����=��P�(��}�R�W������,����L<�L��Z�7#����N�t�7�<� �T�F���$ֳ��0u���w���iq	�N�5�US���/�O�V]�E3� ��(�NRBh=K���D���E��~�[�7̂���k��)a�
m�k<1�O��a����Ԅf����k�*�$�Z��\�̈�/��x�$g�qga������)�(��t>�Y%e�Ă:P�t~WqH�V-Ff�� �@�O%af3ؿ�9?��]��vE�yȧL�<R�F��_1���S&�kh�����6��H&�:1q\9s$�_[�>������L;�K�_L+����`j:�fMkq���;הUѺ��WN���%b��%�(R���7L+���߾��6A�@�/�	�t�ĕm��?�6�!A�81ޣ�L͒�}<���M8�3����$̑�Yx�o�f�4�S����#�EձP�8��Z�zDz-�0��Bp���lH}��z	n��(���*�~$iq�p��������HT�� $E�L*�QD=�b+�3����/C�����:�^-<A��P5�I��} ���Sg�����r!�&$5��P�!6@���ł��x��P��\���!bdZ�*�A^zPEpyZ�"ˤ����1d�+�!b���WY��S��P����P<���(�C�3I����b4[��j�I�h�����q'�$V٠*�$-],�_}��m��+/�Ks� �i)�N���M�:&z'ٸ�T'��z%��f�	��SU���!E�D�A��V�~&�F�W$�	$E���v��x{�M`�������7��
��M�ݠ�F���󶪔� �W��"��^B� I�������Q`Ƅ��!6��F�m�w�6�9��9X�ᭈ���+ܴ�%����[$��O4�7�~x�����ܦ����n7f�����ӑ��3,�܌NQem\EЃ,�9���i�Q���{���e�y��7]���&k�AtI�F�Id�"�p��&q�4�� ��р�1��1��� ��A���^���@|mY !	���Yc>�_8\��}��7A��w���/N���"\;���CT�JAT��Q��E�
T&Ń<�N��	r��-�Hz"�A#b�ϵxT���$iՀ��+�������q~u�g�]�a����1$!��|?�E�o.§1�Ϩ̖�+Ș����lg+ǃ0�]�w����~������:�E�޽w����1� � 1��DJ"%+۲���䤫SvI�dY�J���E�b� �af09��t�q�޽�>��{d�ֽ��ǷJ��P# 3ݻ��}�{׻��.�)�u:鴛��F�����T4�w�{[&h��~d0Ӏ���+_{&��mJ��]\1���bOXm�@Tك;@�����>��tuv���� Cڙ�������Kw�R �{���@��<��S�z��{?�n=t+c���>�����K0���G�:��s࣋�#N5� j<;Ɵ���躂�}�8���E���E��>k�a	�b&I��{�ϰHi)����% F��?�=�s�m�<��q�bc�[�~�OO�0�v��Y��c�^�P������z��q�j
��́X7+g�	�w���$qo�P�r�,�����P
�+��V,l����MgL�
�z緽������ `�<�{������xW���)?c�V#�l�w��.0퀆:�6+ ˼�|�W��� gq`�,��C���諯D��M��� Lף��s&㗾�(gAkz���� 	�U�m(�L��1a�V9a&s�W�x0%aYT���lG�0������%ʲN�(�~)+w�}���9w��L�#�V W�}<������%GFq���X7pv6 ��yk �Bc?I�b,�Lo?���.n�HtZ��mf�_�|ک&�p��q��������@&TDVK}҆�Y��f}����L>����֩,�(��s�뛑9Lc�a3L3l��������=�Pa�q+Xd/p?�4r�v\H5|mCc��V��Zd�7�s�V�M�����`��p��N�Q�T��Ƣ�ԧ.LVt�ba_&�wSh?��c@��+��Әy�~�0~F6����F^���80Ņ����"�<dYJ?1KF3 �e��9�ZՑ�!��FL��Kq ����
�};���px��� ���@�#|�0�6}�����9�~G��سa5�����!��V��Ӎ���G9�]T9����2�n��Ϥ�4�����0��G?1�n�����W���:��o���=�,�����!q��ٴ�C���d(l�qJ&=��Qk';7���=�<���qZ5l`t��G����Q�� �@`�t7èp ��~��~!��nK��;r����o���	������Q9�"�ԚMo|��ip�n36r8EkSA�-b:���k��?���= ľ����T���fw^v�@�!�)@�!�b՘�<N�_�=�n,�tR��Ug@����<��p����� �Y�����W���F�2�H�/�;�T;w�����o>�U �)��a�p�B�ZIS0�t�q�^~>�H���}�؆1�|����6l'��)U����̡9b7:����>#��f��ξ�X�ٰyG:�%��Կ��	6�AZ%�fB	�����`r\S=�<��-�ڕ�`g���X���h`�g�U���n�Pc�2{Q��F�`��.�6�l�������{8�6L-�Y�	�r�7����w-�Q��O�����wc2ٜ~���I:�}�?���K��sKz�/�������G[y��h�8�ګ����?���T�?��Wө� 8�h}�s�x�]Lc��Hcb=�L{�ԩB�k�X�5W)� ��gb���~���L	�uֳ}/C�����`�dG~��~:t��X���t=}i�n����G8D-����/�/񻋲�3@s� �f�*{&�$��69�Ȓ��Ʈݻ�q4�^��%�Q�#@�]�鮜&���^��$�,E̢3�Х׋	���[�n��wE:�\��t��-\�Z��#�@D*�u���!�҆��ͤaa�2ܟ}�Id���֚�D��Z����mF�{���{���v��N�X�����ґc�9;���ɉ+P,>�Ki���k 띟��?Ð��c*;AW�c�輊�ʽ��1��G�*"���_�����>	���}���g��p�w� ��gÂ�1XY�L���4,�	��ř��$4G����;��F3�H'�Xz��c���\����/R�z9Ǻ���E�M�|M�e���0p>��@���Otfbw#��u�q�y�k���,�y0�9�ѯ�{5Zq�ߵ�5�z�l��e3@�g/�fa�X $��n�RbraR�N�*��N���`t�d����<�� St(��qm���A�	-��z���8x���`rs���V	{�"	]�uU�@�Ir܊d�ۿ�-����o��o�|��d�f�1��V�nC����
�P0^�tAn��>���O���<��5Rr^$�h,4�
�t��5�i��[��G/�A�U�@j21�Y~����F��:���ade�:P�ع�;jz�Iٱ{G�E�~���[�2�d��us�� l�æϕF��,<��f	���b5��T�<��5�q�� ���n��u��$S�"���*K�D�_�/L�B���G�z,��9hf����S��X	8Cmߝ9~w!��U8�!�0�eC8�C=�Bu���A�ˀ��\<}�y��ϙ���J�d�l5��M_fN�car��"��l$��CZ���v��a�*3�tR�!�	@
̗x�����*�mO������>�.6yW��2��	�қ.�x-���Q�~ ������s���q����Z�����+/_�A���Oq��#��� �1�
[u��/�z�Aʗ8�`:��ttEՓ�Cp���W�~)�up3}�� 0��l�9gK0��2*�NH q8�z�]N�H` s�?7�n���üKʯ�F�h�ހ��e�0Z���)Wa��5�/2V�2�(�k:�#J�cŠ@}-[Go{����u���Y�		�a�������$�(Ao���Թu[�q��('�`�B��>�<m�GgW��䐑�k�~*������D}O8�\����1 ���3k���cd����M�:��N��ZZr�����a)����h&?e����'����Ğ�=�a�6k��w�Sv@o|8��T�|l)��ˊ���ñ�=|̽ Y9��h�h���{v���G���q�D(�/����[�{ގ<����G�O���)��v{o������w��oܙ���8�x�/ӽ����`�����,��"����bR4��N/�Hk,��[��9� f��$�A�����c�X���{oz���N��[���~5���Nx�m�\v�� G(W�I���@jOU�1��9�m�}�8ԧ�B��K�^{swL� ��;K�_����a&���ׁ�=�`�������t�A��ҳ�M���y~}$�G�>��ë�qS�0g-�E۽o?�@u�BǬ]t��93�Z���=���9*�M"�!��w@�w'��:��r�3���v���[&	���H��DV�W@�)�L� +��)�wS���g��0T�������M�m�g�ħl�ß�'�4��_�G�~�)�[�d�Z<0�����c�)1�f�?�W1o���s�%Y�6~�4`f�U f����ߔ�c��͞iE���u\W'�R닟��?��d�9��H�j��?5��.��$�y�I)�L�e��]��v��X�w�&Y|v�k��^ kIOy������w�xk-3V�!�'�X;�c����I�2��~J�t���$����F��j��J�)�T՗�eOz�����&�p]|��'�If�s~/��v>�W��T�4�v������K\sK� kf����D7ù�����$�'V���B��w�l���GC��Pvu��,��cUK�e�w�sb��-�[_����9��CT�V�5��K0�T���MUv��>�4���!�[!b!:@�˯m�f&��j�]ņ�l� l+��:2ſ.`�cG@~�8LI����*�s �(�0��2�B�/������2�c��j%XY��a�J��6h�0�"����"�RI_)@�]��2��_�ֳ����J�b��@�a����`��]M?�S?��l�K��iC͍��D�Z���8�߅N�E������id����S����H���9u��a�Sݶ�zJ��s��tz���{Jw�v8=����e(*��MkL��+Opld���>��Ҧ�pǰؼs�t� Rj�D�� 1}l�Y�Dz�a�����GlHӣ�����Ko�+H���ֳ�
�ϟ�<��8ڇǇ���4��8r<�f�P�>��r��i�m
�;����D�A$O�+�=���s_M�g��fL�JQb���	P&�P�Z�3�)���(�	XT�@�jPR硸X�SG2��|�����ر3�Ư��t;����y�����t����ˌVڼq+A���Va�.$��I��Q�߆����w��`7��>��/������ �iIUaH�6 @���s��[�^�J�m�#MD(fÚª��qr�����Q��fT�EK�����ɞs���!~Hv�T)�p�(��K-��q-f=gRoM�Ԅv
�ø_#���p��2���2���vF��!����UT��*?�}�9[X��Х���*�k4�<��9������������X��O~<�����k����?����I����CwH?��M�0T��_x4me�}��;����7�g�<e�.Œ�԰^�(9E�'#+�k�>,��ukz	R�{ӻޙ��oI/<�-����?��.�x�lz��K��y�5����'y�W�}o�?}�'S�q���{�4�a�4e�k��Q���x�����^�1:�7ܙ����V���~s�A$��O���]��><�5��w�;�[7�=)fn���	c~`�^bȞ4�T�7 p��Ś|���?=�`�e���G�V�U�0ŮS�f�v�&�����&���ɖe߂"s��4�E���}��l%�l�%�%vϯ���1k�Zi� P�tn��l�]�p�I��w��yN�^A���xt�Z������I�5}�wgڻ�FΒ���?C��"L杔����#�h*�&�h���e�[q��<���z~tӠU�����0���'����_�|Z�}~�) {(��tb�o�sbt
-)qe�h�(u�����QZ�^�|��#� �
��j�vI�ԯj�ʻ����pX��ž	3�s4�]�j���bhh���>��O��x'�X��L��NVVK� �5���?�I�`����:�"e�Fb���˾q�$�\�S
2��}؀#�ێAw���(��������Y�	5v�U�$�u��9��@�.0��c����l�����m�\9�B]�3�q4��QnZCz���8.����#y�L`�W7�<��_���T"�����"�}���i��Z�
�1�f{���Յ��h�b�|��d�
,S���̏,s5!`w��ѓG�A�4��,Hڬ�d��
?��C�㡻�9j���/�[T1fq��\����[?�`2� ����1=�pt:��;�ږ��Ԃ�S�u�	�Ƹ�F�1j�t��FFɴQ��b�j�ڍj�t�4���V:�}�{c�r,h��p�5c�`� [K�Ӯ���1O�>��F���E�gSst��ca��׾���GnI?���O�q�t[[h4p$]^Wh%�ي�3Z&H��ٺ���6 �����oB�{G��p������lx�6��Xj�����i:��~�{��3}Ƿ��Q'�#�J����LO���,E�<р��=kF��0{�����],��U�{��R?_�՛w�aR8��m;�G�2�����cUg'$�Ҳb�R��IV���߁�w���`�$s���o�
_82q���Y��h�>���H��u(4Y���_�>���+f`n�w߳}��-*C�/�#�h:;=�6�����E+5m����(n����o4�]�Q~^�y�d�md�/��0����V޵��^���*H�� @.P�� �c�uP��ơ�jL�:�.IP���q4M�m�6n������%��˙u�T��� ��LU�a�̚6({8g=�쓘�'H��!�d�p�(�MV�h��`10n5��8|�������u�A�&d����lc�Գ�w`�9�&��������u���]�գ�]��S��QD�_Nod��Ç/]<KY�1J:v��c|R�Sr�h����Qj��g�D�xY V��y�����=�\-2��i '�~��_L?�#������gB�T�Z�?�2f��+�����!ڔ~����t�Bc�9:o�ډ+C��Q|�,�aR��N7ߣϝL��;������Ʋ};��2پe�)X�/|�������KϞH�q��ɻ�	���Xq0�K?��� �$����ŬW�W�X�-�N�~o�tQZ?���SH��6=�#���Y�6�I���6�QdkĿ1I��Jl5��٣u�l����
��&��d� ^d-+"kxMEbe�����y��
𳵬�;9G,���&��?����owL��an#�}��IJ���ṙϓ���uc?3IR��E�gg�*��Bا��
�d�3�qC��ɻ�Ko�Έ�/�wBۋ�$����t��O�>�J�,�<8&Fh�ۘ�9�Ԣ�2B.B�0������U��F�&,��8�(E�G�b��q�����������v�*E����I��q�����t-jG���ORy�a����n �W���Jk<��N]
Ʒ3ۦ�.��jϱ`5=Z-��g1I���f^��6��1�f���+u�j�#i�5Ļ�Կ�uoi��f׳��:�\Ӓ�SQ8��s�'���	~	�z��'�C̱>@��7�4�Ru{h��qp�ݡLl>�ֈ}uT}V���\a��Z�J��Zcm���_7��RfY�*-�G����++M��C'��!��ǐoK2`d����04�dA��Y��V<�8W��A���R��D�|i��j���܊�ey(��q�(Z��F��{���3x�>^<b�[V��Y�
�[��|_C�2�p����Ws'�\���I�����`��z��; ���ɝ+�LIa�eK#f�h�|"��z�:	k�
�P�<4!���a��C��b���)���_���w���|���S�hpZI r���g:Z�A����0XM�)e��#@}��K��s#t\���aW �#�<���{��ߌ������H��[7�I];� �j $�l1��Xt�'��%CTO����"P �w �F�d�ξ���a�_�l�Cs#�`5�{� VY��A��B@�>[q���-}�.�n��:s��XZS���`c����K���2B$Wab��3_�\��`� �˵��%J(���1j�����CC�2�Y���s�q�1�z��s{��������%E��D=��d� 3Q��;�d�h $��z�%���/��ˬz ��BU^t����lFɡ��y���|�a����:�7��ͪQ�Ö�4ղ�@�l_M�)���1�Dɡ�1f,a�Z~� &J��'|�^_�������s����2ƥ�rkZ��)�~��8���v��
�(������Lzû�Ӳ���M����O�����L��	ۘ?��c����ksoz�Ӕ��]�8dh00���n�i��q�q=B>���k��	J[ֱ���q��H?������W._M?����ӯ���J�)��w<���=N����� �o{�����P��5�'��l�p2�k�.f��*��SxZ]�kP�"	�zY$��:��5,�`b��У��)��!�a׬����p"C:c7-��)J��w��Ҵ6.&�Jv���ܰ�!���E��^���j}�f���|�<�E�Қ�0�#Y�S(�YN�w�c��;�6�BS�@��1��?���Y��3�Xۅ%�X���ruX���*����R2�M�[=��s���i�A�S:�G����J��X�2�����x�  S�;�nW��#�Lk}R!�1!��Yhs�}oHcM�3ʇ��~�����S���_�B�1��}@O0#�S2�<L�����.bQ��k�D G2R�kl�y��;f��<\�#�Q"q�!^�H�V�˒3��631�	=�l%��L�Z�{���J�����1�2�`G���4����/)���H�%t]J�L�!K���;قtb��e�ޙ��3������=wHW��T^������_ȷ�1��P�h����e�5(���S��.�H,�./.`_�䂵�:rL�������!�Ab�]��n6`��oP�Is�$;���^0z�*!��[�����M�0�/ۛks�j���P�A��@����i��U�t�*�R�0�yc��ҭ���������`�Oh�WXS��;��ά��{��-���6����Q���M���(-���DgTߎ���y�]w�2ӲcgVم�(5�F:�Jdlͽ�u����C>�%�/h��EsH���6�)*���<ժ{�3�r<<;���w�y�o��`�  ������z��_�C�}#�24k8S��[��w���3���l�_K� !Н¬��7����w�������tR2�i�p�����錄��!;mM��{��~��Tz��ߙN���;����%J�\�-��}C�kPH9����Pp6b�!�M��E i�'��P!{���)���v#i�p��FϨ�x��'�8-���� �ʪ%��:?�y�赤�͈�J�ek_ ���_|!�;��+��_��s�?��dG),ݦUD=� e��ߎ{�<�<Z̖����M�~h�|O7Sv�`s�����Au;�4 �P�<Qa�[Ҭ�Dw�{@��{)8c�E���3E���6X
��:��p��Fާ�L���L]Cd���55���H �p��I��5�nRc��g{`ʂ��)�>��f�2���2Q�4�a����L�5V��cg��U��C��}s�ji»�#rf|(��M��ї�K�oK?�c?ʡ��<˯���7��������.�<q-�������w�G���>�մ��Q�:�w}��0����'�NO�����Ke���`Ł��}�Lik|�>�<:�(O��O)�<SK�5����[����a��:�u��b���p_�� ��M�6�_���C�O'S X�d%�\�}x,�E،&:?�#��#�{X�g����
���5�&֝$[C��c[;���hz�5Ǆ}��9N`w�-i`-�a0��dK� e=��Y�&om���Gq�������2�%o7-���c���A`�#dl�/������R~dЦ!ȯ��L,V�p��4���ʚ����}+�w�څ��Q�_��R-k���=s��L\�Ya�5[^���Htf�E�l��`��W��̆�/ߧ_ ���3�qA�5l��A,��HىZ-Y��V��q5�OO��ۿ�����A�|��_�f*8H  ����O��%�Z �ФD��5�֊��ٷ#×����V4�����k ������*��*b
���7�_G��D���>:1gIdg!� a�K�!ی풜F��.�-K���6Y�씮��i�&��,�]�J'�fG7e����x
�<�ߊ���ksP`�&aR�x�=$�x׷���0�~���$�Q&�%)G�׼v�r �i��E�f�<�Ԝ�j�vnf��.1eflM"��� �2q�YM;Ċ	��-�1��uO���]<�V�.��3�z�FR�DW�<������T�kc�/�u��A����R]��B[S�*[%��X���@�y)��aC@��z����]'�y:����F}ܩ�0JK)��x�B}��$���0�%, �\ۧ@�]t�UȀ�|32?P�������+0�2,�S�_�՗�B������F��+GO�O�K�����J-;RCw}���9:�R��Nm�-��<$NY2�!�7�n%�+rX�ԮrX\#��ro���C�BW=fܰ�{�94n3�`P4;�S1&�'�W�(��, tDY���)k�n?�O�lsڪ�nP�k��zr<d3��\���Z����_M��O�d���3i#��iƩ]��5� �h����M�[)���k��s�7� ]{�8ƕ�Va�)Q�Gqlt�s8�P�o��K��J�hd�Y� ��s|}0D���8��U*�[`�L��j�]x�����iy�+��YCy[�E@��7�N��VC���q��&E�<��t�6�8����~�7��?	xZo�Eas�հV`O�^=p&'��L�����5J�y��d��e\�y�e~�3�%��Uܛ��KK2������W�$�|]��L#G��JM����2�7G%�`�����y��$'�ZK֎���
��B`5&�7�x�<�
�8rVY9b�2�lu�QZ������{K&T9خZ:�V��ү�H	����" W�ni3G2��*�u��賔(?h����y��.�,X�Cd���ʿ�����~�eXI�([8w����oD�w�$a,�=�j�	G�����M{���Q�� �eLU�<�.�J��/�W�O�q`��ݝ>g�Ѳ����|)K(dIr�
���Q^��Cj97���4�7m%vi�2�� |�Xhl���&`�Wi�	SD5AzV�\���JG��6��u�C��]�y��歷�D�$�5��G��C���^��`�f��!�}��a{˔z|�65��v��]p��KWa��~`/�}-ɉ�{�&�1��cѠU��0�����d @����\��$K�S���@��h��y_�=�ϓg�jْ��	$qP�U�=�5����LY]����0[m�[���ߚ::땪�̵�h7&��5�ͩV����92ɲ���2�6P	��4.5�W��$��. g��l��G" _Z�M/?�?��������t�2����W���t��w��2���nR�l%Fi������2�yVM�m������Qϙ��u���P&����F�'Q<�mgyV�7�}459I[�|I�q�ĩ�O>�5���	v����JsMW�$�	���}۷�vGҞn�0����U�=�ӱW^H��&n���h��&c�I�,���؋x&�umƦ�h'�@(���t6p���~�?�ۦ��R!�����+�����s'c����@{�����LpB��i�����5�e���g݉���G
[���̊���D�y��h�ж�P�:���Ճ�,o��5��
+�4\�x>V�Щ��0�d��ՀH>	koc�[���͑Y����0�
�yIvH,�vN��%�|�٠c�%�{Y�@���rԏ�xc�Ȥ�գ,�!���Jvշ�� ?xna(Mx]�r���]�-@��,�=� �w��ml�4;Bͳ,��}t�T:Ω5���҃UQ;�������#�moؑ~MXa1�sxO�S��*	
�̄g�iV#�h��څ�B6��G�����^~�O6e�Z/�eX�#l���� Tj����X#+��MB8��%mZ�lĝx�`Xa󷲑N������ޞ�^��F�3��̥�!zq_>r$�rǝ�n&��,ो��n@Z+ϡ�Nk�f���18�,3l��78G�"`B�� �H��V�� wP��!�@��T!�����%���}��7L�0cR}x�9�ʎG��aE�¡���驀X��h�4K]p���I������C/�L��8P� ͮNKI�|�����N��ad*�S�a��G˓v��6�(z�O�&�J�X�>�^�v�oExL�'�KIfR�0��5�e��E�U���8���i m�ҿ���Z�ذ�*�K7 �� � e���Kst�i�a�p�$V��e~��	�U[Z,0@�ϝ&��ܻ.� 6����3�ӱQ�[��fƜTʰv�W�����`0� ��z-�S^p.�%��F���������-��q�47��%�+�o�#G�d�j��:CBs�A��1�qzzkɰ{c�~~�h\,׸��8�.��N=;�ט�72NR�c-�l�g��f�a7uEa;�|���\�4��6�`Fa���w���b�]h�<pe�e��M
�Օ�yf��$�=��i�ۼ�&C'S�^F��S�Tf��j��(�#�V's�O6���4�ܸQw{��C�]�>��8��d�?W���-�7�^�*ɠ�����-�����U�e��fv3M���/c	k�=��ts"�ؾ�/ƫ���c1�X��Pv2�D�ױ����P�(��m�`��J4��o��p^�#�- �4e�@�q�4-���}]�U�y�CK���v:�Ѻ�	Tg�
k&c�t�Qg'����5�j��]#��nO��@���QJ���  e��������mn���3�]�|����a�k��3���n}�Ж�{`�7乫�l��(;�S�LY5��U�_��D+A�\�*	�	�q�鍌�ж�N�afhN��a]�x^��,�C��8�_���؝XZZ�,z�1K?��Ho8�;u�\T�6�H���k�i%���e�} ���W����a�-�i&��[�_���w�!�g�R����y�g���DL�C�1�Fd��\��ٲ���y���@$L����$��"D	����CBE�ų��8�B�F�y'��v�v�!�h���,dM;%������ݏq0�Y��J��.8���a�0��R ,�"�v,�Ъ:6{.�&Bl8�ayrt"m:�=m�o��\�ř�u�x��8$�ԍ��m`f�frS�J�x��T[��[��,5|X�1�(��i����O�#���>̡Z�������Ш=[ӓ��80.�1��N��Hg����̇�0B"j�v`��B\��2�z�ܞ����������;COq��Xz�[��I�J�������̨s=r0-��� >�ߺ1�]̌#�ѡ8~�3��r�8$/�R<F�!�L� ��|��R�F����~��<x���["ñ,���Rӹ�#��nF�_��N?�^{��8H���w!�b<�c���J�����S[�^h��x��8ޏ,r(",'p-b���r���#���Pv٢#Y&�pn����l��=���� y��}t�foz�;	���3gɨ�a�.�j�HRSJ ]=�X7��.�ڦ�=&���Q� ��CJ˳ �Gk����2��#3��m��>JY�:�SN�#m���= `~��̼�6F�����H�u��Q�%�4S�C����Z `ާ�ӔS`�MDQ.��c��CO/:�I��9�)AX&� ��C[�y �����2M�\�-kAg�Ҏ.ΟO;�k���n�f �g�k�|�!\�t�qu���]C�<�æ�nj��j��� \�g�j�s��(�����Y� ���̽��������M[�Ӊ �KY�n
���-ߦ��񳂞�L��`AX':��4�VG�F��(x�M0?z-�!�oFKe���/�	��4k��a�g���c�R(�e�T:����^��켃C��W�`'$�{:�^X4��,b��Q��E�qj�;�Ѳ���8$w���H���'�f�����U��20h��q8�86*����Ĳ�"i�h�R��d��k���k��yo`�&u������7J��\ ~��i`�Ɇ%�jS�l_�
����ژۦ�-	��u�/8˞�+���t`}4R.��-W�5��_�Kb�1M�`��exG��	�M ��}�*6����b?��w���⛖I(e� s�w�T#� �����Nd!�ь.9Æ��k�.f�α�]�vb�`=*�N ��o�c�����ձ.����yi�~J�N�XH�1nDGx�EA�{C���{-�.J<7;���ְ�T�xZVӌ�;���Vh�	N�X`�MP>��z��44�� S��oa��U(��ٕn�+�����k���NǼ�6��eJ� }�q G=|W�������-���,`����,����6��+�g;�h0)aB,h<ɤǯi��<h�=7��5�>���ؚ`����s/�Cw�S���H9ѵ��^���vD��)����?�E������~��%יeٟI4�G�6����2�փ�8N��_���$���sg�7$W�x.Lg�T�B�"^��n��r+�ɇ�,����k��f�:�גѪ�X���O~?u�F���EƑ����5�J�rU���\.(L�t�	�Da��9��6^?�rR�#x���<�����nt�P^Xb�H�Vi�ޏ��Yp_e�|������QA-���p��ք��vX��]���j�ta�.�� ��Z�q\��~��f)��}�K�s_�|:s�thz��S,@�����#�QO'�0���M���k�O<�}�.c�"-��+dL[�1����ڵ���c �Gf���#J��/ �����������8��� 3��2�3����[ɲ��]b�X���e3e�96��ׯL�Т9O�w��m�A��<�hN
d�3��
���G�Q��l��>d��V��H)���c�-�u����G��8��r0f2/�YAg���͕�&P�����% �ѧ���`g��\��Xo��_�TG�{-����slF�2bS�J�O�~�Z��e����8|�p������ ���\f�q:�;�m,7¢��	S&�0�P՞�4 �\X�~�hy�w~���� Y
��&�a�z�.�^�x	�3������eN�L�5���H�$��<�N�|Q��	
�58���J�wn���
�X������}��-=5���ln@ =B&>���X���}ξ��Y�<3[GF/���������	�%��N������j�*ߴA���Ж������ii����>��@&̲��q��k���ϸL�.=yhR:YW 1�� �}Z���S����`Xxeѥ\!	p&*�:��n�q�������&֜��Y��˯��O9�"�X�o�z�L��j6�8�:��6ިT����l�v���wm���	Xd�d$ʂ_�Q>︋qH}̇��<��Z�Y�9����5ʚ� ;�=��I�_�y�n�_u���j X9=�!��3�ޡ�?���ڽW��skw��>JY��W^�>ƂMJ0� �2ų�s���.� ʢ����!kkS��`��p��to��;q��42x:]�t�)L5�"3q9���p�_ N�h)��M 
�i*�i��~�I�}���_E/��}8���}����Y����h�D����X}��,p#gM3����d����y��������FƄ�$^�\y��m;=��-0D�L�\�%�u�2y:ʳ��00���ӏ�Q>Z~8/Q�S˞�3�����氪�K��#?����o��}�	Jʌ13aC��EI������3��g\e�MJ�����㏥[�{�"*��u�"�/�+�������o����^bz����1}၇ޜ��� �:�W�/����g�.��u��	2�/�-�>ٳo��D����|;���>+곰�I�2�� ��A:�_xṴ���`2o����&��o��s$��5���LP8K�W����ZJ��9�gJ�58{�����݅Q�%�-��g��肉fyEĔ��*�oj!�s8 �S�4ǡB�+1�vVc;q��Vs;| �Е�������Ifj;��p�~�dL�%E�j�TK+�s��ow�T���Љ��"��0)��]{�O��_��m��'>�Xtn��FK�$DW�*��]K�ԯ�d+KѢ \���5}��^JA���k/�+�N����f��/=O9����{�H�UD�ZY������qx(Z�g�PLM�JO��!�|��X�7����<�:��*�ؠ�('7t��Q&\L@�G�V�LA��	���n���³O��0�l�%Am]�ހB�������C�e?76����ݏ>�g��v�[���W)#ܴc�,L������+h�G�7OO][����qD�5���:Ã̲l�β�#�<X{za�Va�p}6�A\d��+ꔼ0n�Hx�Iܗ/cŁ�z��fgM�{+A���e��֒C�Y?��<@Go/u]�Q'�N{nf$�f܍���_�1I2
v� ��ݼzwjy��6�v���Najx0��ѽ��i�ZO�*yx���%J��g��^U74 �p�%�ưr pqᑸ�a�� �e�� y ��� �
4[{����Y�}w�gGZ�%�=�L
P[ !���>���9V��{n�˫6]�pc���I'�*�c���Wil$Q�E�Rϳ�k�>�Zt�ɼYZ.&Hn�1��0vs�I��
�`ls����+�)�̍��П���5�pԲ��ѓ�t;���:�p{��.�Q�Qܴ�6�� 	Z��bv�I�+%�9NGp��|+0n+qU;G�R�$���6M�T��%�������$�T�e�\'��zcKʓ�4NY߱Y��a�����c�����iC?`��0f�5�<g5Q�����Y6m,3��8��b���_g׷��&X�Y]Ǵ��1����ͳ)���^��'�@���D���sĝI�# �l&�F��U� ���m�f���V8�a�,�����e�% ���+�����
��J��+�P!����r�� ��|�E�����մ��~�99y�q�j@];�	�V ���\D|��,Cƹޭ�o^�GJ��b�9���Ҋ]֬��A��,��<�&��9ǅ9�xr��	1�q(�s}�$S�M�t舲>���_���ĻmrN*�{�� ��6މ��A�=A����p6�^]N>h����9����-�:?��Hrd�'Uǅ`�H`/1�n��I����g�	���E|=�K��=K7C,�K���Ă��-��B�1��G��0�1e�p���	�-��}��G~�G��s^�<��Ϥ�~�����N���Ϧh�����4�����k�r6���L+�Nz������1ȹ�X�q}S|���5#+j"b�V���U �1gV��&'de"Eȋ$�5�s#R�zbrɄЈঀ�cS�������AXX�X7�^���ö@�.����ъ�R�n^O]��9Tml>����hkmC�ȇNG,�X�* �&ۄ�� ��S�1��������(?i%��y����Fٵs'��B[y�c�� A�>���-��S��S�����y? JM?{��2��: ٜ"��2 p]�Z�8�^���x�`_qe�%�~f:�Us�����P��/?�N{)J9�Ю���@�l�Z�]Xu����8nE��Z��}{wl������Ⱥs�<�v����l��EZfk�'să�#j�p׊<@~�#\��v:_��#�����o�s���=����hK�Bca Y�H�ɫm����� CY� ][ 8o��ִ�l�9e_%�>�|wڵ��@�G�C��rh7�L�m�`���n��1�M�f2�/o�{�.�8�'��A�p��4��▣�!0�Yb��
z�*繁�Y=Y��� 4;����﷓_�<ā<v#�ؓ��`d�㰸�64wMd�����@�<�Rg����� �F[�v�&�e��,?;x{��M�����?>3A��H�V��|/+tv}f)ړ����ݝ�҆>&'^ QG-����e�QD��t���l �ļ��h 8�$n�흢����v���N�>�D;ai��كC6N�X����4W���;P��ݒv;����@Z1�DC"���>{�{ý��9�ޘEw��%h���SZFY<��������jv�R���=s&�mc�δg; 3S��q�]ԇF�s��q�E�k(j{�Al�G��O�W��,���Ϋ�ﻃ�e'�>j ��N���$1Z��)s�Z@5ak|�렅�=C�<�E�.f>���7:�$JO���I����?4)�I�C�{��zsF��-�J��w,���ը�}��J}�s��a��T�<%SY`;ߚx�����<��q��F��a�w�޷s@��iY��ҥz�Ϭ�g��#�=� xk��2�h�C�a���_Y@uy���m��0*��`J���=�~vM���t�$Y��2kz#F�5u�|��C�X-���4�2Q�������҄Q �4�x'(��p�_l�����%&�t�aw�蘧~&Y\<��g=X+�:K�v�k�����a�8�2�T�u�B�z/ >��G��ȟ��`/��������ճ��j����RY���@Z[�b��UG���l-�a۵%��H6И�>N_�5<"5�e��R��Mjs7ɱ,��3B����8*�Y�q�}:�~�ἣ&��mtTv���N�d��}�Y�{L#�߷s/l�Ƹo��������5����1[xw:rd�.�� {u�_��S1I���Ucm��}i3��a�:��q��Lt0��v9⏘��t��ڮ�����}�)1&��$E�0Ш���`�Y��=m-Խ�1]��3I�o�K�rl�Ue�\�f�<��wG��0� ��N��D��L,7���5����吞������(۬� 3�[p}��na�)��D�a�g�ŬI`c'�X��ٮ�6��=�r����}9��'�s���"��-w�A�h/_YIg�>"�2�����R�}�}�Ƣ�	Mݛ�M�0o,z�4��h��T]��J�5�v�;���m1J���T�ء���ӿJ�Ǿ���!���J+8z�`�������d�9/[��P��m#3(r�մ��xe����!���O�g����c�3���}���l�"�\�-�L47v2/��KfŦ�lk�Ì6��A�8e���g�6u=Z��a���t���n�Q������1���^nN�Q������֬-�@�@GrŌ �»D/��8h�:��u�8����vv�`:��Vw��Pgt+��y���.-#iEP�a2KF8Ai�����^?lv��6�����D�!B��ZV��i��߮��>c�yנ�^1i�֛8m�E��m�`��r}�A�Z"��D9�Y�v3��i#!�c�_�W��q��Lj��D3@C{�v�0�X{��-� X�Uk��Z�9/)��N�PK�# W�'f���f�ف��n���e�]��3}�xe#T���X�c�����>�&v�7�� ;��	A�/����ph��^��bI#[ny~�2q*�����Z���P�D��DwX��9�c7�������pس�e2V�6X�ۣ���s�L��Fe
���r8:�����.7j���H����qpWe�9��-�rK�Y�NR5]tޭ*�W7�q���w��?���_u~a�ag�L'k�&�z����a��ň$�dK�r
:8l��#]<��A�	X|ٝ�}G��5�e˧�^ �g��Z@���x��<�N�c��i�dl�@X��Lv�u'��.��e]�`������ ;m9��S�mqJ�luV6�D��
ʪ���d �=<ͺ��F� V�U�F�f�w���?��n�]��d [lJ���W�}����J�Ym������6��^�CX���7� ���k@ge|Y$��U�D��w����K�cj��i3�^|6�l#~I�����]$&��%-�m���rږ��=6b w?�g���
M��G�'���4�$ͱ���ft���`3��-6�8�{�{�9�Z��2�~�1��'{�Ⱦ�gr���<�U����U�5�)[ ��Hd�����?��S\��Rh�JT�����G-��N5F|�H��g y��U�K�r)W�8j���1��e�su������,!󻑟���]�Jt������ӵ��Q˧��2�1ʼK���6��z�CL��v��G�n�D7�y��ie�^���ϭN/���ݑ�]&I��BCAwl�4�d�Z��D7�S���� ��JfְF�z�gi�v�Y�� ٦��C�XR[�E��H oB/�a�C�e=���c��Yw^FRG���5@ք~�����e���g;�1@ �א�&#�2�Դ�kwKw>ws4j�rk��sm�4J��kg������[��H��f�#�qH�E����0�[��	 �OL*zn��IXk��d
4=��(�Y"��l2�_;����>W )c�lvB)���{���f��R�-�y�7Q�n'��^��ͷ�i����i�Q�q�vz�V���`�Ǡ,<l)|5��X�T|:HǍnѝh���:���<4�f���]f�ˆ&+@�j"Ȼ]�ŬV��`���;p� ��!��{�����Au�h���^@�4	�%XՄ�����-�h)a�z=���������8B����HW�ݭ�����x�`@�m�(W��kN��HC�d���ej5�c���`b�����Fp��Bؔ���9��kW�L�YtC*�6co�l�恸�f֭��I��S+����:��M!����.[����'�8�P�n�ڵ�oZ�KT���$���v_dg�	�&�����;�ޙ3��pY�����	��=0e���h#kF1p �5IKAK�#���P�Ӕ��!����)+,�5|�L�ϑ�/z�z`΢�T7�%��5���Vo�&��:(���6"D �LQ��J �Ӄ�bW6�L0�ic�$X��$@�s�djd�(���,��z�DΜ:V��F��h�g�;����Z�s^ 8mZV���$O @��f��X{,F}��Y�36 �.Ȱ/��aCa�ZBH�VIo�%���Om$�[��p"�
Ih]��E���0�Y8��+�˜N�h�Y��u0���s���<1n���
C߀���%���ś�7P|�b��?�6ѽ�	k��!��8��ǚP�P�i�E��I����RQ3��I-�ή���T��ղ�R>{��ܑD�y���dA#g(Vm!��2�4�x�J�����$�0�ug�]噶������gRgb�����&�t�ؓ=��xٿ�0�6h�Z��-�M��-��<�4��U�p�Я9-�ĳ,Gv�������������Z�_$F+������v�8`��}����E���$!���Z�,:c���v��D���<����>�f�:OS�טU������A��]w�ƹ�$k�%���#7���LI5�9b��sSx �qn��5���i��<��:�N�V���X��T��¬�i�ҿ6�w��5�}h��l�و���|"o�˿���ط�ER��<��.�_�����ׯ��G�JrjG{ﾽiP|y�V�;�*�<�v��_7]�T���2nvB:;KCV\��x�,�(I6�}E�x�z�,�w��ΥJ��Q��pjڇ�hA����4<=���SnRhJ|��%jT4�[�v6�5к���A/ [�g����m���`$Hy�g�����������Υ��~��������������Yd�Bu�^�C�������v:RFӱs��إ �>h��S��6K�e7N^��u*3�N��nJ��ϲ ��P,Yo�zW ���-l�J|s0q�L5fܾ}3%��0�Ěc�@>������N��Cn��8�F�A��)��A���g ��Y���;�OK,�D�.81�2@��r}��_������`c8W�Z�S����j��`m˛���F�y�*�`��v�0�A���6�q�����R�����������f�Nt_}��Q*Slۉ�<�9Խ�ؼe�d+h"���Z8�����(��A/+��;�.�����ذ�Z?Lx�z$�8��8�|6�������~W�?�?�m�u��8��漂Aq���?: �,�:7&cc� �r�]P�������#��6<N�����0��M@��o����\�̈(�I؝�?��~�%�M]C�2F�����kv��8dNM4y����sC���f.v�:R����, ǚ�2����J�6�x��T�Љ���8�<Q�M�c�l�@|	f�ò�='��v��1Z�P � ��T�Ҩ;�D�a�4�U�=�NV��+yd�k��fak�	2�0G����He��E����u�{�Nƹ�2s+��E�.�p�� 4�Ӯ�w؉$���d�̶�t�6HV�n�.,�F�h!��m�I��kr6�(i����NW1퍒Y8Kō� �q���Ě��U.˴��H�1D:�끨�+�x�: i�.�^]�јȐ5�~<��MpR�����L�V�L�]+"n;�`.m�H4[���؉X�cE9�26E��� ���*���l�
�X��l�C�����d�S�l��H���tӮ�0_�5Ei�DD qJvx��A\U�w�niuX6<-h=�}9�{�[^+��d����:m-�Q���5-6D�!z5b�{��C�:��2҇E�c2d��oY�"�X�$[V�I�b�2`2�Pܣ�S�y�$��q�Z���{k��'KX�s�l���s �i-m(�jh\k���D=�Z��۩Dl؜��J|~ɡ�����3��3�9'=C���w�<]5}s�׈�j���'�I�`ۺ)��1�`��)k����1a��q��m�k�%aѐ��'�H��&��.��?��?H_�b_��mR2)h㳺 >��*�|�vu �	���.���ٳ��Oѳ}��c��Ёt�͏���˹����������̓���,�J0 ˎg᷋�Hpm�S��V���z^"�c}NaPY ���Ro�2�쥴��|L��7gm��e	������N�3��ҫ�'�;�q!��3cd�x`�mؚ��0G��=w�j(\vpKW��tq�Z�7���'���St1�N�?D�����h?N���B�n �Ui���@�yv`�IFy��K��M��[Sׁ;���[��S�g�0�a��:�tu�a��uk����@�am|]u�.^NG���ߑ�i�a������"�E�_��� �
���~:����3�i/]L݀�I�_��Ud�J"�r��=9T�հ�#E��FKw��9M���:ʍl`檅� ���JJۖ�E���**w��F��	�a�_:߆ ��=�6�ӌ��R�w}�c��?��/aI"ws�6Z�������̐�M��� �B�E؉��a��o�k����f�Mm�i˖���̐�N�������Z&X�.��_8�Χ�{Kc=�v�/9D砺��������Ν�0��D��9C=��eӪ>l���A��� @Q�e�F�W�Ef����0�']@�s�5����?gS2d,G٪��:�D�@m���e�f:Ŝ׃͈��n��w|�y!�?w1�
5z9qh/�{�]bn������j,�������R�N�G��+�>z�0Kn�jt/:EϬy���ȹ�`V	�����cyZ��A�{vo�{�RD-lQ=�e]�%��G�o��g-Gi��SqPܰ�u�s1��`�ğ���?J���[R:�
@g&���Y
�YoX��]Ձ�_��O's�q���]؍�j��}�j��>`Ɣs�ءt����qdR
��0tȹ�I����}��k yX���y�4���ER��2�iދf���R?���i0\1z��I$v��j��S�k�s�A�����O]�?�1Bi��>O����ǃ��2�,�z�K��2���ˁ������]0�z^M�l��l>ۑi�|��Me}\��Rz�a���;���H8`����O�s�&,�*�x�������}'�R.�
�@Tt�'y�÷���Y^)=��$=���a?���IL��Kq�j�#�Lr�I�֨J����k����S*as��[;r�˘{n޶3����WLp��`F��� �ݩ�s�c-���U�{��<��Kh��C	R����O �n|��ػ#H/��o��q��BuGp�L\P?�^\\r������w�1�s״��^0�'��e�x4yS_��^{챳���N,HG/��d!Ͻ���Z��X�
�g��1�����ֽe�v�T�4����?p�@���?���O�8�B�Q	�r���H�r>~��J�z�]�^���X.��#��K���lp\���G5lU�:ݫ�s#���s����g)��kCl4�_6c�T�8� �d��;��mq.��2@����f}աK�3�K3�J?�?����G���ϧY��G�7�N.���8l&򿙰�� ֩R[��Z���x�:A���ԎȾ43Ȁ����OS���ِ8�3��ͷ�m�d�%Fs��h�kA���L`��ܸ'�yoF�{���+GO��馢�S^�J�GAڇ)����[ �,�0d�8篟��;�<�|�4L�l��y�7���+����cie��L;����BiҹX�Qd[Z�wc�{ғ���K�J}�L[��L`�\8��w�a�~��{���xOt�X°T���>�x�Vr�Eϧ�Ԍ���3�,�E/�4���(/�f���~�;M�Ta�£�:����u|w�խ���v� lk��dK������Ջx�}G:t���B�*��}�tz���`�AX���C�$�y�K�t.<�,�v"l�% m�����~'�Z�jzvOKUc7���Y�Y_�V��`�D0���`W�C�Mlk���E9���##p�g9�]��`$� H��k�z١ض�������h��=�m?����i�� ��N¬��E�D������ė��>����2W<�ڮw�ܖ�$p���#��[6�m�c�{��� ��Na�͙���X�hW�Z�k6�!�igh�#���w�����;��፥��-[���z�ϥ|���sXM����0s����(�D�������x#%�ʀ�>����4��xu ��րR���8�:��Cɖ2`��J�{3������-�#<�i�L��.�G�
���r$�
 XV��2�Be>�Yz�C�j����V��ַDg�4�cԝ�u��&��+C��E&(pov��N�3S�9�zvŌB��Oǥ������M�vދ��EX�+cW�,��)����}#(�J"�zbX�^��&sa_�E�F\�|�}��5�o19f��f&8��#��y�� ���C�NkX�tn%x��h0-wj����v����.�F�����ǟ�z�C�8��ɨQ�R ׺g� �脄r�A=����sh�A���.��1��t�6�$v��=��_���v/q湾"�(���n������=��;�M��;H�������WI ��l�T��������n������7�YS�&��}��]��6�����w���-|�v5�^h-9��b�3>��ӈWֳ�P'�Y�TY�ｏ��ӓ�%��m0(�e�mG�{G��"6ꧨ��C|�m0��x�>;�=:t����Q���n�d������sk���$C:�se���G2�f�a���5M��N�d�x?Ә�w���$Y�&^��m�D`���y�$�)�]�"�&�2ՍzڝL<�Q`�Nc'm����f�8l���lʑ/<�l����1@W/�O��ގ�d���@/�K�H\~�[ �)��?���),}7gi�ݹ��Q�%W�x/�fX��<�z�O0K�޾-�^ފ��ߌ�����1Σ+���_����7����t'��1�:��$�6\������������ѣ�������?�>��� ����]=�U����_7̈́�qX��חqG���� ,q�$�Q�SW_@�>���K�qǡ��7ܞ��[�QY�,��Y �NcVg��2e �_���}��5��Jsz���v(}��gӋ�.Rf�J�d���_e����qx� �]����ݽ�C��� 0�X�t eW)�M�nAcrx+682KC����ߕ�P#W�N�V&��r�,����f�t��sہ4s3������ԍ�{��a�P=�@�fT*�Kq�ҹt �ڃՒ�T0O+�4
%̐!���|dN9�]y0;�;�!3sn�u�A�O>�4� c{��{��ձE7�����݂1��lb�J+����� ��d��I���T�\��D��s�g�y���p�Z�� m��2�쉺�>��p��a�P�L��ݣ̂�MО>J�-Tܷ9���[�gÅ�c�� ��RKġ*ݯw�F��qؑ��=���{"�:P�CJ�'�;1�Ιmk4Iȋ�,39�i�6��m�w����w4����HO=��O�}Im�S��䞝��{�Y�\���^��%J��<���F �ck��S~\w��� %Y�:j-섌��uv^Y^ҿK�-�׋��:� s� ��7�s�/�1��5@"%w2�EN
4���������C�QeRHD 2�o;� ��z�#�.,�)}��x<�>��/G���hK��V.\d��ګ��5[�ǡ�d���z��Prv�!�0�ftj�R�,]� H�g9b)�pP�(G:�,�1_�Hwt�R�}`?��mh]����
���/�S	/�w��F��EK]�����
^��Z�m�	��3�g4���e��9ˮ&�N���D)�KI��̖�����pe�dM([i|ؽ����Ӏ��)�.e]g�+|A��%��ɍvƖź�c����H�g�~*������gf&l�fF��L!���x��n��٭BF�:��:Жm�A�u�
C���= ����@ۧ:�EM��_~��;H*ٻ��_X�Δl�L�;�Ԏ��ӉҦL�(,S���{� �� ����da{��9Lf`0����Z�P��^u������0�v^���l!	ߤ�k�qmk����~�h��e�%�O?���zv����^�q�g0H#�7��H�!�Pm��v/k�$l�2#��5ک�.�鸊yc�ZJ�$p���8e���+ �=�D��}S�!�t���H�N�8�>��/�g_8�K�|��Sy��6yt���4�m�C0"�4>9L�݂/�{CG�?�]�����*�e�$�R���|���ƜM��9�=��d��>ſw�����nJ�S��3*�����L��	X{�}��:n���#����z�V�I�M�QI����z��b:�M��L���c'�J	���7����c�p���3�Y�6�g&16���a����N�KG U��\IGO�阯��`�sa����D���h:����^m����η#;ʧ�~�q�����q�8�o3����r+Fus@*��!߲P�lc��b�����ɴ�u&��-����|(�d��;���E �ͼ�C�a'}�-e�J�봽L[F�][;�XTv��lO�G>��T����G_L����"�'ǃ� �س1D��}��Z�QCF�oO��B?�F��c��2�m��S3�N�̈��c3���e���!�lD��aQ���-�d۷�������3i#u�~ʏ5�d=l.j�x1u-ڣu���@t'V��ZF�p�N͡�'�fF��]��EZ�����,�pzv�Es���4��%O(~2V�Ÿ�%:hA~�����J6e�eQŬ��Օ�q�R��p�ld��Y\�~B���O��;�c�y|j�f�L��87L�F���gP�Rog�k��ZL{7Q>��(u/�?��E�Z�Ƭ$��F񾃿=����X��6�V�d��(4|�y�Oa��xdW
�gM�mP�TO6s�ʈ�Kb�P���Ǿ��V��q[E�m]�� ")�Og>���Cϣ>%�i���A��H�m�ّv��ڬ���ƖU∝�cK�S�M6�(�����]q�v%�P�Z+tĖ�Ar.���QA�/z�N<���(mviӞ����% G�ԫ�� �l������Fr�6������3_�a*����fQ&�]�ʳ�=�!�W��Wt��p�dr�QU���f
�娆F4y��hP^B��+�� 49�K���g���RF����zX���{�.��?����O�	m�>J��B�]���x����� �a�v�ɲ�����o�9��J������!iQ�A�]g��씴3N��z&�d)�f,���OOcf����a1�|���U֎�jX����X;8��Ԉܠ�Y�m�R�L�8{k'"�]��(�E���'��
h��o�-�7^��S��0�� =�x�C�x��N����1��o<؆�� �3^ƛoFyL6�y��E�G	����fL��}0`�]h��wV�]��V�^J��x_}���$����޼F���^OB��q�����E*�Nz���	�2P2��G2T�5��I���'��;;
k�)�Z��\�¡`�&�+8��I2��)öv��st9��o�J/�$��%����� i��{������Ύ1#��MgLQ+�M�n��Dqe+c�z���i&]_@3��c
vg��:J�V��N���z��#�לo���3{�`�l�a�S�0���Nc�Y�NPK���:v�DK=cA{b�%�y�����n޺�5X$1،���9�u�s�s�ݱw�b�'��4�et��4޻Cr>��Q�$R�v�<�d��3��I7��O��w=���6�����Yi	�@�˜GU�-�y��kh�x�Th���[6S�<��`!gJ˗>}��� 
��}oz(}�>s��	]�?|�����x�B��Э{�<&e�>���̀�ﯛa����3�֜9W$��sā��-����;o�I���t���}7aħ���``�'�V�[�h�I�˰:z����N4�H��U @f����k��������H��?��t�	���c�� n��u6�#A,�0*�B�p�qJ{"�g6m�B�#*�`��i���Se��~ܨ�f�%�_�ẃ�j�o/���5X�=�Mf.BI�a��!��ŵ/�2��C�Չ��؅�S(�*iH7�8z�C�Qm�d��֓i� hל"g3E�hh�fw��.�P�꧚(l�m�3d��(�B'K�g�D-�*,]? �A���ǨU��nFL��@�S�PC�Pt�F�_n^�Gv����o˞��xm����h�`�Fq���et"�r�[Пm` ���
?��D?�F;*��?�[�ŎLK
94�@�Y�����H�g~\+]�%=����i�H0Ut\��\DXCcD�n-�|�����y����{G'T��$�=�Z�[TѸ%1;�d���tս�N�ڰS�&��@�}���(����9L�+k����r|'Y�F��#h�`˻e%e�����X+����-���!HOP���;�A�3k�}�ň�y�v��>>y�a�+$8���:)�q`�=��v��X�ljK;�wQz8����IUA���������E��2���5�5�I ��ӨJ�/[BYʓ��Lo;~"/��J0:9��\��M�F̔�'�h�v���e߮Fm9�
��u�Y�c�Y�fk<릩�� @LX����Z�lx/�B�6���~�
5��Z���9y@+ ��Ce)�4�����犲M d��a�d�e���
gr\Ot:��I��̺q��e��wvĶ��ta��$��^"��3�rB�n�5S*Ĩ9t��{���3�eX_�} C��?�	M0(��
�A� 6h��SCS��nޕ6ޯsW-�9��5��5�Z5V�ں�g��h�k�f�i���;�F���-�7�X���;6���(��֑4�)J�'޹ŵ�Y 	*0Z��ݙ�$� 0��q�QW�t� ����R�|��; ��� HZ���0ֶ�s|�J�r=�45>�Q�mf-(n�R�{ ��hAg���E@b���\4�4����y��e �NP��E�<R�5����Vt��a�gX�l��v���͸��8�����.�NJ�4���2i;{�t���!@{��82��%�Q�^�G�T�����~�8?)0d�Z��yj0�@�]�#X�T��n=�x�&�vǆM�U�Y�A#U��� �5��=[&6V�l�QO>~�4�y@�m{6������G�s����^�)���A$$��_��zH��ἷ8�`2ux�YA:;Vۖ�}o���[���ޙ��_A3�>��Ѹ�f{���z_��Msq|VVi�.�9�����A�"1�Ԑ�/Y@L�f�!Clo�c�v*�y{{��7�J�rxԲ�8����i�Z2�Z6L��Z�w�;�b����ӂ8�������  �|o�=�1�xC��^M��մt����e/�(h �x���5[��j1a���h�|IK*e�{�;���7���.MZo��tˁ���Kϧo~�3�8s9ua�I�ڂ����|�dL�_���֬B	�P��ܕ�h:O�@�n�O��.N�[Gϖ�떬.LG��j} t� =��-�)$�~��ĕ3anz�� �^O�<)S�i@�L vJ�
t��w��_v�8�Ё�jH�G�ґ��	�h(�����6�)_��4 �:�"YJ9�tF��p�F/'߃β�@m
�5�M-'���$�ALf�HP/���ax��p�V��v�Ì=V��DiS�$��-�e`m�QcEǰ��Ȫ�뢌����8���%�0�";X�%��fղ�	����o!�I�/`�\¡��M�?��,X� ��y��g8sȴ��j)H��~h�:�� H��Xg\��yuh�)���C4ls� ������8xc{�H�9(Va�,9��F&���A���e �HڸK���5�%���`}�E�Y��U�k�ky-H#�v��h��c[�RY�*���p܃קX��.-��to@�v-0��}w�I;%�I��3�����y�`�>�GaalM����`��M`=u�!Կ��	+���İ�SRsh�y�ދ��U�N9���g0�G��Ck]�Қe��B��|��d�����n��ܛN�\��f�37���QG�����7�������8���`<9~%j ��#�X��Gm�Є���ug �}8�D>B�Z&p�m�%j�3��l��<{��W �Fr�;q���IGhY��j�cd7[�5����q�2����4�9��J�M��c�݉U�eJ�% �#ut�Ws�t�& q���/$[I"&X��m�a��k�"e+���h��#�_8�;Sx�O5a��2c�$K�M��I�z�| �����}o�&��4�X0z��uH"�d"�xg28-HVIH�V�;�븍�L��'i��g/]bRȅ���|9����r��y��.z����Ѧ�:tQ-�e}�<L4d֯]
s�{J��6ޛ�ܹ>_E��F�6�X�w*I0�X��9/�E�?Y/<{�{��ڭ�N�Qk/�x�߅� ����Eمfl�f�`�!_Y�$WmZ�Y`�ϟ|%��_8K��Q�.���� H&�<��7��4�L@j/��:��#&�- h�2%cJ6}eޡ�\k+��[�t{��O��=�-��H5}�fΎZ��z�P�F��Q0�0a��l��L�3J���!��5��������?pk:�4�O�������}gH"�`�/�,j��j��p�"]T#��y��i��Cn�1�_,�V9��u��s3�ҽ�k���}K����=M D�@б�YN�C��K���B��jך�c�Xh�[�m���֑M�����ff9y2��^9ܕ�vޙj�g�%,&�[1ʡi'�A�a!�6�:�h�9h�Q&j%�t����=nڋ���7@���0��b��b�y��7!�?��2�.�fTt���έ���f�fHڼ�}}�K�3��Rhvt�ހ��Aѵ��M�>QӣX>��,�P�apagh>V q�l�B�r�8��3Z�(���ۢ-�)A��	נ�K�5j���R3�~Im����jC�*���5��p��FAmC[���e |-@;*Ʋ�4���t�� ����2op�Ԅ���O"�h�<��	��V)I[��"1��T	�ֲ#�n�gh6��v<�E�� .7��)2� ���&���ac#��)y*X-��G7.�������"ӛ�Vq۫�	���%_��3��0��@��T�Ym��A=���R
ӗ�����Y*!��ڊ�V��	�ܳM'��'�,�.kQ#�m�ʼ���$�K;k�lX�xQV�#��X׎Va�t�3OPnV3C7�l9P}�d"��&@w M�ucc�E���8 |6��j��o=��<�s���E�z�R;�P"!�lR��Rހ�V�����*�Ƌ�u�����D��5fJ�(��4X�Z�Z��&~�������7��ˠ�Üqlz�q*O�W���R�u4Gv�5���&�a��*l�:Gm]dμZ�s8�����K�L��� ��^c`��O$A���� �p*��jj�'N�hk�E��Q{Vd*R�����3��&� �9�j��א�_d�G1�QD�<����Lg(Y��yG���X�~jk��')!e���k�2�cr��-5v���,�#����=���X_���ͧ?N�4�((/"ɰ�l��dJ���-�k}�Zi8([�=� ���-�\�� ��~�iX�͑�̠9:}��:f*�w�qbU�݈�67p0k�:_B����h���w�"t��>4_�1ԩ}v ��u��߄.I}����L[.�F{(�+��l�kL/�H��h�c��!D_`�`a_���A��L���CK Y�Vާ3�Hc��aL"R��g>�roh9�`_>�Z c��C��� ��;z�1`MM�z�Ô�����o�#�^y�<���F��s��W_�������O�Oׇ�W���R����a�H�� ��0g�v~vE��Ch\�p۝�H�������=�3yj���R����H\�d�aPg����y-�t�v�E�~��C�7��~O��I�i�ef6��h������_�,���iXt�vx���Ť�8��s��e�P�_me[����;�>��7�5ے}�e�b��
�?|;�wܟ*���Z�Z�vR���_7�8;֖�K�ֵ5MP�+0���އߚ�4���G��v!������e����ОAer��S�ែ��P:q�ſ 3�����l� �|aw��ߛ�^{	B�L�ϧ�N3׌9��M[�`����@�C b�k ��HPh$s�M�R�ë�kƇ��+`������Q����	-�8O`WS���u�����/����0:v�\!��,����~�@d�����9��P1g3�B�Z���22z�`�ᨢy�d\�9�7/P�Q����lߏes(���c�*55���a� t�:���PE$:ϡ��jG�ٻ%�`��V��L�jH�4��gM9���(]YUܪ��@���i�g�L���)ˌ�K����ޕgICmXLY��Ѷc��!L}kE*�ap&�%%A��:B�a�碎N�(3 xj��򗚴������s�zT��E�|��D�J�:�ίs������};�ZGh�_Wh�\q�.�a V��K�����껍wbBVތ�<?߲��,l�I6]: ��Q�ԾA�P���ς%Y/m��1�������\���]�3�\�"�I&��][�bʘ�+';�6��l�)+��ZzF�ً�����Ͳ�4&m � ,i|�7�M��u�e�Te����v,�||�Jb����=��o���𙳄�R�$TS���D�㿬�뱖�ӯ��ih뻬Rz�f�c�k���h��ޣ�;�5�����x<���٪�)z�x��2���]���D|�i��7�-����߹�J��sW��fRes�2:"?���:��T�5m'ʬq��U�DK�A�뿘�=KV��x'��X�1�������T*OPV���h�Y_k2�فI�f6���-8���V���1��*�@�k��2�T�j�5p�I��)��
��=�P�g���`b)�������t����K0Tķ�e�L�e�߫I�2w�����8�W�������\�[��U�2F��R��M��A$��GD)/p���B6������Ala!iCq�� /�k��4��}G�
�;�BɆۙlW�	�`]Q�A�עb��3w�����q�9�r7��ivC�v6��m��bbW�V�a`/�ˎ(cGZ�Ԉ��&O'b��v�

7oܚ�h��*ցIG��C��fl#���,�����������M(�WO��3݅sAvdGă�y~��i���v�Zm�)�5��5`�_l �ma�h���ꈳ�F�Z�Q��[7�O|�[�B���i�ikHkNma�]+�V ���f��_7':˵��j�R���ܳ�{?��th7>J��yzzGy^�Vn)p�0u�m�-{Pʬᰮ�eQ�ÀLB�^m8�V�+e�UI�88<2v�j��5���H���]��/�IZ�Ֆ��A��*VZ"`�Lc��8^��َ��:�Zz��ʩmh"Xq�8*�=���SQ�������}��F�n�k�枥M����Li�"���%Z��nh#ٹ%�8X�6ن֡�`����U�� F�������D�f&d�2e��6��D�.��dx�,g00U[�(f ��h	�E�e��Ժ) ��G�(փ*@�M��U6��}94b��I۫���@���.����M?�g�����bR�?��1�
D41V��.XpX��e<S��|�YT������.��8�@!�p�W���W��m�������\dZڃį����@�|�\�|o��|�s��s�`�8���E�Wl�
 M&����=�+�<�l@�%��>V��:VȊ����
:Q;���=��~��I� (�:�;�����l>K�˰W��h�&9ҥ޲�e��vت[�e6��|b���`���.θ��c�F�H���{5����PcҰnÐ�5�Q��G`a���O�,O3�Z�{Ya��O���}>��2�9N��D�?�dN��t����\d�y�-'�K//�tKO��@~$A|o��u��֔��]����NJ@��iJk,��)���c�$�w6=�uci�w&@�\[&�c��[ p�V,��?��n��?ɔ긦����UH����#���41�RF ��#Q��HR�U������Eb�{�� ����G�4Þju�TGt.�DI3\�]ӂ~>'��wb�D3�ٮ�'�S��Y�p��Y�ϴ�܋���jĬ�Y��}w���B��~1I�$�'�Ǥ�M``��ͯ��O\�d��8���������^üV3^=�^�<Xݫ�J��u����G${>�5�8�(AF��T�`�h���!�[�F #甌��ZF�1���U�%�� �0p�)Ve@���DL�yk�SK'��gU \6t)�3��7sxvüMT�Ky_5�o��{ۨ:�N�^>����-����3�k.<�z�M8y����hN��|al��q$_h����M.#rۮ���P�*��6�U�vpo@^��%3��c�@�'OP*W�c���?�&b�D��+W�V��n��g���TjV�J�^���i�j�זVs@,�e#�A�P�S6����r�=ăM��,��ANSV(�"iJ8d�:�{��#�2�����_EDȢ�5Z��];E��Y���t�];��;��G�-���}&|�9��94<|n�.��B`�q�a+h��$m
�e4l��A�9F[qV�Ŏ��t��a�D��MM��@�KS:U+Pd�t�����r�W=Y_A����Ȓ�z�� ��$Y@���Yl,S��urL�_�WZ2vG��|6���fk=��>�,h�������9�n �D��b���h�d���n���sq�G<*��]��:$^��<<�'6�r���8�ʁ!�X�2l��쟚
IN��[�k��)R����9�9���$�H��؜���NC=�jfdr`=;��}��bv�����R����{H��p�f�Z(����y�f���C@�0���DC �߷M0�Mʼ���k�m��`x�1M�$^��(ʀ��,�M����A�(L@��o"����1E�ØL&UQ���Ahx(�r�y�Q.����Y�1I�[0�;&(��aB�C�!����ИCEf��`ȉ�����Z����S�&x^?,toW ��
���5c�9X��9�ouy2`���
]�2����W����^߭��}�M�%��YV����&/�T��������&ǫ��w�'�U\,�L���,S��2��:[T��Eַ>rv�o{CcV�L3	��R��o��n�-�@`������\W�R�#~��:�q�k�un(�XZK�ha5ת:�^a��B��k6�X�q$"$ʮG7m��5���n=�d�8֑�L�F�)���NVX�o5�>���e�!7��@#�4׃?�k�)���+,}|w�3�Y^���+U��c_Ǡj���5��̝$�A��s�R�������h�i0 ��|Xt�� .�U��̊�u���3�?�,�}�*�F��*���m�EpJ��p}��V��o���1/׽��n�4��f���<xp�`�p�߁7ᥐh�-�p����v�a�s��7��c/>��)'�,��쵡՚�+�Mw�H?���@wv>M!Ϩ�a�:ox��+���ں�bۗŖ �3�Z��M''�JZ����J���ʋoG�����2�R	�%~��, 0�81w�kC�%�
�d�ޙ�����p���G9d����A��ڬj}e�\K���}-�災�S�ưv��=���(��A����ՠq���΄Ԁ���(dv��o����49+���e[���k�P���y_S�C��L/ݞ���t/�Q�Non"�T��.$'��lf�>Wnƒ�1�.��{�g�-��4{����D�x��Kt4���bĈ���]"� �(VE:�d�ܠ��h�z�d�B���R�������ȁO��p�_��Y��r�����(F6!�2�,,�R��J����j.���sd��:�$E�
�c�� j)u�i�
,FV�S\l�#�~6��k�-���(!�
��W�� ���-K`Q29��(�%m�o8� @�O܍:7�_�sL
P��E��2(��UDXg��}���Q���@d������5q��i���f�*c���x�>n����@�C��@����FC	תh\@$��9��5/�NA��
Zp�X?\��Bw6Y"���P}o�!�e�Ӓ��J����B~�������[�T�lI����о�I��hL��JvA��w�A���Np֒eF�S6L�B��a�i���ie\�>' �c�\ϖ��#X�+�>ˤ�t��}���,����r�e��aง�a��9+ϟ5eg���
�Y`�S�P�kP���6�k�g皑Y�e����6,���z���s����%��6q��<��8�ܘ������5��"J���l�	�e͜O\�:������^����3`#k�b���y&4�L�=KVeI��)�j��,���~?!-�c.|��\!2굇�->G��u$%@	)�F>C _�� ��=�`��L����iMƿ&y��ѳ�X�W �U+C��Nt��e��>K��D��7nK䲩�o�}c�@g�߾�&dg)@��[�749���zc�`���I�����'��$ec��R�2�����4�#R�R��e�5k�pGGYg˳��٠���Wyj _U�_�T��c��r�˽e?SV&&��r)0�|��p!5��̄����v�e���������Sv�th�$Ǝ\,>�����&��(c��Py��ĺ�D������O"ۡ���\�`�,���	�?Uhh?�o���ڦ�W�u#<���|_@���_k+#kjZ/��J/��.���0�N���Z�1��.��;сw;;|���鍇w��.s�4c�PR�R����R#0x����3���o^_�]m�����shSK�����s�J,�j%ۈU��j)?�	T�h��P?S� �CW�r��ξ`J20f� ��7���2�o��ԈM�չ��E��0�o���ti���P�$��uZK��s\F�Իچ���t>y�5�rڍ�g3],k��n���6����7�����D��XD�=tוKh�X�-tz,�8�"�	�K��Ƞb`�(;("��0�\hJf,��9UԤו���5d��Q��XW��@̠�i^<t<}��ϲ�oD���c��ǥ�	�=�p���u�0\"K�}@M��:!��砡�{9C���\���ywq���	
����gf.kᳱ�@�.'p3Hs�y��z����Qm�Z@e�&����c9�C+����$��!�\Oh�d����:��\� w�U��p�@+HLU"�	��B�\w�Ό1}� m�l��.�I�ӐZfמ-��Eiݖ@�{�s�`4C�� �C?�oh�2�#˒u����R�eF�7��n�l)^�R��B�/�%QAW��4�:�OQ�D��E����9P|7���D��5����0�]�R薴���լ�*]�2+�`V\pQb�s,����k�!19q�S$��Ö���al�\ؕ�
�����Gz`)R�4�Y���,H���3RSd���09��W�4����t8 �Z��x�)Kn�DG��a�� K,e	�_g9
��r��3 ����痘͸��p����[�M��+ƑM�����p?xi�K�1�B��, @Zg�
��6m_>��l�VĤx�t)��W�{!;�wR�;D���vK�v|��������ږ�o2֗�bޏ _����9���N@At�]��aD�@�.���%l�[��Z@k��w�q}�}��x��-daEC�:��uy�v��r�A�6*F$)Y�d�{���L'�e^��Ůi߁q�Rc0Ů�Б"� ƖM���m�Im�K�D_���+�D[Ɇ�X;�y����xn4,󾔨�ڐ����Ӌ/�B�B_t�_��1���VF!�3��(��;�n�xi�UoO�$6<�z��43�>���{mI��Ob�j܁�c��61��Z����KŖ�?�7���
]�s������WM]�7]Y+MN�6����4_*-�}DyKM~�-O��Mi+�6]�����i#���Pz��f��T\�S~��k�u��A�a1�����j'��0�CM�	Z�3�>��A3Nq��6ѝ�����ŘR`����nP�ܖ��cK��ZO`3]3������(�^��@����C[  ��IDAT_fwa��D�c{s� ��҃��IˏAǒ9�c��@n
�)�8�)X�����ӎM݉F.t7W);�NsgG��uN2���hڹ�.Fc�4e�罊t�t�F���1��<����HI&�c��L̘n��຺�I�U�Y"Aï���5@Xֳl`�5��6��Ĳ 㡨�#�~�_��,Dd�<��E�K�T�����<8����1h)��Z�K@�F��qp���7J��d�tL��3�L�bʹe�"�SrQ�/�d��_�K9�-uf�'�G�ɲAC^����T�ep
�,��Ս��̀����A����f�Ϟ�~� f�P�L��*h�2n�����o�kB�b���}�DZK�����!����,@Z�p�{
+�CXa��� ��T?�]BWe�r���L�Cu}7�pw�)^#I�>B����1x����d�f�0�v�9hzU&ͬ���o�OP�8����@��.��!yp��`�U9׋��T�|� u�d���Ipxc��({��P7&�(��<�����~�Z��eK���@Gx�0B�q���OϬ��B]���)�>�L�:&����:��A��U�%MYr#.��ʁ�n��遯�,��6H�lC'���Q�a����Ĭ� ��|����癆0[׮�8�5��ή3Kb���#�
�p)����,޸�o���f��:ӫ�kT��:�#Ͻ{Śv��k�}�3enp|�����9p�߼C�����tCg�I�@#�DX׵$������4�b$Bs_,�̛��y���E��_(����U�M4c����&�gM:YRzC��1��'cA֑�f� B�T\�2��i�yb|Yfֱ�B���x��D�n]�v�;R��2�c�w����a��i�6�������t�tg�hpY#9���\b�=(P.�Wg>��O^r_����l�e��H숎j6A%�p�~��h�ـ1���#��q[���Db���5}�{ޓ0+oBo6r�(�fTr��,3ťs�H����\}��T�6�������輞�����J��ke5���F��:��`�5^&m��~�N�8u	@��o��$5��u��A�O��1L~e��A+����U�B�+��%�:lP�U�_�ڊ�!��'��3=HP��V��%>�;:$/�`C>��@��*�0 ,�g�SۮqDe�W��bg���v<��d:��o�N|h��Z�g��y|W��S��?L]��67o�Q�/N���eI�ƴ��0"R\�1����5Z�ϩMa��㕆������k���ܜ��Ps�f8;���i�<x�+H2к�Z���5�
��	0H���y�6(���!�f��c`x�����E����:�cE�����W�h��/fK��d�3���rHd�v6����Dp�>Ԝ�pƶk��\�$��i~����DV䘢�f�W~gj1��ƃ��Z#�h�U�
uC� %��L�f�T3b�?���+�~�@̲��9�{��u����SV�bp��nX/�e���
Yj-�(>+�Z�UsQ�"ߛeO�[�׺�A����)	��:FDO���|���lf��/�@�2Of7"h����p	�B�&pg��=�B�m�\f7�]$T�������?����i[��_��)sG	��ʺ
]ǚ�Z�� �6twꇲu`w����&��lW����ug�L\�%�`b2F����A[��N�,}�Ev ��r�7<�H2d:���ꚋ��=��O������d�=�e����G���3bS���\�&�Ǯ�N�Ig�2�݁�4�]���`�P��-20�1).�Ӳ���':a(��	^�^�nP��eD�kh�,ĳ��O/�"
��3]7�܌L��}���e���9fL��9t�2V�*�6��ZwH�L?�q=Y�@&��:ι��6u���k��Z�ˊ�YCH fcL�			A�I��	�BK�0l��]놐H��C�9��,����{mSdw�Hĕ�D �����|��s2`[Y��{�sL4"A�g�5�d2�uP�ܸ��}��YI���2hY��f	>t� ;��C�n��bF��]���?c��z�m, v��9����B#k��Mtn��\u;�����y^�$����HG��mM7�Ϝ��%����O|<:ͧ��i;4򕩴
�Ѓ�#Ϫx�56la�_,{����{�&���*���~em�2���~�gzk�T�%6�D�����)�yP����{s�c�J��� �8um�ϲ����Pz��M�0!TA����֮���\�67*�,�)�t
�\�[�ɧ4s���LԚ	�#۳�4К#��Ұ=A�����b�T?;�tg�H�n��J� ?N�~O���`�zvl�.�I�3�2Đ9��Z�� �_J�O#d ,(\�i���D�G�4?���1�+w����4�fz���GG.�3?��c���������:i�b�rGFwdnv��"(�ob���T����Y��'� g��'dvo֫A���X�+�!���&>/:Ђ���,p�gR_�Uf�>y�S��(���I��=]w�R�pd�� #�t#��x=h(B/H0\"���:㥯x=`ɐ�.����`��w�U<;߫�u�;�Uy
�����O�+e�]W�Yp��8�0&� nr�KY��~2��e���z9��`o[��" 9�u�[43u�^�Q(�ZwX�)/e]�Q������vͦ��e�j�н&��
,cP�7�ՃK6a3T�:���]�������b	K͖"�u���%S���G
�S�V����9��,)
x��D�U~7X�l��=����TOF�JC��{�2	��De�O ���F �x���Q���Ưu��{�9��o��J<�����dk<F��ɒ�fK�62P�o�yj֌Kރ���`�,mʈ�?;������bw�@������l�� �K1ן#�w����F�VB�����@�#X�`�łDWq�>3�0��7�D� )XŨ�/2��mtS�5���rm�i�� 3>�}Ŀg��Y|ɞ}�b��ǳ���3F:P�z�D�(�&��_4k>SJ����=���H�Ze��S1k���M�g�c����cƎ ;�ZA�{���3N�8���Rjց��n��>#�� �jcK���|�yd���c�
FՅ�ub��#[�QՑ]��j+�����~\3�rf��.ٸu���8��?W �;��2%�{����4>w	O��d������i����q�=��|_z���ҭ��¸�k�,����f��kd��M鎻������{s��Ï��I���4�w�^�^�R�gZ��̊B����\]�s���
i"����_5�������\����Z�],=ʒb��r$�u���TOy�|_89��!L�\D�G�����k���]7��9�
���z|;7��Ԁ���P���#��!�
6�uin��S�>���B�ɫ���0����3a>�n>m��m5U�����'��ᬵ��,B_���5��M0�kEt?�v�y�i��<AM}`�TfQ��~%�_KE؈�6���/��������Υ��C��4�'�`9�)�S�`�p���ȸǭ�#
݉aQ�2�sc$�"��s2��9x(|V�a�Y��g���1hF�%t7O��$+����`��n<��7��+�β����lQ�BYhp�,���gU8�3=�
.ۙ���o6j��?����8���(a\2g���e&lT����<;3�/K8 	��L�u�)�4 �D��о��$���J8d�X ͯ�v齦7��f��F�\u$� ��xЅ^���%�pqY"Y2��!x�`����=�JY����,�/�N�E3\���`|׍}#c���pT(���ħp��g
C�uv�)����2j��(�e+�)�e0Dg�^�ߘv�n�{�D&h��4;v�`t��Z���Ĺ��׭��s=áQw���i���]/��"����j	�j�,=�ֲ�&�����2�熭JX*8V�p��X���"��/���
�P֕Z�1[�QTmrx��"��`*����C\����+��7e��Y~Y�H�,�t����LG���ugfI��E���-��1ϥ�ΎGgv:P�����ޣD %ۃ���A�k&t�QB��*�Q��<�W͵��b��c|��l�<�<|��D��(g�Yt*F��=��^��e�f�1��}D�Dh�2��8�)�^��*��Y�F֤QBx6&DZIx��X$�����S��솊��˴q����ך�0����Ǻ���we]�[�F?_+T2��3e�g��M� ��qY�M����?�=�i�n����`G�?����(�*O0����n�������`w����Zv�7�}R�aԭ_|��������]�������d�U�hh���C0>�ٱK�֏}�#�#��>~�w�:ͭ}���Լp=}���#��rh��q�/L1	�����}5�Z_�<�+�O��ӹBG�0�'��&kj���j��䪕m��j���j���I 2��:��۶ޒ�0ct�2��vzp v�����[�m7Ru8�5�귱�76�XsF��Yg��
,h��#(=�c����(�U3�=�j<�_M���50^mat�2�kU̩=��NJ^����� h�_�T�w�SF|����c}��/\M�;�;����O��N��c�����`�v���16�u��.Ӂr}��<��of��ƚ+́l��ʠ+RkOOZ�6��B4ٽ5n��x#1AYP� �4�Q9���=��g@QHm�d��{@F�7�8��Ӳ�u����S� #{��!����[��lC��_c9��A�|΢/�ϵDf6��W9�.!~��,��gqmjwx���c�U�,c-d+2�?{�c�9������S�a�F���#�z���k#��p٭�s�,��#���NY	���'{�;�e%��T���Ŗr˖"*Z�X���=�4���4���>-����=$���K��#�u"ˎ�eY>K��X�2l��$%T d�ݿ�0�Z��s2�{��eg4bW�Jv+0���Ě��F�ϝ���U�� �\ J�>+�8�<첲`� ,J1���D3����e0�V�1�o��	�t #��@T���o�J�*�{��T\et�2�Ig#Z���3�7�`ߞ�����M��?�	F[�O#�B���(��v_z��A��B'X ���L$'bI0j"��.y���Rl���U�����Iٻ��МU�V�#Y�}u��s��~���Q:��� �F�� ��=���s2�Jd4�$-��X�2o��bƒE}��F�%���葱���랊x�i�BCi��OZ�"�0%����ʸ`(0(bY0�Y�$�y�Q�C�qj<���"c��ōi^K���/��:�}�Y�F2�O��dͲ��ɔ��L�LFc�7�䕡^p�;�^+[!3�މ��F�6K �8���gR���b��)&�Y�W�>����\�g��uTZaV/l҈��x}2�T`�HnC�i�fm��q(ʚWg1��dc�&�*[~��~��y=X5-��>�`����?���3�����P#P.2a���1Q^CG��p��E�W~�7��#O�7ޜv����O�xg�f������|Y� ��
�o�W�XS^[�����DZm���4�l��w�D��g�N���M�Ӗ�\:qvr5�؊ZA�M������� �Uc�kmh�u�$Uײ��R+Io��}�ǘ�{��e~�#u�^p;�=���Kl�W�:;�_:�ȚS�!dd|?,�����"��wT����b��r��G���87�\� 0�ϧ��R;�#�wЩҞF���s#�
>O-�=�V�])����Z6�z{2G����4?��a+N���i&��7�I9�o�,�Zx�ȘȲx��%�8����8��O6��3ȱ"�zP[ &;��D9��Ʈf�
g2�a=ρ� ���2G���Ѡ��=��»G@%gc6Ĭ�\�AH��F��~Rd�v�Y��̰n�F�<C5���7{c��6�3 �� ��U@�ƌ�l3;\|Ǟ4e~�",kXX�
m�xPBb`��#����Ov�ɹ7��g�}.aÑ�(_.}ޖ�j��݅g��_<3��H����
�Y%���S�^� �G?��r3�x�EiӛR��4��Уi���F2IBwO'���1�8���A_o,���\8���gmD�����9����2fނ=��d-���U�e	qU�7ؿ��d�Y[�e��(�X~�.���s	���%`ɦ@8�2��(A��ۄ�>@��\@���� �n؆�膫�޹���л���5����d~p
���R �u�� ��楞���\>k�ȹ?H�L\b�o( S�=bl���}e��ctLA�	z�����P�r��X�t��$<��e[gA�	.����4��1+N����ԛ�����F1ͬ3:��HceN�? ��JdmHt���CjG����#��?���=����`ia�Y�&��`�x>/��{�Ͻ��f$F�!,�/.�)�K��z=&z��Z]7���9���!�V���žd+ �kW�}���8��u�uW�۱N!���`(+�����������s�d�G�"�7�ZN���lv�f�L��B��lȈ�&B�rU8�+�"�#)���9��j
T�C�'WǬ�)`Ǆ��;4�^L/CC��y�-X+M���~i�P�S׽�U���6��CDБUjZ���? �,D�����<2�v�b��i�d�5!*�X�L2���a-��WؓQ��.���m:�l}s����(I��+C� ̧�B���۴��,��ݘ���n��`lns<�6H5.���f��$���;�m�gqf������H3��'y�#,��BD7��=w���-���e��!�-�$�FUDk7;��dkl�E�m�ܙ�߶+��L�RS!��R���5�U���\?�˶��z�D�-�2�ds��4Q�	����^כ�����E���&G��R+�N7�$�d1�FA���L nGA ��rf�~=��;�%!��:sљ�3�	�3��1�4����K�W��5\��۪��A�E��zI#�s��� ҫ31���<�3Y��l�>9 (D�S��4#����@I�#%���sШ	�eZ���қ�_� ���u����>3=��-,,DwOox���7+N��+�փr�Ad������LL�#����2�#FI��pX h��Bqp	�a,�hPk��,�D@��{��R.�m�s��B�#{c�;ׅ�Z������X1D��3?��	��1��"P?��,�l���JnYiPM�@o,Σ��J�䦬�����N7Y
�;D�qvY^���z�{�h׿��wZA� �R���73_g��́�^����%�%)�9���D2�
�����-!P��Ȫ�YD�\�Se'����f�j�쪣��L3M���3����z)*�֢�RИ�#�:o?4��g�1%\ .\t�" (���S�'�	�S�۠��C:J�|W2Mj�2�I����e[;W�����\��J9.�,�7���n�x/��aכ�Z���;[���Q�|XO��Ygi�L Cb c�.����p��ʮ��^�������\�0���MK���͚�RY������d��+�yk��O�l��et�Ee[�a	򣔙5dn��Q��nb<�X��,�u��0Fɖ{X�Hd��:�ܻ&�.wc[`n=�r�½_��?Z�d������Sc�^tO{��+o8+cZ�t]ús��6�ho0�!1�i�~�*XMPC%Y��X'>�cfNl�� #ŉX�/��s��]n��(4ذ���@_���x���m��M�J}��/��λ5�x��t��U���ӏ���ӝw܊y�%y���s�4$��O���j �fuvv�®��(�A-�q���q�zk�k5E@S���=�������e�+�#<$�*K���+0��Q.���Y���ikVOu�F�Z�&�[��&��R�+Wyg���� ѶRn���ɢ�AQ�/}��/
�,k�Ȕ	|��B��;R��������u_���Ά�MG��Y�՘�:�%�}���{n���q��N�<����
�k� e7Ė軮�#�JY�]��k�5��B�!�c�4L�q�2K'��[�`��di�E~�Ȧk�l4��u&�s.!ya�(�P^������n��`�s�l�c�]�TDʁ����F���o�}��(uݘ��80� 5��m��[��U|�qg�Ҏb��ϲ�)C��d�u5�u��;������>p���+�#���5cR��y�M00�fy�� �2c�~M<���t���Ҧ���{1�����0a�i)��'!��Y���L�S	�x>\�m�m��e� "����p����>��댠g�߮=�4�� �	mٶ�[�p�q$��[d����%4�st&�5�o� ˋ�%����?:L{1$��[<m��k#ip�vv�)�5<��������� �â�y����a�47����ݵkWz���y�H�z�j�����䕁+��p����,�@�|�{����nY+��mGً������ը�@��k�Rec�ZN�P˲:����j�V/�?�q�����z�]\�8H����v^j���α$*C +�%�4`��I�֎f�Z~f'f��9� ��j���+[dL2�c���`�pc�Rgv�Ɓ��}���K?�J�Bו���D��0���-7U�#���l&�i="��6����ؖU �tEI�2��B]QfΜ1���3:v�!�s7�ژ18�g����;,�L,�s���nO�������32��2��Y���WZ�L���)���<�l��1.J������*lo���o�ª!i���b.���:e�-�
��\�mᗕ�=��S�fBa"���lH_�ܟ�\�l�'�lDSA���w���QUO������!�|��)Sc��ٓ��ɜxV3|O�Ip����N��i%����u�Mܯ�i�R$�쿫�Cahb�x�Z�.�eF��h�^��mbz�<+�+�x�9V>q�� �N Y�@�xIg� �q��;`�7o�����se��s[L[c���w�
5�w�q[:�� ���X�siﮝ�����=��}�8�i9�S�l���Ao����<w���2Xaޫ�G��Vr D��M�*�d��xZ��2�* ��� �2��J #�f~CO��n���m���auǸR{�cj�p�2�rd(t֖�Qc�����\������j��%�+�Q������6�׶Q������
�f�HpE����>;k-D���	�K3�8M����Sc��5 .\�u��7 ���[����l���+�im�n��kz�R��I���2pS
cSŊ=tRr�ϳ��Gp"M@'Z}�Ǯ�;�mLvn�+�1J�K(۶n����C�}K/�  V��t���#�6�BloiĒ��Z5��Б::iB�>�z�	س����D���a�/�~��������(U����調�S���e��8��6���̀��-=����ynE��660!� $�8�Gy�w�DY��4x]&���)��(��4S���0�:��Ȇ��������<�.1м��v��u���4$ρ��gֱ��A�;��NVų7l x��Όe�x��49����଎�~j[ �k�^�k�1@nh��G�|���d��������t�����`ڵcbwz�WҨ@k���?�Հp��a�>'E�3hwdv����03�A�)�u��������}iׁ�i��p:��+a��� ��弞�4K�[-q�7^4�X��4������iؐ߶;ؽ1Ŕ����Q�6�J׆ǳ���G�8*��yeq�\צMQ.ͺذd�>n;t�d �g��:<2�0�4<>�/�s%��U$7���k��n�@]�:sD� �܄���9�&�5,� ��`���<�?e�Y��c��IS��yL�e�Ӗ� ��N;v�N�vn�R����}˶��y��ұע4�1b2`|��sG.�yh#d B�$�y���ߗ������<�ҳ�փ;�8]��._�̲�
����ge��`�$>7}�l�b����P
M!���fe���t�gJ0q�B��ܪ���C˩������"���\D��7ݟn9���eIR�-��Mi�
	�e?5Lؕ֣!�DM�<~�#h_b/�E}����G�	��/8�	u��}��"��aЂ#��55M|jx����4�브V���%�}�mi떍�٧�N��_H��q0�����\@�SΒ)�s�P )��Q����D���OoA] >�݉�hg:|`O�v�"���zz;�}%�Pzsh����aQ��<g�v�����%���|9m��N{�������B�e��1��dk��!�j�v���.�1qo���ͅɐ]��/F2�8�gϮ���D��KϦ��=Q_d�[�l��*{h&���ٙ��Y7���1,�\gCm%I��|Y#��ϼJ��CK���,��.�n�F!>�@ե��|� B
�inb���Ժi1 �4���K��[Y�NN����O���D�M��Z�lʜ%fC^Je|�����=�A'�]�h� ���:t�5$h��ef�љ�
�'��_�f���Ԕ��
�B�A��Q"+�l�3�aO�8؞8�R� �m��8( �����_��n�I�3U�&f�������R;��s��P+2�umX|���ߡD��(��$cus��-�ƌ+a�K�د5=�2��MAj]�jo�����x�fIE�Mw������)q@�2������7o��O\]t�v��C�HvrGjr�w�p)27�T��vD�Ԭ�7�v�C���|��8��̩��+G^JO|�`�J,���.6>Ul����^v���mؼ�03%l5��·�G��;6�\�Al4��g�-�P6|-s5R:��a��F�c���U&�7f�:u/����;���� ��j:v�xz�c���%�+�]�X�ب��R�v��:��#Tx�
�72���x[:pp?���̳Ϥ_z	껛{$��ܴycڇ�����t�܅���5PʾHPo$��D���!{��0����i�-Q�!8�684�5e��R����1�h��K��đ*z��a)x��mC��7�'���d�PCW\<w
�n[����!���3"y���zOz�	�����a9�����[���a��t��#���$�r�Y�	K���[�N-�V2w�ܸz˘u^;?g;vw�yk�V%�AM�������@�����_ϹyN&p�*_��L��GE֩#Q,�߻3=�� �t�{���ܺ��uL�`��r`��%�X�*׹$ c�6r�����c'�|�z`�.֡�y@`�.��KW ��ρ\��²���!��NvW���mGGK:t����e��'���m|n�>ku���A���N.�od�L�`�d����uKڳg7��a� �V �f����l�(]89�1��4j㡹�ل�� �{�{jb�T ZX�M�ˁ���L�gϞOC0^�lZtQ�}	,�v X5t��ɰY��gi9�Hhjf_�,vw���ҕ�#|�te���-<_݋��}:QfIϭ9�U7	����}{7��˩���]�=�������~#=�ܑ���oG���j��JǷ��L41�z�׺)��}�]Xt��Z;�&���I�b��/ʮd���pԏR�Z7�R�5{�Zd�(^�%!kc��+G^$1&�8�{?�y��F�T$Xc��4<�,e�4��d��<�i��v�J7l��ŋ/��0�o&��,���_��7�cO>�Rc�
 ��ÿ�F�t��r�\/��C��[��G�+�O��|��?L�����'�������Ͼ�s�i��ii��g���(� e�Bz��\��x����;Hlܺe��h'x����k�=˨�,�:�šAb,]�]]Mi ������IS�F��?c���=�I�4s?�d;w�Lh�jH�L
�a�KhJ�
�ƹ�u�?1s=���@�D�8��5�F���#��;*fU�D�f)��!tkK1U�s�~Ű�o�3Zn��,�)����C(�	h��o�B��}�M�0x0�Vkuf:_]Z�O�t/U��n-^�XA�B�3��V��e3J3j2���8�����*���L5�ZF�A�X����"�������ϒ������������yTt+�9�m�"W�fq�08yb�?m�[ϵ�e�̯
��
�YY�:4Y<� ��᠑kië�H���1;
]����?.��<�H��NSW5ru|�%�9LYG��\P�e Q���[S��^��v��TE�
�:׮ӑI��Q3�և[?D���l�`:x�v�5�E�u۶�i�.6�\:�A}���#��IX�L���%2�VHA���,�y(xp��N�g�عj�޴a׎T"0����HO>�lںcgذ1�<u�D�6x5D��(�m#T{��]0�k� �n��nI��~�����kW))�LC ���� ��������Zb�~�w��ճ���}lH>�`ڷ�v恎�{2��\��{9 ZS@��lv���ޠ�A2�X,˩�d�Zi�Do���t߈�t[�<ڶ�/|�굘/�H ,`s���4�v��&d���=�%:�A������������l|�_���<e�YZ�s|^��_�������%:xW�B�L����ؿ�΃���nK�t0������L���i�X���\Z&��hDd	��dY���^ذm\���t���t���X��̸��U��샚6��2}3�_��753le[w��֌9�5��Sϥ��-�	�"ˑ�E�l��{=�y�D�.@c3����}=m0M{ӽo�?�~��<7XX��)��r�A��0�U����y	f�O��\�Wa�1�
��ϡ��#����sg��J:�����+��ZGK��p��L����,��S����{��m��� 3}�4�ΝL�����3Qm ��Ye-���T
e�ڮxpY�
��߱�����n ���= P���}b�Z^T�-G��|���d�����=�-:O81q*إÇ��|�G�b��?gb�3i���yk&Z�b~c� %�&�g؏�	t��I�����'>�abUg:y�l�I��1l$��>���i/by�	svK۬��	�c�D���u�B�n�����5����{�(�+<"�D,���z(�@�p�;��v�򾆮�׎�]`g0��i��6��U���.���/cL�d���O�=\��f���Yd���^@���R۾�ӛz#:�&ʻ˔޻��}:�
=�g���3�>t[]HB�a�GI��z �	�	�?���f��d��x��A�W+����@��5����tkMB��z���gM�Lҝg\����ĦɄ�gRO������M��݉�T.�96�kV���������I���-�:��9��7Rś����p� ̗�
A��ظ:5���7X��҅�^Ss3�<录
��f�veyPf�ʃG���pn��~�i(T@V�Ǐ�?�R�7O0uNv��LQF�ڻٷ�����|�J:uv(]Z�IS�PX���3�*V�V��TK6c[ t��RVO�Z�J�������T����E�DI��B���S���͕,�?�\a�d4�F.��P SEa��E������]��B���#�>f��<@a#���L�чk���S�m-N��M-��罡Gj 8:>����Zd����c���:��>`�֖4u�[|֙��9�)�.t��
�<��_��y�[A��&��fc\Kf�O�J�QEז�yJCP����:�n�v�w���@<<`��0ja�^�Wߟ�If��]�Q��, ���K�@�^\|��D���j���+�AZϟ���������s;�� �KSuM�0�����ԚF����z3�L�㲏��֑<�B��% @����E���gi��V7omMG)ɍM<M�M�GI���}���y���m���y�R� /8PZ1n<�(�wQ����K�d�Q~(���ݫ�������,wl���?�#֭g���/Ƣ�QF0a�~�3c ��ﬃ0�C5F��(Õ�h���)~����NBԂ&�ϙ�8ٯ3
��5\��̡as��'� 1:FYO�\�#jd�:;��\Q֤lg��ٿ��h�g�d3�h�a�d�ֳ1L�v�\+��z[ڽsOH!Z�9\�xv�(�@��#o��̚_�0���w憚H�M�:8d[I����G��[����Bo=�Z۝�IR�H�2ecYn��
���|��"���Q�<��{���C��;�J} �C<;��lF�X�m���c��e���/�N7Ǥ�rڻwoz��o����[��v �I���Z�M�/�A�g��@J|1"���� ��@:x��4��wt+�����fHZ�)Uܾ�G䟖���S�{I�	l�S=H3�����u��ZV�6nI[��H��]� :�������u�;*\OD]�cb��X�;��������#>��rg�P�k<M��3�V�u4i�X��\oÜ��VAo+f�\�E�f��@__h�&F���%��51;3�.���foo�CW�v*�{`�w��SGYM��mL p��c�՞4hn��;?ϦJ]����b�,�A$�
�f��	%<x������5&Ԭ���$��k�^�ق01$-���&Lm�%h-}d���E�����Z]
r`��*�&���_�~� ,���N�쬎�UҎv�H�;�M{�Pp p�To�`�0J	��It�(�_gd���7��ڂ]��=A�g9�ǩ)k��2I�M"C�(Y�A��e�:�-�)������qc�Y$��_���{<��Bk>�V~���w1PHm�f�q�[^��_�75{�ˈ!��� h�
:7#�ܼy[:}�L�5�	Jm�*�S&�rg�Ri: ���%4��P��!��9
�in"� ;vlI��J.X���������ճ�9��s4o��9�ib����}��k�P�]�t��x&c;9ݱ
�g!f��1Ӏ,57fpm4 ��޴���ڽ�Lt�C�Z0h[6o�j�DY���*(��h�Q"l�V$���/��͛��M׆	�M�l�v�\Ϛ�d��e@�V��>�N�#�-���B��t�K��%$01���p�Q����W<,�b�l'V�TM���.O��A
|v'���Փ���'
[
��7�÷^o!���@�W����	Pv����K��a���6oݖ���t�ҕХ�꿦��/����ek��E�C��:<S��f���=�)�J� M�t	��Y��:8���Q&����%��]'ܷ -�TbĒ�GF��{���p;�|�Duz��2%m׬������6`��Y�Y@u��=�-��z��e�s���+(n"����eE<�]�:���.���W k���~A�4�	����*Ò7� ���hA`G'�z��nF���6t�ܳ�:�[	� m-�_�h�KS+@�Ɯ6V�<`�I�
�vș�ɢd��l95�$X3�ܼuO��������j���w��seA�Cս�F;�V�� ٌ�ք�.W0��nmS2�O�]�i�L>b���r#�5!Ղ�g��\��5���A:K� 2::c�� jm�����9׺����f�V�ď�{�����X���EX�^�NGG����1���}�{��n�U��K�윞�FCq�"��	Jb�mH6l�N���H�C �5A#F$FL��G�M��!��!����������Zﭺu�%��yn1���P�<r��]}���}��9��������oFP��.,oC��s��$��Dx�M6M�(���i¾��H�qf��p��k�u)�;���17O�T�¾�f���(�3��
F�x���`X vB)P�'Pw���!����h0�#U��e�`���0ױ'�&(�Q�>�q����D��V:��?DPi���~-�{�F�5ʬ���ގ�l�&�fK����g��jL0��ƚP��I�"�d`]c	<��v�k��N9�=s��q�՟@\���@�mFԦKL�q�7�.z��(�KL$��h_Xw�����j�.Tޙ��9���ӑ��0�ҴC������DrLń���Gat�"^_1*��� }2-�-�tKF�2�};�h��tNF�)��4��X�h��BҟH ,y4Sb���c�
D�e�V�x44"k����;����9H�:�$p�th��4��b&g���I��FBF�1��q�QKyG\���X��d�8�t �I>T)�!bs���F>���g�ɣ�� �~sz�<H-�Џ1���Ԕ�m��Qj��(:/G2��}H�}��-���m\3L��9����d�A|?�P��"�E��Eu2s�L��)�jc��8��7�iy~ ��Ѫsp�~p="�E�SC/�@~� Ak�e'���Þ��1��+oG.s��������)��+�YҬ��)$��8���-�+�F�� 5�v��gDM"�`Q�R�1��LW� �r��ެ����T��.2s) K3O��C�D!ZQ�L��s��8g
�JzJ�;�	���5f�a8,͓���<��t��2�����ej �uu�H�i�0��џ��J�i�:�b9�l����3��
�ݻ�����F�,"�o���M��W9_ftZ���s���٘,�pK�XΝ�R��:O�c�<`ٵup6�ãh���n0�S����r��-�+���w�	�M|yRu�ȱN�Ѥ��.��Υ�{��,)#���h,��p|������Q0 ����d��D\�{�2�eq�o1&��`�r=�_$+ky��y��JZ�9��$��h3�2�<{P�&g�l��U�s�q�ګ�5�3)b7�|��g���&HH7�$���`��Jh�8��!��+`�I;"��D_�6(��Ҥ��W���Fcq�� |�Y�6���r�sMf|�r�mg�"�%7o�g=����	L����G�!�q*��ZF�ǌ'�miJ;�,Mm�es˟��d�y�R.@�y�&����-��� �+����{�@caa�{�g۔��<�%�����nG�������E�:_N��.%�[�vl�R6�R?{��c4̐9$d��q<��ܷ��g�Q{��kA|~�)M�?R�B?1�4���V?��e�@��'�����Yړ8ϙr��߂K�t�LP6�k�@qEg,]�pG��:ΤY6l�"e��\*.f��3�,�}{��tBe�g���Jv���-h����s�;�S�$��C:��9&s���Y0��n���+g���g6��_^��ݷك{��#2k�i{�����+Ο1�
 �:`�nOΈF�~��\���x���-ޙn�����p87�6s�.d�#�"��o�d�Y�e�yf6s�����
��HU*������ L_0)�����x���1F����3Jn�Γ6W�%C�}�|��aj�Zg�fT��:��`� �L�!	�BJLKo�8�b��m���)p�[c�qN�����1�y"�5	�d��pH��""'�6���le�h���a,A,Q!5`�XN�>���]Q�k��N�
�pf�����ײ׿����a�Z �X�;$3�V�� ���9Xm2�-"7�&�U�߁+��7�f���,/���ۨ/�u���Dz����;�N�G1���U�L�7�.�5U'F@�*OW�~�T��(�i�4��2t�tڹ�O�7�����/�!2ۥ2���1�t�,�7����ƭ[d��#����
g]U+(�5I��)�����&��&��kS�I��2$�����+ٕ�7�>-�YEB�k]U}n94�߸�{��m�I����f #�hQ������_�NK#�P�ƀ��.y���'���k8T�{��Rr�v�4�;�-27��������x���>@*�(�C�Eyy�.S�U�n�l�G~b������]��k4��?�9%�v�n�]����A���J����|=?�bP4�]�k��A݊�ٲt�q�6����e�� P��i���tjUU��!�l�a-��/L�b�kz�U��� �S�y{P���9["�T��� � պ6x)j�ٚ�9x+�y�L�Y�e��8��wފ�?�h{��Hg3���L��'�N�����$V�i8}�U�'��o�y��1�a�G�ڦ���jن��M;L�yx�2�� �?�8,��w �.n ��o��un�gz�����#h�� T�y��2����$�K[0<��U������+���~P#��$��;�]%�8d�i'�/v�h��yK-h�֟x�r����������]�Y��B�^���A}5��sS��,�Du#<j�����DY�k;�t��i� n��.�q3['ӫ�ě��Y�2{��Zǜ	��̩�ĳm0����OLQP�e�&��*�4R6,�~����@���]�����L���	�as �%2����؊��e��� ̵�~�v�h+���V�"2������6�p��ۜ����Q���� �޽z-�
KR���.��\�`��(��s�iӑ�Y��EY߿�a���U���Ҡdy|�"%E|�6���]�PZ8䖙���Y�	�F��#��_��W���Y?�`�>��Ogt=ۧ��>��1�xi����� �o�ޯ�������Jv�{�<�������'X[ix���	�"tK��¤8������`�~����}}��I�/e��	6>?!q���:o��Q�VY�8�wH�T�֦t��Es�����#�0�[����V<<:�_����A��e�@dW���C����]X�=�#8I5��ԬC"�������NK�
5ne.��U5P�K��~H���
ʁM2�k��Y᧑N~�����L|�Z�FWF�F�1�4:ΰ���H�,��@g)'B��3�v��|��F��'!���=���L�i�o_	��F�_g���N�}-��L���!\�5�����������B2:]����ɵْga�7�v��)Fi��MJfvg�晴F��1���F	Er�:`C� 1V���u�Z� ��c&q�	X l$���yH��)7�|T0��ev�x}� #ju�4�sD�q�O:B�.�3��=Yf\Z!��,���󯏁{���ϲv�K�`pr �������`6U�*�R����G�A�Pp���غ}/��D;�t��c1b$V&�:Z�8fTP3�:}� VU����ZD�f&v᳙A9��%�d@e��@�Gd�$OM�J�WW��td������,���(�&�f���|>��9O�6����	���_`z�S��3�E���H�k��pl���Uзb�y.���.8�)S˽�Y||�C� PpI�je,�;��by�ϼq�^D�]�2C���4�U��Ҙ�2��sH�F�fq&���N����q,i"`�
N�̃]���1����$�mu ���H�L���Zvr�y]d�8W%y3(�ܺq;�/Wp��8���:�^�E��v'+#`�GqNנϵ=z�Cyw	�٤4��ڂ�t��]��q��o��6�Ĝ@l���5SS�� 3�v��P�Z0���z�ý
N�ه�o�|����r�8�r������9�0'</�gf��,^�|�G��n�. A���4��~p�\KKif �w��
����(��	f�fn�>>�v� ���C�S@��"�@vƠ��
�"��s�soi�L�A�`��fw��@.�sݿʶ�'�p�� ��� ��n�?�U:[j�����y��kA�ei\~������^���Qb���Tk,�N/a��K�nZW\�s��'�Q��?�۝��aK�r��>4K+ph,h?R����`0�*�e���Uli��6Z]��؟��nd�4Qu�tl��B���8@���[� 0ʰj�P�̌��G�;�m��޹���Ag�5@� ��2��٦�������a��������N����g�H��d����d���`�/���G�����b�.N�_�k8��xԠa�������	�F̍�Z5P��2{y>k!5B���>�裣la�s��4K��6D�����#������.Lu���s87�H�X�D��v6g�]q=��;lZ�����FJ�R�\U����9��9�,;�3�Tp]��Ne�F	`�{Zn����C�_\*{�M���P��q8bCr�H���-g@�!;3YEj�Һ�gJp-���pF�n ��&iL�f��J�%��IL�8�D�KDS���U�Cp`�dL��s���#q]WB�<<0!�⼊�r��̂4��T���uR��*D�u�NY���@�0����@�z8?�atIl�����LT&2��9�Cf�	���ܘ���;�&�����*��@�Jߏ�^Aˎ�H�\�#Nx?�Q#��S�2DV�� tZR�� v^C�5H�C9:d-���׮oo��ݜb�4F���z�;mJ~�t�Ƀ�x/�c�l���@�x@�~�O��6帇8���^%�F�����|8�0�:��q�y�\�*�� �;d;��~�	d�莵$i��@��F%�%�3(h��ا�`���Y���r^�\;��7u���>���{t�Ή���{�g�r�7�B���呜B�Ȟ�����7�cd��t��Y=�_r�tT�S����Y�.� / ��F)E��6ch,i)jk�.a��f� �o�yF�y �Rdt����N�����\#<!@lQ[�k��ε)k`�c`��e=@7\��(�:򺸧����T� �8͘H�Wt�@��2����}2wR,��s͒)%r3��!\���-C�l��.���,p���4�S;pDv�쿥c��ef�tKv���~�Y\�[��(rd�<:\���VO����ђ�J��ׯCF����HX���)LK�*�3ن*�U��r�M!6���~Hw��o��̤�Q����F������v���zD�)���\�X�L��r�Y�P�+g_�3Ȗ�|](�ۄ#�
���J��s}U�O�W�2m[�õ|/��{�C��i �W�U�cK8%��3����
ϭL��D��iСP*{����=���QWrY
�,5nf��f��D9��g�}.7|dl�q�g��\���v}" s� !Odqz�2�g~g�6���)�aQ��ɗ5�R�B�^/��M��OHB�B))L����K����y��yt�-����)jevy}0,E���nf����͂���_���Gǰ��h�h�ڟY~��=>�6i��W�<͍�KNs<�a��67f�����P,�_�_�Y�Y:>��F���4{�*�A��cp��Qw��dyJP�q��� Lc4.�{�򔀶2����?����<~�
��@��e�o��b�X�ݲ���P���J�����s�9H��1����.#�0@�F��-c�c��1)��f���^ͮnQ�� y8�"$�F|L&�+�P������}�q�\O#FB#��&�lj�w���c��cʈaY�������8�C�I-���Jy�y�R��!��=2)�$� ��a�<x)��h�4%���O'�]TD��d�#�l�7��tZk��)h�.���u�Es��C�)*��3��#Ca��0�g���X��1�['�"b38���N��]� �"ѣ5�l�6����\�a�Q#�5��vڙ08����D��#�p����L8��X�k��:H�/8�,v�*�@�gi�$�ЭARД��ʥ���}Y��+(;i�E�ဨTf6�Ϻ���r�?N ;���	;1�\W �=Ui�k�疈��o�H�״r$Ͷh��p
 �528tG�f/o�>#��;�C
�lƊOŬ
�c�o�̌���r�}�v��XBT�i�� Et��\	tʹ�{����ڎ_�UB�\�� U�h2�*q��T;�^U���T��	�-u:m�F�F۩��?f
���<�ݲ|d�9c��.���<j4�y�.8?3�ip7B�����1�eך��,�".eSBtS�]'~Lf�J�q��HO6�lA��	Ϣ
X�	��,%��͖{�#nP�U���� s��@kG��2�U�@�F�8���9K6�,#���a�T�f3J���U�A�٥�Ըf�f��: p2v������;�W���u�>#����>�q�}k3���є�O��4�(��W��wl���t��r�a��W�9.��{6*I|�r�O�G��[z���{9�<W��f���`'\���<�1�'�-y�f�GRXG?Wa׭�)�=J��yG,q����ڣ.�.#h-Iv����
��p
�����G
b2G��1!ӞFё�^7#����ڬ���:g-Ov���:LR��!�L��{f��l%'����A�Fα�R3�mޟ���h���Y���S���v�Q~�Wv�$�>*�R����i,��03�vwï+�l�0�;�9��\�&ze6�~���"��3�5z��Eyv�̹��v3��׮d��s��~Lt�.vWH]���Rr�R���}ne�YX��{���v.���Y!�NzE(�Mu7��珏�� ��t��I�y�܇�m�~aK���ۘ3}�z;�#���M�v�����țTF��Y���6�eG��\�ٙdo�mRYʞ�?F3�!"k��ė Sǐ�0d@(Gز�<.%�,�xx|��HP ؚ0MޖV���#5��Hk���ϖ#;�a��Ⱦ�[�lg����,b�
�C�(#��UN�~H^��i�X���,r��#3�D�8+�E�{����S�y�S���z��Q�S���[3:��HC�UW�C���p@��-�F�V�+es�"������x6���e�#�}�Փ��!l���П'����-�0��c3@� ���a<"��J(��z�J����ѫ)q����<��6]�dy��9ab�2�� x�F�r�e������dۂ�� ƟHz5CcFD�8�~�HfD�c�ڏa�,'F�L�!�:�<���̬#��7ڇ _�A��� �*HK@`�$�*��:H�UM�MVm��\/Q�4�.!]1r�b�gr�O���^)��e��P�����v�l)�< 
��k��(�a]:|N�B�ZK�8[r���F1���b��i����kUq05��3�1���Q]�F��)���@a�i-w���а��B�: AM���1܎iѨ�Z��٦��y��f>-�Y�20����8/�� ω�qJ'� �;8-�y��f��of�4+�o��3>�<Κw���,±�[R���{}j�)���	��\��ueq��s�� <1�=��p�r���L1�g[��{"�F��fr��PjI��JLv�E	�g�󕒚�]�x��e�y�D���A@/`P�:�~�k(��A�X!��4���D�k6fh����¨��O���� �A�a�Q &��Y��([�7��ا�Eph�%�hRZm��N5pj�D�
�3�>h�<pfC���9��'���*�_��_�gf;���;rJ.���A�"�1�[� �XS��P$\��`���4V_$��'i�tު�1�}Ƭՠ��8�L{��]�� ��'�v��y��oXw����@��r^L�3,!�v:L<��`���uho��N���-�y�
"k�s4�`o@�W� �<gs�V����ҟ�js-���dճt�t�b�{վ��T�4���C�W�g���6���뷾H�N��KYO�,��y|ː�];��]\�,�+�9�w�[*�B����_�g���l������C�>g�����^��g{���ܰ�xu�����7��j++��'�*��H�i��2������=Ɖ�{a�=������a�V�F$�!��V��rFp��6x��{{ٽ#�~	J�s�a��<D�|l�>r&,�v��{�;�6�a+f�A,<�L��2�Ǵ�G!!Rϧ�a�J�d�x��|��d�I͆�:X�T$��=C�P�E!���(���:+y!�8Bt��_�t~������+��2�{FN>Gt �4��ٯ!<�.����3+�rb])�CD���5F�:粳�H�w,�@������(-����0C���e���>�*���M��T��C���hI�!�`�4���J8�%f�ͽ`H�i�K��̳/dϣ��D�]�r7$�z�Jkh�4��н�Pz�]g@��c�D��hd,奄m�	޹��4 �n�Q�=�����X "w௎O�$H����k,�UM1�ȇ\��.[�M�w0���ɉR��qDv
�v(�	�t�)%��-i�g�K��;��Kf��?�� �]�c�`�s}�:����}�H�f]lM��׵��#Rd:j�ϋ�5t>7Q�2NԆA���B�m4{瞔_�:��แ���F�\����|7�F��Q>CiZ}�����e��!�@L0���-z�#�sTݟ��3dH98El:k,4��Z"6��c>)������יv9�vbY7���j�ZC	L�A۹�1��N�
�\/t���:-���6���G�X�\:���*	�f���s�$���YڑGJy�ޟ�� L�����f'�xu��sv�a�r�Ik�]t��:���(G���7i�1�b�{�SO�0J4��^���J�2`rߪ�F��"t��f4��,]�Y%Pd�[�]�t�@�m��e�+a����w�~]��85�r�B��g�n�3[����,��

|^�ָ_��!j֦ks9��3�3��R��3n��=�H1s$�Q�Ptls�����	�tm;�L�yoK�vq
�lj%a�B��.K��B�e{g+J��7�}qO+
Vx
R����:l�$ϙ��+ �;g霔t��='&�ėR�ᰫ�y��Lܨ�����"Ȟ���I{��6p䓈�s| �ᙸ�
��_}����N��R�(T ���A6�)S�^R+���P��2��?
�*&k:ߠG�T��.1�͹��!��o�����������+�C߮˿�}]Xݏ��l�g��?4�g�{�����'Ǡp�����7����3���S	��|��Ofw�����P��@��gf��nf4]���$������?��Ʃa�J��7*V��4�<?>s�z��k�Bm��ϭ�{��z�̻������h2�jP����jo2�Y������|�y�k[.��f@����!#ۇ^&YZ��^{�V��7?�J8���L
��$�Þ���u@n�}�X��w����I?W��sE��ٻ�:�F�(�4ð%��#*ʀR��&~COQ������B�K�Ct� �� �[¬�)��@[��t���B�&�AWHi�c0� �B�s�{f�p�Eߟ�Z����	��yL�_�R��,��f�Qρі�j,���B_��4�p���?�����ˎ)	�0"j�ۦU82/�!��G��ˌlyuo���{d�t^j�YuY�'=����m�B��7�G鄬����(��G�!����3�2`��0���mH���>�Y����`�rvo�p�k)á���������X�2���=��̤)�`A��~���§�Ւ�0�N��2�`*�f��p�?��_`-���dZ>#ݖ1��"��F�yOI���=}6s�
�:z�f��4�R��n3���}���'��@J�sH��ggIZ����z8�#ʒj�m2�Ҧ��[ ng�S}'��Ȓ�U�5��--O��u�Sb�Jt7�1G�QP.o��3�u|�lr�x/��ߧ̖3[�?e|MHn�!NA@��ǿ�}[ϗ,�O���j�_�;�����f-�Dz�Jd�4r�l�xI�%��[V����uqm��0)9"K�a�ir�C!�%�u*��/ZDJP��}9�Hf��Og���=(�!��2yt�Ej�,Hȍ,	I
����C�
�.�f�� 6�K� � �N�N�P#���"?��{j�uZe$���@�N�.��C\��{��8�c2���
#�{(�iIM ]%��y2SU�1��Ρ�jp<i�?b�f�Us���1Ġ��.@5�oC�Nu����[�6Sｪ�s?����t������r^��]�X/��;nh��oS�^BU��eJ�g3N�{�Q�M-{�Bp��I�ͩ#֞�t��e��p�mި��38��rO)svZs��tz��)r��z^����`����b�ر:{ڭd�e�Wb���ʄ�xf��ϱ&6w|I�a�R,�\�'���� m���-�1�: ��gH
��d����*ݕ;I� k)ـQ*���c �6v��gQ!î(;d��*	��u�.�&b�t.��t��ebu����.���B��Kً\�: ��W���N]��i�����1��y2�����_�:�d?���ѣ�S��d��f��-u��30G�0��Z��!A�K�x�N���ײϼt!�MP����H�T𛫋�jc�{����<��z�XYm�7zչ�NnB�K���Z��<�붖'N���D� �E��˱��2Av�spw� ��w�����K�LD�u@ڼX�B)�8+T8��1�������ʕ`����nݢx;{|��l}��
������ ?
"� �WRd g5#_�U��D��[D�
G���5�ϑr�qPM��Q�/�Z�{�����z5���"�H���`+/'M�ɟI�?�>�^��������sV�j��h�>��̇��������B�V)����~����IT��qF��ql�T1Pcy.�O<���
�w��W���ƌ8�:���c"E5}jQ�ȓ�+�mr�pl���y�Q�y�-�D�r��(��|��h��;�rdAp4!��}��]���f8yy.�j�����XNp���`���x_|�2<��e?3 9ʠ�pwa)R(Z���k�P}v��w��cЍ8k�M-k��L�kl쾔�kY��ݡ�f�ۭbC��&��b��|v}9�\�Y���B�*�/5�!�թ��zs9W�I�=w�!뼯��@gi�+<���b&��N����f-i�@��øYXQS�Ȍ�u� �����e=m(��f��N'A��,C2��}7a��?�3Y~5QB�0��:P��O;�F��Ȗ	�y�c@��� L2 �&u����ǑYN�����!z�����tp<7π]�b�*�W�����g@��Ir�̂�y^�%�	��^W��0 �V��2������<\x�b��-�ۦ��������<�E��U����-%��Yp;�g�$e5�P+�3m&-���#��l��Fw����8�6b3Zv�Y�둱t��ߢ�"���S͜�!���3?�Y���6α��7/�q⃟��j_�bay�:�0ap�sd�����s!gRm2�}�^�f'-;�Z�[;6;��Ȩݥ��g���Y'@2�2|4�Xz��<���q��
��g�����È��'3�DH�}9��|<��)	�5���#��|��ƙ1
#�� J�?ˣ:zm�.����d}b�)����&�-$H�pīHȊ)u/�4�%��U����$���,�a��z�bwjd� ��B�Y�a��"�c�����l�kp����UΨ`R��ɚ�k�{&�Ft�_$p����:K���F3� ����X��<�M-'����醭q_NႮd/1�Dy �C$h�^���vk'M-X�����r-|�����/�ˉ�������Y����o���>�A��6�u�����ЧL-g� ����#��������+��}��x~H�`;W�L�ۇR���&֐B�X�pf2�;�c�A��G�L��P�w�W���/g2iwj�X�(���N�D]���a{���kofoܢ������s��œ���V�Z�7b��2���z�����/���ˣr����&�����W_�>��R��z��赴�g뎷�Ș�x�����8�[���N���|� 8>��O��H��{U���׿�z��׮fw[�  l6f�)�:P��jFKn��Tꌨ��)�J�`����$������V]ޓ!���x��a&U��Nk�}���!7�>t�d9f�U��UJE�Xg�EAcV�����
�|������W�O[2�{�E�j~q={����
}'#�U�b��JEf���p�$���s��	��Ƥ�<���2:�y�<.3b.}��P��%�I��}4��Z��d��>-;�4f���g��:^�3c�ZG`�A�<��hU��Pt��l]E�E��>��*���6�?�Ku��m&�[��)�����X��(��E&��Uՠ�'%#�ѮD �1�G�D�X34j�q�~Hqr}f��l�QĎ�4���=���}�7rt��������E΄%Joˬ�k�"HEJ��3�"fsm&p:��QI�X�ZY��#;h��̤<�OrK�� �}4��|33���|�}G�*F��8xX3	��{��f.r��%F�>�������<���-{���#{9M��g�_Uw�x��DP$��̅�?q���y���:��\��0�z��4��d/�iVƬ�C���	F`8�/���1�sԑ�Z#?���)66�s!���|a�gcX2��Y3��tє0¾�̡�=8���K'����u^�v�q���0�1݊��u�De��})1=ʹ�{���&�`�W##���݇�O��etπ��JQp:�hvt<�}I���z�9��J2�>z�|CAP����1m @��(<�ڡ��o��c&����5�����ly�y�"���p�=	�|���u�	U�/��7�L�9Њ��-�����˿>�G ��_�;! ���̯��ՙ���#�����,�YV9�?��?��?��+E �t��]ͬY��A��Z�f4jE3�<4D�;�}�*(�B��/2<� ��+4�X�v�V���ܿ�m>�5���l��+T���69�L<a �	]�C:$����ك������~-�Zv����&�C%t	Q'?mX��e&�GIQ1�����6�{�{ֈV%��eX&vC:>�����t)���f_�ɴ�����e�!+�۝�s����7��%�y߯I&�3�|���7x{��孓�b�7|aT��Jԩǅ���]����>���������3Ds��I�,m���"��h���K������z��Kl~�t8��c;��_������������	UGpne��@���Qqr�f�t�!{���h�K�_)i�8��(�H�z��|A�Y�p�+yj�4�:N�� �K��l�����1i�=�X����_��h�[-�/�˿��ݿ�k�2Mg/<I��|v���.��{�%T��S�Dؒ�I�nN�d8��ɖJFM3a��1�A�Np��夂0XW�ZC$��_Q�ST+l�i�5���'1�q����,��1�L�`GB��7#Q�h�8� � �^L�#JЧ1�a�K�eD狁�s� \#G��2�O��4�9?�k�o/eJ�+	�sXqM�8����Ȟ��SǤӍ�î�#T��k�]��g��D�Cg��-*o�U t�@X0֙	8�]9@��wQ�3'�1��^obe�0 ������U<5qB,��܌*��0F7j�u*ي��{�@�\>R��k�����H�>C�>ȘzbFiYL�nP"*r�fB<������\�h�����%1߁�9@�qO7[�(��t �9�:(��k���(Sz&��x�� �l�P=�ٞ4%(%X__!�b�	����!��!e�'�И,Q"/���C0_<Ϙ�`��/��!���4klV��8�i�����
@��P&7F	իӼAO�ױwP)�.�	�X����& �_�0s�ޫZ�f�B^A0Ǻ����<\�)B]� ��v�̱�=X�r �4t:&��NQ�u'�H.�؋N�������Ϡ|� M���y�P"�{~݋�����%Nk�Y?p�0�E�L~�6�`���ip@�`��h /�r0	x�f�:M'I�(>-�1%^�ԃ�1@����|x�ˠBO�����3� ��l�&�7�Bs�b�蛏�%�8�>�Yugf�NW l�������]�T�n��E��S��Ys?K�Kex`Cdk���L���z���O��?�]~�B�u����P]\�Ȟ��s��r�>� $�|}y/͡�۔�W7&]a���W��^|�>�Tv���f;%��ͭ��<�Yj�72�R	LN0];�O�LcPXҺ���=2����)��DGS>��u8���r���^�^� ����l��L�ߧÔF��֗w�[����=��?������׏��>O�-�?>����ç`���j����p6�a��]�{��ǭ�sh��|�ǲ֘T-����������&0";Dx`v��g��Fb=�<�am-�C���f�y�^v4�����.輲 �g	� YhzK�t�	�D&A3���AXt�$.�:)�"j�xxX�����P�5��g����t�5�C5���Go�A6"�p	M�����µl�6���
p?�?��������7�\�6{:[a��[��p~��/���������fAX$�Ĥ[�Q"�K �"��VP<��#�t$��f L��s��)���ƃD]*�r��:2�I�C�]X�~�4H��<9*���͌����D�	�p2��<(R&�?�gS��k%�0u������pn/���Q!\J�I��s3c��LN�K �d�NG�(�VaTP�>g팪C�R�3CӞ0��)�;�Q�ĵYI�?l�5�f "�����~�%�5�H#Tt����eF�,��>@
ܻI��r��Y1���_�t��*/ ��9vʲL��f���K/T����I.��[���ϐ�)9v��i�1��yJ5��N]��I�\�r5���=1�c�����|�:��K�������Y�g#Йe ,ʙSwPGn�O�f�]��8؁�4�tD��(��O���I�ʙE��T�#��(f�<FJ��L��j�n��\��;v�)���^k�2\u1��I١ !�����qs/J�I�?x��E���Ȩx�f >J�v�PM�3fke�ӽ��2 =��5��F����
�z6�xoK�f����Eb+�����=�SP!ϭ*�M��Csݼ��n��JR��&,)(�vb������M�g��}�~w/�M������}3�~���F���sq�	�E�<�<�z�i73 vzv��Yz��)��{~y���ݗ�}~ ¸�x�i�~�!�v��H%K�#2�3Y���ڂ�~�{\{���=	�����%Iv��&�`���}6^o���xƎuU��
g��Sv������u��]�FJ1`��؆$ĵ(ñ�ݼ�ξ�O��Ҕ�?�"e�Of'�7	R�1̽˓Q�!rQ���� O۔C�\["0`$��>���3��g.S��e�|���w������:���Aǲ ׍1��';����կ�짟�N'����#a/�s����Wǅ������#6�Ϸ�
�N�C��.ug�&�kم�����F�Ҹ�v��1dq����qtCR"Q8����H�?�����{�d��|��ۅWQ:ǻ�g�P�^�U�-���Tn#�q�Y� )<S�bbڔ��	���u�0 ~%��@\�vf�OA��
�V�XE=22|s���'5��LJ���⿓]~��@6z 9xv�=�����_Ɇ��kٹ����e����#��dTҐ��uy�R�g~�Ht����@`$�2/�?�=;@�a	�m#q4�R(k��<"�H��wq����aK�!>��Ŀ��q;M��+Xt�r_`�W�,c��Q�J���T,��Wr\�x2~a��8����sqBF�~��=#l�3��i	�t_��2�Q�W�u��xt�^���ҟQ8�.��	�$dHʄ�m���Z�Ftl�CjIg�ZG�5���C�B��7�8xs��\Gj ?KyF�|�V�'*�*��Ĉ�(�kK��d��Wc�D%=4� �Mxe�&���cyI"� �5�t�N�X�{dQ^��q����P3���ʳ <)�iF��T���%@3�3�Z	�����:�\yGf��M��s 5��b��͒��$��q�/�{�������(:wW\=,�7����!x�9�轎�,���:��HJ$��-H����$���©�]0k������z�U�!7]t 9���TURO�N���(6��}.='���p����3���>0���?D�-�0�'@?�u5ˉM4�e�ز�Dw�"�I�`����Z�4�k�F�}���
�i�ZggլR�|����=N2 ~.�/�ϊ��۵�.�Y���]��{��$F�)E�k�=�-�SI[;�;�h�\r}	�-��S�L3O컰)�N1Vw�59��~1����j��=��� ����~�f��}��h�bg��K�A�s<���G��=y�g��E W��������9w&�|D���q�Y�����������.!�1"��X7�������c&d^F�f��03��d�Zd��*�i�ؤ�=B����;L��;�Od�|�<E��ص��i��2Ћf�ͪ�1O���˩��K�e�_@W� ��׎��n����A�lH���ר�g�f��A�޹��?��/����K�>�_?2�:}��;�2��>�&�휜`>W�,������������}7;�����`l1�\��.��kg#թ��s���֮�pc��h���;�ͻ{�n���{:���o��6j|N��m�g�A�5;b6H��4��p����!�^A�&�@�C(Ɠ������1i���gg�
uDz��}��d/=w9����f�?q.;�c�/�u��*�����'.f�/�r���L�^�����-�M��2��IG'H� o�s��W?���8����(q`3D�%��gD������P6 ��UHQ�@)԰�2�N )#"�a�G5�@	QI%G��	$i�NP"���ZO�c��JlIO)	K�@2�,�%>�nX+������ٕU��~��9�,�>��d)N�k����oy�T:�P?��M麦[����P�me��-�@X9X~�屓��x:FD'�����Ė�R笜�1��2�V,�\�\��.��T�J%U���e��=�y�.��Ō�C�B�V�I@)���j�F��3��*W.B�-޻@:���{�) ��AD��R6�$M'�OǤ�iA[EM̈́z��:ƙ��sN�n��gdh�ɓ�}\S��RG-2�V#��%�E.8(��ʆ�LR�͊���|����$2$,�X�(U)s�S2�7sz���ٹނ�df���W*�uW�?��"���tm�N7fگ����%w��y�Xj�E&8������5�2X���6H�?�ˉ���S��}yO���u���LY���N;U���eKM8�{?�̜��/��(��d��X�g���S��W �4����w���Ȉ�-�&�*^�i���� j4O��|��,�x!Ck�2�AUp�}}Z[�ì�V�6i��.��!JexV#X��#�4&K�Xs,/���sMA<W?���5�g;[fv{>k����Nq(W92�){��@������l�h!wk ��F���x�6^�Y�2Ƌ�0�Q��\�>�;�8��d¹��w� �k��Q����_ w����Nx��t�k��B�e����{�#��)|V.��2�w��Ѕ3V�.,�=���{��d�^���t�B���s�s�^DJq�9x�T����#;W�q�c��+a�J�:0`$�kN��֣q�3W_�����>#�*��#�V/R��\6��>��������?��~q��wj�?ο�HA��R!w��h�:�x�7no?��k���_z�9��w���Le�����kw�t�ܼ�h�R)��.���\�C$h�VFW��}|<��w��펷k��l[}����P(��vY�@�u8f�Y������4���H�`��ip�Ϣ̈�4v���x @#4���$�!' :*1:;,9\C�m�2�l�>�V�l"�t���_����M�ffF����8I�uj�s�l\���c����տ�������ʕ��`�`�8
�H%��;Qk���~���nQ�HrF&չD��;@`�qX2|�@�E�!���3���@Z��ѱfu���3~V0���QZ�?���
�)����J|�x;*>#�kw�`+����]��(ך�m�F=����2���J3Ge��oZ֢IbЃ� ��0�]���4���Qv�D��Dm���;|C�Ty��Cs�?����G.2y�)X�cVr�F8��J�U'F�P9�0�6{x;3�|�H�Y4&yJE�G�O����30��\3J'�/�HL��9�7�u58�NXg}�uL����z۹��\g`^l�bF)�~��Q?8U9P1eb��,�Jtb��8��aE�Ɖ��R��m��b7��u}���lf �DTۇ��G����a�Ev�_��U{��뢜n�-�,���s�"�^�ү
�SYP�����#��J�Zpf8������� �?�n�Y����M��g�4�9�����H߾_�S�aL��R��H�N��)�H�\�4m����h 
�x������2�������NO��g��(�Aj+�4�٬	��],�c��C��I°A�,k�e��YQc�����^�YÕ<��E�a셤�h��{��>�h���-��ʅ��6�fi�3h��O9d�X
��af6��yvN�HY����p�(�gA���5#Fo�����앭����Y�1�0m�4$�B4��"��ĲFP�ϝr{�$�젽�:Zd�N ���|��z��oZ�Ҳ��*�wlE��o��B+a�,�U��.�W%�9��a�6�\y�2�h��L�Ui=�3v[�}e`&�T�h���m��|��ׯf߻~+{��٥K�J�gk�/�e^.�eDX+� �-�|O�
q�t�6~���f���C(�ќ�!�_p�:��spX�[�@P���}�cV^���6������ל�x���}�P:�G{�o�����������`\z�u�^�r��(0V���6��I�DXX�1'�J%�yT[��D%��ɸ�̙6!W�?�����4�@�b�<�ݺc�.K�`2D	YY��|h���ԹY�<�-����Q�$g�a(�T�H2G��(������2v
�Ch$������A0�����	�}�%C_�^~����g�V˓�=[fq�gZw,���#�u�yt�#X�qk{��իX��R�Lɏg�S(`�]��a���Z�B/�9��3��p����)���$!uh����i�h�q��1e8̖��C��>�UJS8���k�Y�z�e�h��FR'`sp,o�qƉ�M{:M�:e$L�;k0)������i�F�=#�_>�h\{���=J��ޟ_frMf�T_�`Y��Zz��:3ާ�f��.B��L�@���KD�)�39��i��>Rv0�@tp���BK�>�)Z�5dI��"��ݔ�_I���w�����r���A�;6{��p�ғ0�	[:x^��w��R��σK�jِ��[d5�w��(�r��3q���IeE���"˖�G���gu���i�{�x����)�s
��i��8�~�p��>�y��HL������R�b��\=���]'���Ǩ����a�b=x��:E�|�>4/.�O��(r/L�A�=k�̘�%��,�X�	8f�F�1�Y����hw�?�7'���ݔ���4�ю:#�������O�#�t�Ǒ��}�sd�IX4J���\Ç�c����:T9�g�-*`�p�fXY�6�Y�bm���r��\}���|<�Q����fF�M�sʀ�Q��{�]���}7Srxg�_�o)�9E*?�ǐ��<�S?���ٰS^h @^�	՚�I��9�m ���l����v�9!�B������s�F�|Xg��\��Z%�{��f_�p������}I�lF��Ͳ��W�/��j���<�
�0v����Ȅ�:��{��t�F+E�j�I���э�����E&�`)J�	0F�@t�ʯ3k��0�`������:j�n�]ۀ7�eT�vv�j�ʒ�4Y���(���Y۹�����YŖ;h.�.�=�L����]�(S҉Bӊ� ��I�J�J�:��T=�����6�\T�li���ב/�g䀒L��6�ζɨ�	>���#�b	=�ЅΡi������>��_]�g_x��߾�\��dja�#���NW��;��[��V{t���}JT��񠛟:P.��Z>׷B��f��q�h�i4�!y�+��q��M�����RM�����ƹ�\�6.�Z0�" ����zf>qL��0_$��ȷr����I�`�5�(`��S�y!��k���F�+M+����5V8�H%�8<Y:ǈ��͏a�`&�l�dx2�HFY�����z�Ȟ�5P:�>Su۽!���=p�:[�n[W���8�#g5��q�\*�2B.O4������C�HA9A3X���4���1�ӡ:V�
S� ��� c��r!����1��W�gV $G׬����m`��j���"�����ݫ������&�frMG�S�5|���\��xf
��Q6��hWQw��Rْ-��(a�g�G����ZP ����~�L��&�^�N'z8�Nd�|�6���rp�f�`�8ٹi��Lh!�e��o�:������XBv\|�o�f:%��F�Ρ���C�� W��P�IÊD���f@Kr]ޚ�|����`2�a��p.����3|>@ۜM�lxW�z������Bo��F� [�M�;�;�2B0U�qs�8K�3����"CL�i�S��:D�g *�c^Y|Ɛk3�sŁ�Ly'�Y���>�Ϳ��J\g��jI�:[�"�7�Q�$�����EJl ��
��2��9���y��}�8�\Z��Ϯ�.�!@���;9�i�*+e�Q��1��kDe�S�����F���B�>A��2C�xl܌x*9m3,ܞ�Ri�����G��ͼ!=8�ofoG��b�4*�'�x�<��g��JBh�f�4 � <�S���ȋh�4��ɓ�������$�lzHW���]J�T���9)������8Ru��0����\�q���+8U�����Ǥ3+L�lj=!�@+�j*?FS;@������N���}���Tľ�<i��Yl�S���i%o�?�f���hr��)�3q�#�g���,��:=������g��w���]ɇn��y�t>G�^8���!y����Y_��s�X���\�%F-  ����/J����$���).�T�#R�Xb�0֜�X�kw� E�φ\0@�exḘ�8�S	&�ap���U��LyJnY�Xf�{3��Ǵ	��<��wV�!e�q���
b�\���:��եZ����[�>��kh���'�,~���	��C7��N?뵇m��+��4R#$�pZlPJ3�F��q�u�[��jfQ���C�35��A's�D�I��>l����	VC�䴏р3�p�{��W��z�Id"N;��8�6��,q<����}M.E!�d�����1̎E�Y�%����b�:�vh�딸_@v˃$��7N�N��2*�0,�L}���A�P	�>\ь"0�m�QA.��%+<9�) ��D��C*/c秗qU@�}��"�3s�E&�+��1?�S�f�̆��%޿��Z���������I�}�!-�wx�0�Hɹ��⽂�ʿA+�hĚ>�Xމ�
Ҵrh���Z��hW�Fғ�S���q����]��i�J���L"�# p�{��e�D@ұ���g�~:� �|>� 8��ig/����yy�Y�&>Py��� YCfQT���K���rv�qbۥ�(>��������#�����k�z�G����ْ�4�C�8?%���-��J��mj��5��� 7= �YR�uҢ���LY�d]�ƴh�0n���'��H+�ya�� =��̳�����8��؄�ߛ���O|1�S�
��o�C��=买洝h��� �m�A?˝
|8�'S�@0���=in��f}"�������Vc�g˽���s�Q��5|�F��l/>����z�$ߠǍjQ�%a�.�iV���ru�l�6�-t�8�.�W3�;f�F� b	*�K����Z�3�1��I��CS�^+
�x$� ����s��W5.܃����~�^�������>\{�;�P}<+A	,h�6����3�V�⸮H�j��چ%���'�U
ӎ�~�Ŝ�J�%�׃�h��92Rp�L��/x�+>H�=m|4=�؅���FV7�Y�t<f�A�gY��Y�p$�Z��������ڦ�f&�h�<n����h4 9�_�l�!��������
�ؽ��t��݊�gQ�����K�U�v��qF0�9gY8���\~�2�~삷�<�>Ԝ�^�������j�FW����?�׍��`@|�s����q��g�Ŝ�Ѡ;��B�p�C_��Ԃ��=���"w/��n����q�Cx��(��`R*$�<0�5a��Ƞȇ�� ����<���C��i-_�#VcTpy�ϓչ»�||����߸��~�E������@����C}� ��Pǚ��e m�d%�D@9|�wR5�0��2ͤP.M��=`� �k��P�C ��g^d�VG��2X׭��E�fu4a�Oy����	Ș��|&@�LR��(3���W��0����R�S;�@� �$��l����� ��FZ��0ؑ�3���_G�������g�? ��@X�5A�Sp�u(������"]�M�;�� �B��%���n�e��{�����E!�ކ,��Fc������n�jDռU �	%�1�űpWI�q.�j�zD�~�e 3f�" �����([OV����Z�8f�oיO��Ӭ�T�c�0�J d�#(%cB,ϽAR`�
��1?�� ��:<8���xG��_���Q��-��~ƾ������H� �=�< �Ȟ3�'���o�#�/y��"��Y:��@�ǋ<:��vii�O�¸�X�?�g2�;	G��jo�: �ڞ%3\f�Od�5�����x��ڙ4�)� �u����,9���%���t���g��h���FCS^�^���O�SI�9�x��Kq Ó2a��g�]@tJg��k���8s?HzF�3���c�D���,B�C�!� ��g#76a(;�.���$��#�L�N�����1�O?j*�w�k�����zJ�:w�3sv'����fq�zpZ���<s.���*��P�$} ���z�{����E^�� ���հ� �$D#,@����'jɋ墸o2�2�ޗJz����O���)3�������j�^�+���/��:Ӷ��.����'+�A�TӵQ�|�	��yΪ���1G{4)�?�k�o�]$G��f�, ��2TYǹc�1�W�&����>��$�r��>����ED��}HA0��gӉ(�cr#&�����iQ�fT���
�������{���?������o�N�c�fkl    IEND�B`�PK   �cWL̔���  � /   images/37b4a41f-4938-46b6-a864-47b2117c0019.png�uW[Q��K)ŊSܡ@����ݽ��[��R����k�R��$�{� �9�~��>�#�?�1�1�HF��Z{�k���V���,:*1*��)u8�7W��Ȉ�����c��Pkl%%U�$%)Uݜ�l,��|rRӑT5�����ã~A�s~S>��	
�<rH�WI�7��d���O�b��Omҍ� ���O���#F_�Qu<L��@�y�'`����Nwr��*�r��pQ�%�oD�:|�ా_~z����l��;�T���n ��k��ݗ�'@L�X	U�O�pR얏���v�N��{s�t���F1��z�sb$E�k"7W$i�4�ncD(�������n�i�!_��&��������"�a���	�ͬ�٦e�qc���Y*��*�Ln߮''�d��#�|�5�+�J�ȍ�i7�*|�E�}�͡~��5��>(�к���?�F���}ƭ�r݌���q�}9u�ߙCOK[5T���Q��8D��E�9���B'�j�M.����&���cz�-��M�u�y�i9T��<�%����j�yC���K��#j5�r���g�~�9^AX!ݑP�D��1cd����"�����pJ�>����8��=F<����/�Q2����f�@ko�]���`8�z"��)/s�Ѐ3��\�0�R�U�
���2K����&��8lOK��ؾ!�|Cfod�<��i���[Q,	�Qo߿�(���:`ʯ�#ư��*��~�v��5�7��!<�������q��9y�Vx�',���+J�a��H��;H��6UI��J~���	+U%�D9	9*0)H��=@�{��W(~�~E$��"�}<tх���[��g>L�pp?�z �S�d?x���4%� .&�k����'��0T��dU�9yM�*R�0;��"�v5�9�#\�ز�L�A,��{��SLӐ�ԃ�t��<]�q���-�i��h��r��?����f�f�ftg������ը!d�ρыȋ̋��c��I�R��[���M7鎓Ɏ����Y!�������틯o�H����ߋ~��UED���$.�+� � kC�By�+�(�Q�Ğ�!o�TCɃŊC�������d&[9�Qz�	?XR���,�sD
����?�ϧY���~���,/Dٔ�.�)�+qW!�Ѥ�ň�S�A���aUݯTQ�Gۊ�UsB�EG�,@�7J� K�_�ܓ�5�/�/Q�HB�QEkDU��Mu7f�]+�*�*�J�Uճ��ݼq�՗�����ؖ �4'����ҫ�+������b��%�V��Y;7��?3D$��D�q�GG��~�~a��טĜ\=��Ĵ�����"��O\�\��<�" 	{=�~M��4�v�#z$��L��)@�7���g�]�4�ա�-j6����"	6���=%Z��+������K��M��9Qc��y�z������J�Z]����]/B.� m-2�*Ί������T�͊��Й������y�dq��2��5ٲv�D40>�y�f�8��c�g�7�X��a�"髚�k?N�G��Ӗ���C�f�=a�&�eFp�Z8ˌ쫑�����0ݚU�R$�׀~�c9��D�$��X�dm�`zR}|ƧJ�H���������A���ص���ۻ�_�;Z�:�����ԿK;�j^kn�5�q�Q�&�{?\d:�X69�>�=EZ͟�ȥ�iu�ΏA�4O�\I9���\�8-=�V]�90��]��f7k,F.�8�������1���������
RJRyDLy�<E�́O{���/"�j����e���&ez�����эr*|�������lk�,s!Y�r��n���"��c��,^N+U��N��GzKMQ�K���P�vR]�������Y��/���*�p=��зF�8f��Uߵ�#��0�#��qX�k�=�e��9�}_�yN?����zW�Gz��	��\�'I�i+ᯙH$ �E}�y�����X�[9r9K���d^z�2�ҟ�h�|E�Ӑ�_sGs������3�3$��D(D�U[\��eN{��,ѥ%_�'�Ɩ��?����$�7�|1�0��{eC2R\]���4Ӣ�M�[|���&Ǧ�nǖ� �&�=����R�F��:V����Mb�6du8^;�k{g����Ɩy�a����j#򞺔�v���Ծ:X���}c�B���E;��ȼ����+�R�l�P1�����\��i��}�at�JH������<�k+-�;K-ƺkcی�?ׯɬ�-��#W�,:�n߰�2�zWT{ۜ}Z�0+7ݯ5Z�&��R�=�?9]�m(�,)`�r>]�~(�y>��w�iW���@�.��B�ߞx�xz"�b:UDB,��"�(�|`.
aZ�y22��.R^;�( 
t�%�8Ϛ͎�2zz����R�~ �2�#�.E�~Y�@���	�q_^�\����Sv>����L��q?b�>���`��\������� +�IO����w���1�t#�n�KF��{�^	�[�<l�͝�U�5tjY��]\⮆�3��;?��yD��/��{www���g�WB������bL(�y�P�Kp�Sɞ7t�dw�r����/#�0t�'{Car�>_-/� }N�=8�n*�|/֗��D�8��r?AǪ>�e�	|������;�z��_r��ے���8��>�U�]���'L��#�����{n�68o�5'27����;�Z��=�s+Q��|p6�o('������2(��}����n��RrP|Su�����%ڼH�4C�#�}�A��p;T�Y�+�R���G�(I�{v�\���F�[� g~�ҧ����Y����1>�E�М�dc�%`P��7���ڈ�6��KG�V�[�o��Y�'� ��p��� ��9�$b����쳗���?)����x�����BF�o�o�o�o�o�o�o��OȀb�<��t	��3}9c���߯MR�Ynu ��l'��;��A=u�w/�0�?��>$q�i���s�c��'�7TZtu:8#������P���>�"�)��Ν�)?8�Ϯ*x�,`��꺯�D��i4 J�v�����1���VِhT9�$���|��bY��CH���'˖�k^�S���m��!Vsh�[cY���lM�6���� +�����=��ų���s��Z�h��Gx.}3�2J��%|9W�xY]�1���C)��/��R�I[����R���j�C�#���܊tl��e��y7 m�OM����ܽY��w�v�ĺ��+Y�(�vtʤ����\��y-/K<���,&AJa~نh��;�/$!�Mg��������z��&�w�������/���W���*"��B�Me~3?�F�S�w������������h�I��Vu����fc=3V�	*�X�o6` 8�\����u��L;^p���̆;u��=@��&*Lu��<�e��ZZiZZ閻��W��Oۛ�Xz8� �����]�?
	g3�͇�8�;�fԐ�5�iѺ�˰1O��~�`�&�}%p��B�����݄�~=7.Z%����OWn\�*�A��\���p�|ݰY�����j�ϪU�V�s���k��5�t���wBԮ�D�/����� 
�m���q^i��gH �O��O���\��Ջ��v���f��m{FzP\}�&gaU�^��q��s�}K��Ҙ�ءm�{�!�Ni����39$L�{8���_<G<qC$Δ�����w�1���$�\���o6:��v�RGg�x�%�(	��.��LM�WKO/�,�$q������~����$��i�g���aϮ:U�iol �+h�l:y��2�m�ZS�C]���0z\fp:~
xY;ޞ��mPU�[g�U7�M|��ً#W��W1�L�[_����ӥ��������9A?���������9,��(��~#Q�D��Y�p�^R����k�@&ض�`�/[!x�lE}`%��SS��yX���,�*���f�i�A�����rL���KYӱF��b%I����&F3	��f	<�ܧ�Z. c?XN�g�=�e��q�]�:�7.ɒf�x���86U1�7���vC'�-�W|e�S�,�	�������)8�I��5]ʝ�uAn��hϞ���
_p��V��{�"���^��&ҋ)*"�F;+��� ��1V�a�z�k&�$5=]��y��K�XF���:��v�ķ�ˡ�>�d��v�R9W���e����fq����U��$�R�OW�v�զ=�,�]<<"Ǝ���2�l��f|Kt��甗���)�:�^�s<���
=�s�#Sͭ��Y潓j��ɒ��BC@rFp(g�Bz�:˜�4&���h�^5>�ߍ��e�+	])h��%��q1���ݨ���G��¡�4f��ro�sU�A"˧��tO�u��uK\��lmjS)�0 ��t� j�5ҍ��Ŕ���4H���5n��s�����iEj�~��N����V7��@�p�z��r;�(�\Y$I�a��X�j5�Z��&�wy��E���AɆ�������`�Y��yO�ۉz�d3�3;��C�5�	)���-t�X�:��88%ݼÌ��t6+m�,k�iʼb�xVz�5��Kϋ1(0dB�?&b��3HK��k�ái0_�R �z��^H�X�/����:�?/���Q,�X�&ZH�[<��N�!|U�����\vBmn��%N����eO���J6�]��Pr����ZQ;�1e��*�1�n���v���eq�Y��&/%K����Wk��3�A�H/}b�yR�I��vH��z�������v?����gU����P8)�e^�?���T�f�Ĺ%���|9�r��:��	fe�0��&�����8��<Vb��w=ʳ`����N&���E���:rdN7'���]R��QY�ɋ~��D�Au���QŷXR��S9�3E�������*�E���Zk�Y �-���K}��N��9�4�����i��[�܏RJ#�oa�#�<�#�]-.��*���M�I-#���:��$���{Z��MѣOy-�)(��@�*�j��!k��A-"����S�.���u̥�3��"��Ff������F�k�nU=-��q%���'������e�v#�6���w�şG�z�yN}�7 șs���=��(�OH�*�Ư�	���0@E}�,�@*�m�r���p�h��)���P��WU<~��tޏ(]&\j�ԶҨ�/���k���z2/sX8�_�8s��i%�*1��+�N)yܧ^9�mj��>S�v®I�Ζ���E����}�j
��������í�NlW%��G[��	�����L\A��tJ8����$�fE����!����dU83\S�:���J?"&?JO�I!}U�,S�"#N��Á%��մ����Ԩjf��V���Q�qb���r8Ge���ssBS#�Ϗߢ��FF�U�ˍa���i�7	����1V��nG���F��I����B� ##���fSP����	��qFe=�V-g���@�u�n����|ɓ��x�8��p(���o���E����ɪ�E�7�W�c�^LsZ��,�h�t��S�gκ)����P*�d*Q���J#�	����*D�j�b�D��<���p-���� Qͮ���ws
��it���n�4��
�)��Q�x�ȤrT'f���ťW&���5UVjn˥з�nLI@�5<XRIt˅F��Y)c�u{1b�7&�3��6��{�Ռ��ZE�Y��������뼠�yjO9B�0P�!w�- $���Ŗ�V�W�,��a`r\�Ԥ���D�e�~�����}si�
hk3+ HҰzޥ.�x�\\y�7,jL
�v��0N�7���D���ecg����
L��kPk��WLa�$�@޻j�V����Q�����oz�'K��w�霶��MM��<<�65xEq�:�o��5r��t��w�8����h�Yo�Y���j���뚹�!�Wp.����m_��K�Uөԅ�W���L�;:&�	�כs�'�W�	I�I��a���o�y��b���Hٻ7~K2Z$MA0�Jl}�+F�	��z������i�56Z�� ��+(��\��� �#q���l��%�!�H��UU��j�
��Rf�v�w�j���X�mR��53[!T��f2�eڇ~��O��zmg,�@��A�4�/��gw���A[yg�]`j�q���)�v��8��d�"��n��W�V4}n�Џ�6۹밬$�v�{;?���d�L�s�:�g���>��0�O2���yE��>*�˟	y`|b���mwE(RWe��W�p�P`_!I�j���$�y#�}��b�5r�^%D�s7-;�s<�w��b?���y���_Qg� �+k��vZj��ns4h�>5|�)�4���Th�ˤG��|^�F��R�3J�j��HwPt��{݊F�G:%�m�k@� ���y�B�fT������+�8�,���t]�^d?hF%���A$��W%笮�T���oI{����e�^ى]umZ�}/lMA�����Nsf��~�-����Q0��<�-P�u{��3�,/u�ذgΫ�FhJz0>�a�v�d���q�e�[�$��uMC�&~N�
�ܜ,{�9l�޿�i8��e'WuL�_�'�qDF���-V
mg��j� e��L�*>��o���h�D7��-�{n���~�m�1�.�G�9������9?�,��<[p���C³�����������CP����^�ݗ��_�Y���܈ qZ��02���-�E��J��2V��"B��V�d���۩�)B��<.��;L��j-����b�5 �L�Y7�ݾ��>��miKg�*��Oh�������K ��G!t54/u�X��-c^��0I)
x�W����<lAU��w���3��۞#�Y�L�\�8�v_V1ye�'��(������T�uU���-��+��Ω+|�u�d�]jE�8�{p��Z
��t_�X�Y�U�)�Y�r��8e��K4���O��"���F�����ܚ�Y���ŭ	r����yL���o�Y�/c7νOnMY5�D���m����-������OcY	��=#r�9��O�"� +�,����sd�|�S�q��O�`�wH;Z�F����f[%V? �Q�76BX3؃�M<�a>�����^1wi�+*;�� �H��o{��	�C:(,� �Ѵi>f�4y��$q|�!�,�|���u1�o_ߪ=�D�v)�X/r\�I]��~Ԫ�}��|W8Y�M��O5�߇ �N��?���{h)g�|���u�{u�n7w��K�z�6�nh��S�n�؄T>T��>#鷣T��B�E~�Ю���Q߹�縋�\�?���*�^��H?*DW
���?��\�0�n�����j~�����t>�gQ/0�pTUͲX�����֋:&��ק�6mU���qb<n��2U��ݷ�oKw�~>����G��a	}!$�~8��"�_)ʁvr|a�����G��?��OT.Cd�S}:ƾ��\g�	�Ϸ��&�Ag�U}<�3����E�끰��ݰ�W�!�۾�s^z��W����=��B2��J����oR��>rj�%�� �vD�n��+�>�Fđ���a"f� !��.��O���wX���[͕ڨ��jW�ZhR`� _�M ���k-��6�X��`E	_�w�!r��Cw��јr��mC�lՓ�1�Wn�S�k��ay~vɡ�5G���ԘM��N�/�4�&<���c�?�0�7#��e)=�_�wO��O�e�w��ϕ7�d�i���	�+j������R�_d�A���ˀ����yc)�:My<U��Un��P~�x�r����h�'4�5���^�AMý�u���!�4���Gݻ�?6�`��[��wt��Y�yC���İ�7Y������^�5���<9#mW��I�=����=eD�e��s�KWZ�?y:Z�w�u�d�z$���<��^1�@L��ė񭋭��bq`NH�~ygr���7R�%^�}u~ej���~9����4�JO*�
�K]�d�#c~�-��Cճ�>��m ~Nq�օR����-z�3*�p���Y]�;q1b���>���q�RoO�ߴ��*���.1m�
�|rT��eҟ�yv��2C�K���ӳ�ĺ��F�g���\,�uT��N����vf٫(&Z}�	��:��I~A";�!Däo�:/�:��_SB4^�ͮ���b�s�_��J�,`o��>����΂���l��>�P%Z��R"�"C�5��e�}-��S|I���9�`T6�_Ka����d&�c�{�^�;�A�"-����yw�$��&SYc$<r��ʳ+�y��#0F�<cljJ�,6�U�Ҽ�&���$!�P�L"���?%��3d!o4 $շ�u�����Ō�˨{����������hd�H虃3�K�<Yk�O��O� u*�hO�oՀ�ȯ�5���_[��m�c���x���Ƕ�� X7�\o��x�<߽LM�����%TV�����nØ:�3%�LMB�'�)tq�$���Cu~V�VAK�,K���7ԗ{J)&��r>bc���Y������w�@S�ٚoR<:��xC��B�.v�A���������|ŭ�G��+ϝ�Z���_ŕ�U9���w�eBm���������X��:)�݅^���#s
��9��É��\�S_&9����e�'���W��݂�z�0V���J~ò�i�����$��#��!� ��q9l������+3�؛V�qE��nR�0v��Z�?��#��@���%�=�$M��&��NC�p�EW�ɷ�y�,lK�� 8�ۃ�KXC�˯%��Ək%NP�!Sf���\�KSZh ���&'i���X:�z���{���ko?(
p	? \�G�!�j��e O����YO���c��U}O���yW~0�	�n�lN��x8��"L���(�VH������*����&Xז�H�b�eA.Ġ��n����	6�.�.J"����:�"�y�W�H����oJ�E�I֍j%�{�BI�τ��3[��¢����CV�nol�|�޺��`�Z∄�ޟ'jT^qw�P����ɜ�y|~����Z�;�酧?]�.�$
%G����P	F�����;�.�# �h Dܔ�J��i؞� ߉�#�B`v���9'�
(.�M���w�aq���2�S���ྭ�3��n��*�UT_�,���K�xf������E�R,l7��!~]�9�W����N�?�Y�f4o#��~#�sek��V���v.�?N����`EI��V��?M�_����B7�����%��Z�˓E��&�C%&J%1L
�6����Ÿ�'�����>�}#�J�7��ՃX�]�Q���`l��m9wڊ�����&dW �bz s�HQ6 �"�E��QY��'5�����n���U�[
Μ���+|�Rܺi�$8g,�K�I���y��|�Lv��}�݌$�z� hw�Ao]��4X�䀸bǄ��o�yRĿ�K�[P�C��"*�zQk��}����`Iff%�>�U��7r��?��ڙ���6grڊJ��7����̮@�:"��g��`�H�a��t�S��m��i���e��XA`���> �%�jd���#�o	���r������mL���.�p�N4[���(��7�e7؆O��o�m���G���;�p�Լ|�W�=$G��Qw��	��(���c�񯘩����'���t�r�xS}�[����oP�������1!�N�(�e�e���;(T�n�,3��C��F��gP۩M�$w$��%���\ƺ!Ov�l0���]�6R��	�M���K��m�v�WRh�t�䀁�����g1��[�}Ķ��թ��On�T��Y�|lY�+��E?���E(q������;�o6���#�n���p�^�(F�m�s?����Ol�W6��=tʚ*�]�_�X ��c+��ϒ~���W_�|��X�m�aZ��vI�2��c�����cVrT���?��6gE=2
'�QF���y���� �p|(�dv��a�#cp��rd��{�2�.�v�"�����F�m�ҥ��c���%U��*�pL��R8>3��^�w��e�������gN��2�Q�����s<Y���>�Io8����D�N�8IPT]�5�>t�wTY���	�Fh+��j+��n���� X�q8n�cr�W�;36ph�&A�(b����t��'���:�~�8����`�U�.4����Ǯ5�I5t�elj�茔�'�.�mޔa��ɝ�`fdi�=+�A�����z�jp��Ԧ���g�b�nCU��j0㹭C�j���$� gdW�'Gk�a��l�>_�Z{�����Rs�������f���u�Nʾ����'��ێ;�\#ᄽ|�ǧ���F��U����r=A���LttOh�%�%3��:<�FwX� ��a�+�3e��$`}�I�9r�)�=瓀䓗"P�!�
ߧ�����/�uk�u
(��<y�^y�����)Q��Yi��:~��)�dy'r�$�p(��|7���~qi=n�����=��N�?�^=���A*_�:��k9����Ǯ!C�M8u?�VW�w9���>پ��m�?c���o�{E��斳0������E�d��J���u޿�IP�%���=Mi��Ia�!G��Nn�
���H㽘d�@��7���y �pH!E
GɄ�	C���@X ����q�_��Ι�F/6W�tϙ�x`j�Hlh� �+��pB6i"�  :ςi7E��S�=�a�� ��) �J��Rm����k�+d�Nkx!�m�w9��� �:�s���)�$��G���G�J`��8���b`k����_6A��o�Zt�v�K������ҫ����D��k[�\�巠c�mU���.��Ft����U_�l�neq������$�Tn_�7�j�t���.1_��Q%�BQ�`@@��?~F�`ڙU�G�{?�&��i2�uWX|-dc��a�ײr�9�C?=j?\�\��qZ�����Y-;���>�64�?P^�![��>���oQ��uHr+FY�����P}_��X/��Vz��Q��Ͳ5�;����Ab{y뱼���	eNE�5k���?�d�<8��n�	�+v����R.&_�u���m4Rhy:_��%^�g���;S4�n�dɴ���\~K��U~}�]�,��9h�O>\D���e2���]�N���x��&7���7�)ݥċl:�0<�/�Q�-���DE�η+�����+)����V���X����7���A���Q?�Xq��v�B����2�����6�#r���dhO�G��� ��lJ��) ���V�M�Ej0����֌����z�&�%��9/G]H!���j���:A��V�*]�2ڦ����u"^j��s�B�z� j��<�	���J��|܆�nc��#~.�-W�d�ȝGO����W\�zh���޸��b��2�_�}=Ƌ����s -1��t0�w��"PTV�0șPC�_�4�� |=���x��j���~�R�І4�&$Vi��pS��SO��ϵI,���GZ��:��zo+����zl�m�;O,�ɉ�3�;L���Z*�AК��R��*��Y�^I�r����C���A�7�o�jEs��.!M�x��<���̢������cwI�;L�!?�����TVsx<��!w��K�A��$f�U�5�d����.�t�8.��[A�Oj�4�(���6G��?�L�����k�M7�hR(>���0��ghS(��_�g�$�=9`�f�u�E.������MvC��>� =Щם�L̔ER�j}W����m��M�������T�Ֆ����J���i�N����h��q)7���U�u�LZ��ۑhC�(�f ��~a����[�-E�`��ðc������� w�k�?r�Q��+X$r?%,�2j�N�~c����g��7x�@DE�k�3�3_�"ɦ�VhC,�n!�R�L�_z�O�|6��SP:�#��k�����}/��,|:FǍ9����Z����I��٠�*�x\�~�u��s����N�����'����?�����n�xQ�2%~��Z*���+�7%w~�7�r|[�-Z�kb��2�N[^RX�����Aq�E���e�� �]�ai�� �R�0�j�\�6s��_�~1��,]�5i�"~0��B�n�i�K��+9J�@F���<�{H�+�87�ϱ8C�U������5'zd��P��������R��v5�<���}|�?5��2��zo� �ߖSp�Ө�WsW��S�^"3�v���i
7������X�)ID��`۵g��^ �PW���Ey��$�?ۘl�Ȇ~���	�{��B&��ټ��N�EU�?�*=���:���-	�� �˾�F�����ׅN���p�S���D����lB��u8��R �E�F��Z�#gR|���EEG/9������.�ZcZ�V�`u�!Ki]L�9���F�a�&�~�p�v-f�0lW�W�a����;�d�*+����]��� ^���M�Ib�ǡ�N�a��0h� p
��L蠻~r�XS�˩�#Z]�_�SV�w��r����%'�S�9rx�������y�E���>�$0	�X���ˠ�t�$�?n�00�HlϋP�������#��=k[R�0C�i�	��N���QI�	�]���BRAZ��%z��M:!u�}�];��rw��c6�?v�9	
�`��a�iD	�D��t�v?�}^p5k�p�4ׅk��#���7�G9·�"���ժ�G[��m����S�!x��O�"�F�i�����������Lt�|�@w>pm��@�����8:*�=>��:qE�E|e�'��czP��*��},�\+K��vhap���d�8ę�����uݦ���C�X?	ҷ���-͎���X���?�����%G�E�·�s� "��܋ZnXa��&w���`6�g���tkED�8,ļ���K�/ �N�d�S�>�Ne��`�$�o�'o�+�68	l<����z����&������a�9������_`���>챲eK����1��)^:ު?�A����J��O��Y{�9��+�"9[�s"N�����hm�ґ]���,�mH�=ΠI^V��fS��s�����{���,��#�V���JI��5p��`��yq��VF>�`�d>�������k4��(V�T����~EaxI���J�M�� ��ΝhݨM}p4��e�Py�4pN?���b5M���/��o�"6e'/t-��Sm�(_`T��l?T���Qf,]�M\=����+��z��%�#v��S�ٚ�}g#����e�s�����0ON�M��}�䩙(��C�N]���/Z�ZF.F�P]X�s ��+�MO蔏�;�}tGqy���WDI�X�}n`�tŝ�xע���4����2+sʋo�����d�D�Vi��O�6����,y,��n�J��uc���Dw����n��i�˂M�<��(-V��]I)uұ��]:�ۧ�s���h�yFt���[��"�u�=mTm!�������J�Zw��3��}s�u�� ����z�."�u�/�HҦ�h�t��;�[�Z�v#��u�Rٮ��\���l�-��$�1�y<@`�x�We���[��dg4c:d���
��{��}�����$;����a7MQ�Z�BeIŬ�
L&�v](g��h�K䒚���p��0	$���.��������w��jb
d#�������ݓbb; se]�e��t��w��<�j�,��y4����Z������A�Pb~�x����qҐ�����@y��gʝ��~��&[qoN��g�\Dq!�J�>��q,��15��0K��z٩�Y���m�.�qĲ�C�s�&���а�g�m��΀n�{��|B�M5iI ��K��r�kq�hhu�4�	�Ry���/PP�8?N�QY>�=�U>p�H���drz�-G���6~��X"�i���U<�ܻO�xܫ��[��h�s�=a�8Vpu�3���N��nIQ��O@��cyeb�Nzg�gJ6�,
�)�T�5�Ϙ�}�kӢJϖމ�?����r��xBʌ5��̋���+��1$�<E�۹��R�li+zn���V/pz��6ya'W���#��WF�$k���(���n�"��5�����]� �C��s .}�~��%*��������\EB��]%�%Zϻ ;���Lڹv�t�	c�B��b������lJ�M�~�F7$$..t��g�~�սM8�V�6g�'��K��j5"}����|�����P�EQ������kj��9R��s�\w+�0*��E�?|D<<'O.G%�j��:G_�����/s����>zw}P�+ђ���k�$�d~Jvl_��<�0?���];Y���Y]{�.;��K%�v{B���-u������vw-[m��-�_�z�"�J�2��W�Un{*���6M���x��`X��Xj���1ً���3���?��<�����+1���U���+�<�2�b�?3�2ݧs۰ɀ�HR�xɯV�l6����E��r*�nޔ�k��<��v����&i|����)���É�T�����9x�S�;�b�v����765��7�,D�����UԞ�詡DY�qҚOw"����7U�}I����Z���#��nNHݐ3�w,�Y�q9x岏!8~��N��w��̙���tا�������dt��4�}P�m�+�z4�L��)������>�?Ҟ�����iY�ž�aAb�����|��]�C�8a����%��7Cu��4Z�Ҏ*����
�����FDG�SB��#㞪0G�d���@ ��h���|eۖp�I�(a��<�Q�� �A'�F��
�q���=��宫H����y'ּ���0>�c5�.�*�\!Рʾ��[�����NZ�s��f��5��ʮ���9�v��t;�٣��[_�I���gޔE/Y�!ώ���W5�Ӎd�_~\eܴ>ͬꡒ�N9{@�S���!Ļ`��(p��FLs��cj{���IV�I�����(<�`���GB.V�7x��{߭�T�uN7��`�
`e�c�pn�}����׈U .��%l�h����oSwA%&k'P6j���m��J�h�yM
{ӊ�K���\F�Ɠ0<�Mw���U,��]F-*o��6F#p��F�1>&S��K������4<.�����(�{�nwY�UJ���.���Ī�{��oR�����:~�W'�l���,HRUR�ƿ���5/��ŕi���QНe��ӣ�:�����|�0��p�Ir��l��ێ�U*x����[��4�?)K���<"aH�Ŀ�}��uEI��\���Zz2|�⶟������fѺ<�Fӝ���p�A��E�S�p�Y^G�rmwM�;�3�r
���.ͽ���e\�H����8&����P`��mi7���v��������a��� %��l0��yڠg��ı��x����"�qwq�ѝ�c�--_�,�w��g����T\���U�������D�Q� �	���=�-���i>�昈D'����Ck��O�.�O�F9'ʨq�Ї����g�C肣�O������HOm�&ͧ����D����۞u����7s�A%�����v&�w�����-I�~Թ͚��~�8��L�����\�YS���)9j1=�8.(>�B!�K9�����l��<�:�U2ʳf����K.�ޑ�4N>~!�ҙ�P�)egQï������H��mQC���2�:����%r�t�˭��=5��l�vK���x"g�6�O%\�Bnr~�rBx7W�զ�]b�K6C��˯kuŉ��#�M�<D�e�W$>�G����?��:� �;���4n�S\Wbk4xy�NjT�G��s�t��e떜���8[f$/���*�C�����B����|��
X-����:A>W���$
]�a�8�f�~/A^��SJ����⦽]#}��\�����~e~�y��3�Q��K+|C�+Q��8j�&RZ��p5���R��Bs�9.6����pХXR�w*�އ�G�J>��}��B�GV�ݙ����*�Q�Wʀ�5�	��Ms�d���=������x#0��JB�5[� R߲�*)^a&���u<[��b�[�{���S���|����S�D����I�"&��!��(�E@!	��rU�T��y����-M`�B���x{�,�`#��8vZn@��P#���ٴ���w�\�>iV�9������SSqw���p-��cZKF�Nf5��/l.��X}+��z ��s�O.�^.ߎ;10�ǖq$�J�l?�޻����]ӵ�m,��ӪM�2;��8�R�0>^��� �G��Th���_zh�?�˕��Dx)c�Xi�? �@R�|��eޝO�m��w�Y��o���z뭗|�*>������lʕ67@At�H88eV����7S �Z"�GT��
P�����o��ؤH�Tes's5soЀ 7z��5N�)wQn{1N�H�Eݟ�g� A���$]Ժ�W���?;"�YC>�<Ͻq5��P��1iҸ�AYUֶ]K	N�"�FY�/>o�ƛo�h�:v���>n�i@�S{�g��9�����,��y]��3/o�4�f���jrVU=Y��캍�p�K�BC�Xc�@`�E@�ief�N)K�l������oL�O��Ь�kӆ�1�U��^{�*o�!p��6�وnσ���V%�r�f��������
��"��g����}���[�Z�ps�!&��GAd��:��@/k�Eb./sw@�I�.�3���"����}ݢ^��-8p����C�a�/�'b&p���	ܧ[o�=��m޼��2L�9�&�'�g,	��ƻ�R������)�LC��,����՜��z��x�kժ��m�nܸ�|�>+~��#����a��i�����Z��W��h�}�IZ6$�T��3�6��;'����[m$��{�*�)�<��h0�sN)�z�H�M6��O"��)V��_H���ǿ���ɲ�
���k"C�hu]$���$7�;H�~sk�E�d֭�Θ���~��Q��ۤ]��s!���T�z"�R��D�V9f�f͚'�v�]�@��:Z�jc�G�GT�#�@�O��x]��5Z�\ok&
�z�W�����a�F4�����;����dE����V�4m�����d-i�q�%k������煻kf��ۯ���7���4X�_�2�  sL��~�mm �7mr����C��D���Jc� %�ܐL)�l�H��a?��O��& �`�HMR��y�$]��4�^���!4G���� 2_��iyPWy��݄�[�u��⹜���u�Q�����_�Ğ��%���n��9������}�q� ����B�{�������]����R��V"s,%yF��1c+%��!B&�Ʒ"�OD���Z3Bn�q��ceq�{���}���*�d�YA���:�	߬a־]�l��]o����uޥ���C����@ ����k�
pר���"�l��6��CO��J�&m�:��AJ	dG$�H4SX"7���r�q������}��^��=��c�Zt�����;��U��i�=�Uvs�GaCj.�b0���p�=�������u��y�K���h���"�ǵp��^|�%度w�ڋ����,��F3�ߤ$(q�S����{�5��3�!����K,�5�q(U���ov>�{��4��%葴DJ�N�C��������b��l��ꜷf���9sǄ�>s��Y��<��R��!B�T�U��ͳ5�X#友�V��*�$d���/��B�e�]�̶��!2��i ���"�A��N�馛���w�����gU�YwE�o-�^�ggE�χ�Fmt�t�eh"3�a�b8��r,sE{������!D4qƱ@������'kE3�F��A�q*Y�(���X @`p !c�׶��1����kp�>�ժ�k4':ޡ�7ѷM���k��aٷ�;���+��U{�[^H�,��> �Q�$��Kni��4�+���j��|�V*�k3����>=(�1��<��4��D��^!�jja
I�9Alΐ3DiB�"�����u��E��;�c�ï��Hy�"\�� }v�����'2�!4�?��%����C��4�^j�b��l>GG�pP�	���6�{^y
Y�z�'H�������B��	q���G��x퇟F��Z�f�.��Z�R�ܱN0p��B;g̟{�q8��xjʒRKo�dmy�>����x�ɽ�x�\3=��A�a.={v����dUIB��F�g���<}'�ӇS̓�W~�j�go��	m�70O��M�)�g�qF�kO�<�)>riމ!Dk�h�"���A�`����W^}��e�]�����8Y V���Cj&'�@ȵ��C��t+��I<UR�m���Iy���>\�� g�?�9�c�L���c�@�s�A�͛Ϛn���>$i��ѱc�� &`&̋sF��2,iǶ4����z�R�g�x'M��ܩ�|�]p�y_O���q���@��w��<@.�<����Fet��GYX\0�I��Z��.�7�����C�G �E@)i�p�!��:��c�M6�,��{���w�W�A�L��5x�u�l�=�R��ǳ;�K��%34z|����R�F�eW���?����o�����-��Qk���+O>���;��W�YH=�S�}�	�"W��w���?N޸���nyN���Y�겲4L��&'m�i��C�<s�q�;�˖�w������ڴ>�ĊAqu�է��� :[��)r!�a	�:ߑ�#<��>č��ƌ����oPV���k�}����_��&L�cF�r��f����w��(k0�	&�9���^i�	?�D�r��F���������@ 0�!�t��E G��vk��-��r�*�'Zpl�hې(9�T����M��H󔗎y�M>!.-�i�Is}��P}�%E������թ-��b2w�:̣�=i���wε#�!0>s�Y1�̩k.�[��K�N��v�R��	�9�6��s�Y/Z)�(�z`A�[�s�ȧ��S�p}�y=�Ƈ��}�b�-�Z���.G���`����J�W-��sKCC��J��O����w���i��t��0.�3s�����E%��7���<�{:�B�N��@`^A`���M��7�nw����RK-�4m�F;��K�:ks�!��U����T��w6j�@�̘�!B�͐-Ģͼ�L��Kk��pS�GqĚ���\�a*r�t�j�B(\�mK]~Brp$g���L�ώֈ���{�ɾw��D�qNK3�ƻ���x�aL�2�t��]u����oij@]M1�^�iR �/�9Z2�����2`N.��1�[�%0J5Ζ�?C]�$L�� w�Å�L(z=�ۙz\���`��`9	�%�9��?���>'ޕ�S POx��P����t�I'��2��w�}�<�f���l�h[��3�<�ʷ�YC�h����Zj�ϝ"%�N$tV�~�=5�eHck�6�}��?q�5��!�B�{�V(c҂݇�9�� q�Y�u���u̾���W��[�v��y�N7�������O>3Q�v�Ikw@s0��݌h蜗�eO�L�}�]��&�3�Ҭ�c�&>!��YD�����<ET�����M%u����<eE,���E�c����I��3ں��~+����V;cDP܌�Gs-J��#=Mļ�W4P�M35�HĀ�eR�8 ���)C_s��4��!u�����5m��������.P��?��=����ȧ�"�;�	2�����rM8oNb߼����5�R��g�7>梦�xk�ˤ^�k{�0a�hF�x&`J͂�ڪUPh��״%���:,��:�"d��.��b��Yϼc]^b�X��v�}��&��5w�3�   ̩zk��]Y�cz~�"�=T��$�X��?L��{~Od2��h���qŔ"��S����y�19���/!�  2�u��_+R_ޕ�~���%�0>p46���(!Y��	t���FM6j>�_
i�4��D(�D��h̙EH���>2����۾(���C��幞���� 3
?uk����s��!;H҂̬���x-V�+^�	o����?5/�k������k[K/yq,[�6�0����+'��9��1�5��N�c�D���=B�
0b<��Q#�٧z��>$��v��C��y9p�1�b`Mx���=AH��k�>?�g/�"��|qr 0�#��SO�T���J�Z��J��Β�mBw.6� DH-��o�={饗�cBeG#sZR�߶�k��fY ��i�S�C9�w��"���#�����퓆�,,�Ո��9װٛsXsd}���$V��mn7�ɵ������9ޟ#֋� :2����1-�}�"YNT��^��Fqiּ��>}���4�y������� �$�� G��S����|�"�u�x��!�-�bA�'�5�����L��4/~c����68r���4g�0L�s�����m������W/�r�)���n�֓��*aK��ӦO�:%_!�>�@�]פ�A(|FМ��AK���?�TU�^qŕWx��O��ʫ�oԨ�;��K�ڿ̵!/b�yzj;ϩi\ Q^3y�'8�f�A��x7eq?o���'�)�@������w��Ұ�H��M�E� �u��g�6.r!Pi��O�@K��W�C `L���yT�C3g�h��w�Aʚk����������R�����~�"1~@�\��22ɧ�Λ����u���ʎ�E?�8�gB�Y��@`�E`�ͷ�������[nӦ>J�N[�ЯP�Rg囿#�pY֡c��A���#�v�-���/����dmڶ��,�'����d"��s��	J���j��|܋/��A���h�=�O���\r6�v��L���x�)�t�<�\q�͵۩�Y4[��x�X����6㻻D�| �"qKDHR��A�y�7ך2%/�:yr^>��&o��������)X�z����M c��#d4JZ6k꼒gO�<���k�$�|�i��F1��g-�յ�Y?և��s4u��tD+G��� ״is�el�sϽ��N���K�o�V<��R纥6�x��_~9�Ԟ_y�!1͚5�Z&fk���~'o�}�KI�R��g��_�ޚ�s���_�A��=��������H|���+m��HM�M�k׮u6����� "��|�-"�ϴ�7�蹀�z�s�q��w픰�Rd��d�|�F][4G�w�̋�a�����i='ة�Ɋڰs�9�Z��퐛����8���pm��5霴��}|��M���1�m�g�$'�ɵ�� 9��_���u=v��{��j}`G�����)ڵ+�9����f4)��C���!q>#��� Z~:���B���?�ȣ�;��=�r�[���)���#�� <a.���<	�|����5qw`�ܮu����Orٌ��y�_��"��s!m�'�o߱��vXҲ!̦�N;w����B2gC8�D��W[m�쭷�U��OA�!�kށ,�9@N<�w[���,X����	�H����"��~Z>g����&��}�iB�h�n�Z��xcM&�q����\�p�=�h����9߾{��b�2�Q���=b�$o��X�ݾt� C���r�y �q/�����:�̑5!<踵�������|�v<@Ŀ�R	;s�	��Y��	��J�+���ﾛ��s��%L�pq�W\��<�_l�\��ށs��bR�@ 0�H�n��nw�(6{���v�ɁI�,)�f������=��s&U��+�fؠ!t6uþhH�>��RJ����! k�&?�����bZ�����i���/�"���4I_׹ю���l����Sʊ9��Htk�*��q	�����ͅ0e��þ|�U[$Jwj��![���2��Ʊ�P��w0u�-���O���.r�s`����<�sGP`͌�{ŵ��@�ʫu���<��i������p����θh�|ƃ15�D�N���j_U���6�3����$ �������2��)-���S{�����ڟ|�Gg��{o��f�f�W��DBD�Wʟ�$H�Z�&j�C�����T�WQ�v����Ŋk��xg�}_mb��n���6ǚP,�'BI�+Ͽ7A��7���6�5��\>��ڞ���V����G��%_@�=�\��O1.�]��#0���ꫧ�6��q; �u�8�C�������y�"���=���2?�l��Xxc�v�������y��[o=$�|��-A��Z P�(�h�s�=�xi�-��g��LZ9Z�X�(��*-O���g�%O�j͛�̶�v�������3����m2�&��ݚ�	�h����g��-��;w�[�o^��]�S�a�S��v��#ާL��,@��=w��q�M�|���RD@�� M�xH�)e�c�麩�BgNX�r�����3���%l��fh��
������tL���U���Q�>u��̋�st?{�b�<��K��1篿P�n Ɩ��U"�m������z����B�̀����BࡇZ�C9[���9Z��f�L�3Z��A�� ��,Z=f`6t�-�;��U��&຦u�̋����_4���>����o�G���>ǂA1G�1d������AtT���I��_��s���Gk7k��	�0��7GA��B����lp��ь���=��5���fo�s�{��rA�Z6��h���e.������ u��Ksc޸�B(����j���}p}��cܟF =~��<����_���|��c)4or��ԅ��8��Z��)�k��&y�ԂgcF�*�zg�����*��ح��Z"sJ�����g����Ec�y��L���Zyќ�S�^$u�-�i�K�z"x�1x�\ E�@�iҤq:�&{�ܽNL��%(J�j.�
�N���9o�f%��G���9qOЄ!\��#\9��mڶϜ�9ps?� ~q�ʸ��3s�YD��c�|���5�~���}�$�����yX8!��Ǝ���>�|��w���k������%DP�\y�bҁ�T{�������+���IaҖ�i������X�$�	3�g���߫���\�qQ���j2S�Mn���;@�Q�Y��u�i��]�v�U+��xM���W�ċ&x ���w���iU���x~Ϲ��I����yz�^�>r��)%�yՔ*��O��:ϔ4O����ghĐ �dh�<$������s��Z.����-�p<�s����X����&~����i�Ɖx��g.������o�!,������q�q>ǭc��G��]w�u�n�a�۰���Y�@���2F
f;��^G���Y�M�V42�����)��Ax���>���Ak;tIս���(VU3�ҲX`1Bgs7��ъ��l��y��H���{ܢp�6��F�M���8��Y�G��QNܼā~��(�W��/��F;�1��nB��"X���>0/�����Ƈ�CG�r^�Ф&�!���;ײU��Q��sѰ}�ꫯ�H�Ný��\��k��X(����ܦ��9�����=��s�+����l��/��?�@`.E@�n�7�t�K��L�3Z9�斡hf-[6OAnj���S/6d�ֆvIA��_��|���-K)�D�9�ł*֦s��5PS��9I�5���\;.�-dc����;ư��g�8V$t��
�`Ʊ`�9�H�UU����`�<�=o<b!����1oS�1�x�Ղ=xzm�z.X4��p}�y��ٮ]��Y��ك�{�;��>n��$�@���X vỸu���|{�(��g�_p.sf��=�w2QV�7��������f.�o4OM;4�y�v�b~+�z[3�Ǿr��![�Z+�H5��F�CmLSmv���vZ�4!#Ȝ���Ie�2�1��`r�5c��AR�J=���<�����&��Z߯��s�ټ^��[c6I{<W���B�_�w.��c�[o��BDN�yZ������ArW@�h�N��1yC�vp��a|4�ƍ����{������qm�:Ǡ5#��[�p���>g�"�1\.ŠA����7�83 S��wn�̋D��st���+j���QG5���nN_gh�s���uP@[c��u2�o����Ϫf�o�rcS�;"��A�͚�y�ӧO�,IisN���ba��FSˢ����'?yA�69Z�q��}�E|]�.j�����7N3I;��d]�|mN�`�ql�7�9-����z��F�[P��r-_�ti����@��ՠ8W[k ���Fg��s�}��i|��1�s�	�`<�����d��}wV������Ʋ�BwP�r��X
�͗,�%^y�������t�A 4�9�^�L��E@�CK#�F��F��;�i�.id�bm�uQ����['EB;���0��g�en)u�H�cl��i0U;5a�ti"�kR�_�&Ydg�0i��=��&����LD֖��c�.�M�}�%�����̂���s��Ú������3�kbGC7>jQ��-����^�;�h1};�=σ���\���BL��7�a���[�q~�3�(X#w�����7�H��ZQ��K��g�q�lG 4��y\0�9������f�;W�f�m:��?����f��n-Ӥ�cD�/$������_3�+���Mۚh2�gDZ�ᶠ6W'M�drwʓ��z�Fm��I��MKK/�h�����yֺ
�n���/v�Z�Tρp"���W,��}�`ia��g�p�����?��%��*n�o���6�����	�#p�c���D��+�g~.L��d�Y��e���y0g^.#���"��v_�FL�E_Bd���Z���	p������F ������@��/n�ni�5����V`�ujm�9[���3{ꩧ�Cj���w�}�f�f�������h�-[��:��EV�H�<9$�ʔ��#���K�Ӭi�YW3.j���C�`���y1M�n�Y���;E���j]����`7�����\��5������v	pݼ���D�.c�Hn^����=*c;��qvqp���
1 <8��q�C(����0����}�9 Nߏ���h���w�G3�s�Sfar�M@�.��/4�?��6�r�hch��&0j�h�ͣ���.��*�,��$>����j4�� mr�N֦4I�4V�	�O�&Z�ͨF&��]�NQa����<�8��û�������v�)���U�'r�r�UWWJ�ڌ7i���'o�������C :'{��RDn����b*y�/"��]�ʑ�u���S/t�?�H��6`�q�D]����J���1��֋�_����Au� 6�x<|�o/�ȭ��3�W��d�(�{5y��yl�Ӧv��Ns΅@�7�z��s�^�Q�5!|�ދq
\;��g���q�&[1��.k����:�+��zu�\��a���yfYA��̭�=Qi��"��2���_��|n�e�]X�DO��o�MA�}�*m.�ڨ5lX�Te��Ⱥ)���>o����~X�b��5:mPUڴ+���ӟ����9S��M��D='蔉:~����?W9́"�!�����1�{
O�3�0{���W���2��Yc�5�1��Zzu��#iM��Ȝ�&�'�T�>g&r_�;����N]�"���-́T&-k�U%��T��Z?3+��;��VZ$�"I�X�Zr]�z�- ����n�4c:Z�d���y���3�L��h����k,j�E!�s/Ω.�����}�-�x�<8��s!m㗏�w�������I�de)�ܹ-����_ֈR� k�s��/��b��/��U�.�5���@�}{~��)����~�Z��3�<��6���0zhØ"m��6��"�
"����
�_��K���yS,n�^&�����Em�Ǣ�X3����C<E�i��3Q�	����� 'H�h�\��:o�H�mi�-�Ԓߨ��x�	���k��9��f�mvS�����f�
R"��c�NɄ��g�kM�+'���� Z[���f�����VF�op�d�SҰ�`j%�MЦV6}�ZMI�-i���hO&�R�������Y�̤T���}�t�Zo�����t��ɿ��/γH�Ӻ���k����8v]���8ߗH2���RX�X8��8X8��-ا��'%��5l�����f���I�+�,�7�^rL�od�~o���]��EJ��7�����E7�>�*.i�Q
L���_)�uCm8�5jԤ��V:���ڍ�EM��B�	ȗM3��?i޸��x#�f�@����yCo�^#�{��f��O� =Fݼc@9�A���ֈ����(L�g��Z?S�����?P��E�O��2v饗����q��7/��?��f�yH��>���c��EPƏ� �Uڑ�d%a3ǜn��Q�9�V��&�c�2��r�(w�����W��tO���Ԋ�����-OK����I�^Ԁ��A\�Q��n�C���%s�i���<�b��e[0�{��ֿq��
q����zP��� :Ux��~��wxu�������=����3]����"\n�����`_;�ڷ/��*�������~��<��q�Y�@�, qnB�\q�]wuy�G�ʄ��6�62�v���v�UW-�n4�5ebO�=6A���0�L�jѼX�?�AC/jn|W�d�ffM������xoRE����޴-L0���/u�¬?LD7^��h��3a�4�w�;D��o��&y��zz�zꩋ)g�J�Ҳ��4�|G����m�'틵w�<���k�\U�uq,�A���}�E��5=ƵU�,UD�Z���6)�C7i�
�1��޿�������5d��؎�F���������\����#����o���Mh�V}|�߱��&m0�7�7[�Xh,�.Ƴ�c#�<���������l��A��M����k�3�7�y!�☣M�\J�8��*}��~������L������t�J=�ם#�B�#n�웄v4Rg�.z��p+m�]Ux��b�-�X���F	��q#�+��9�g+���D;��{�nX��?��$_�!2�52��������&IkE����󔣼ʙ�>� �{2k�+k��l��yРo&�����YN�X?��O�Z�����A�V�J��+��i�?�~w��gߣ��=W[m�Fh����F
AMS&W'�47��z�6m�I�A��U��Ҭݛ���܁US-'yn�5����D��e�4mҝ�@f�/Z\|\]�������+&<�a�{���/���٪`��\�fL��^׍g<g�gư��jp|fa�����2�5��fqά�ߡ��VO�,0X\T-P�=!����`3}�\2.k�K�F���S*S{����믿~��g�V\/W
B�X�A�m���v�s���ZZ\gul�!�hL�ir���c�f�y�� ��,�%�+6���My���x�iכ>Ģ��q��ͯ΃�5��$]4�����ps�H��P�.оc���>�tk^�5�㯟�9�ӆ9R�W�����f����_�<Fḱ+�����cW
�]o�[{��!צ�)�lc	Y���ߩw�ީ8�ii���Ŀ�fP�GM�AnM�6S��ŕ:� �@8����æe�xMu-+EB�`�p(�}�&+�I�����|�Lv�U��&\k�|_7��(x�Jc�˥z�E+�-^sQ���c�JMK��	� ������>�}3���%^-[���ieNcݮ��u�q*s�8��w@�^[j-'�1q��Y�,�o��U.�B�v�Vdޱ&s=A�s�-������Kʬ~���/����e2.��O.2U�����fP��pmWW��[Qk�%؊�l*��Uz�Mn2o �.�UU�n�"A��
��sҮL �Gmx�8=j?���q�����ڞ?��)2Os�5��X���������������שЊR��R�e:���+r�T_K�����*7Y��?H�#$�k�n�`�X�ey�UW=����{�=�����mps��S��{����4��M�v�~��n�6��[o�%"b^gn�	��ۼ�g��E��B���ZSu����t���C/ܿ�c�ԋV�/ZbLr����s�S<���u����L�8���y�sl��5Fu#���?�"�"�R���<<k��q�,`G0��omږ����x%��kX�p��W|g���)s�7��9L8�/w�eGqD����*���1� �>��ʩQ]�����}�-�W@[���&�����A�u{C�\Dě=���a�Yx��5>��VM�ұS�9��Iz?F����d�9D����U�x|����瘱a�I��W68V�S�#U� խ��n�c��vz�Q�]�iv����w=�����H��25O���Y���1]s�5Y�;}Ǵ�0�������q�񃡻�����w�ɶ�n�L���;�s�4�������'��:v��˿���էdcƎS�����;�������o����K�4��'�ɵ�I���%J�l��L&�b$���Մ�9�D��m�6Ys=O�m�|����E뀉ʚzn%)�5�#���㍹����Z;����iA�W��-Lx]r�[3� �1;�1&t��=�p���:��&}լ��N���>�B@H�t6�G؏�y_*3Jk�N�ݮR�����<��ŒJ��C?m������WĽ�z��I�^#z(S`2'��_����9��M�;�ե�3�&����Ňz~�(Z���8#�1Qf�4���ϴ/��n�^{��P�V�T*��5U�|2?��<[k3�_�n�̺��Ict�Ukm�y5՚�	�������U��dr��� 7g�fz�x�]Q�s�->s-n	Xٱ��y��ƿ���s�dx���S�V"��~�tѲ��D
����k��a��H�����^���l��W�\-�X �HƘ�k����$Z���`kͼ�tn̋�m��)vEs�T�K>?�瘠�.ƳP��ob R,2�p9��e_�ߔ%�+
x.��r�u��1u�;��&�'*>���s_:�����
�h�]vy夓N���1�#�>��{ｷ��'���H{[�!w����`���ɯ��_�v�i?3d�&�Y�����FVU�@����}��>�MbR�~���S���K��`J�>���0�M�����G��f�]sǑ�Q���3��$"�I� :�)>�h���ܾu����\���!̥�����?f��k�M6Ʊ���.iN��H�c���ٳW
�i����!'(*��,�nI�.���l-�k(j�&��X&W�m]�e�ZGK!��H��Ҿ��nӻ��㋿��<�U\���q��|O}]��5�j<,���,[hh�Y�#ȼ.���^[h��P��]��..�[+�,<��f�kf\k��J뭒��>��?� ����{�����ԍ���^�ή!E��~��|��v�_��g��P��T�[��i3�0c"��e.�>���3m
oh�xTD�_]#T�d�	�Q~m������TtkE�/(͹��YRk^T�=�Kg�z�Z��Y�u@�b�����f^�4�@�V��n�e2�'���)P1�#���W�M��)����$A����O9�{ s�b+����\4�[S�6W�
7#��@���1>� Q�Eµل[H�u�~��z\S��}c\��s����o��5s�G>w�P���:f��r�X:�����uj��r]��=O�Ӗn���!V�ƳPY�=�b��k,�%ޯL�{:�/v�i���k���Y��Y�c�f��/����?����eV��wL�%��nug�2��l��sk$l"l
%�҆5B�O�)�[χD2߬���#}��_���t-�:��3�?��s�T߼��ً�RK��[��҆9�0m��fgS+��7j����f�F�|e��3��r���Δa�ʳ����V�@�D����SU7��i���O�<�"B4�Y��%�i��M�?�I�����M���H�&���ݚsQ������횠�kʶ�p?lw��'��E���� 4w7��9����4t�g��b�5cX�10&E�V	��\YB�c��I��z6J���1^� ��O�0����0��>��)�SѴ姝v�6W_}��JkZ��k�9�.H� ��FA��}�l0l�lld�t~����Qm7i�a2M���`��S=묳Z�kY;E��PJ؊�{Qm���ݵ�/�������9��s��1e�0Ȏ>��dj����OҴI;�ȝNz�[��R��Z$5�˹�r��+j��x ��\�UԮM(�l^��g���H=�S)@�c�5�{�"�	�x-����	�����㹆?g<������b+b����%ę���tq"σ��)�y��q���rqA��BO�JQ����S���k��ע5����V,�=l��s*�3P�a���@��@�\�S���+�>����f���h���4�w����ll�6�1��"���p�����9-�/6�_p��J����;)�`9mҽ�kkH>z	K��>,����L��l{�wd:'��AҮ��$l��C�1B��s��S�-�'��m"�sW��`�r��i�-�u����ϭ�z&ˢ�^���=�Hf6'	�v�Rq�c���v�X7 ��bQ�t��#8�)�p2; k��|nI ��	D��l"罣����f��?��p׷�d��H��"���z��u���Q�xQ��Z~��*�u�2�'��������wX&���s�A��>H% ��huL��y�I�ٰ�9���neڰh�w��[E������ӓi����t��{w݋��q7�G� �t��&IDM�r��Vp�Zf
4L�<��B�ý�0��琔	���J�����߻�U����n�K�&��c�Lo7Nc�ɂ��XW���+�����[�w5Zϧx��w��b�b�u�9@��P���'�|RK��h�:k�c5}G��������j�$�ap�M�?E����.�C�z�Ip����
	=���O�Zk���=������[@���z���ͣ��>��>��s�6�udbk��+ol
h���L��������g7�٭j����@_r�����[�6�T{�Y����k�W	�j`1�Z�#�l�p��g�̍7�t�O>ف"0h�r����<�01c�����?��k��%Fk��'���eSw�:&���X��[��f]$�n&^�q��x���A��3'p#�n��M�,��B��kS4��͘��s�9D�u�hX��7���{� C����������jX�@H�Z'�p�'�uSp��b��E�|o��^+�7�����{��'D���f��{�Gt7���2."�>������l���Z�Z���fCGV�Q8pF��xm����.	�V��3�9��Xoc�Q.7DCiQ��W+��U�6������W�}c��T�[�'�N�7�3�z���@���N�L5�Z�P��6�!�m�]�hq�D�7׹Uz�T.�
YR�x�as���X{Ě9)� ��|�駓��>_�/j��~/p"�<C���\W#4I#��fx��M:%�o-A�L\��mZ����K� ��t��M�+��>4c�a\k���©k�s��8[����-�'Lތ��n��Sz�>�E���"�����@����g<����o�\~+*hXO����@sxV֘��2\��G�����f	A��Y7�6�
�:Af�}D�j.�袴�9����a����hÙ�g���m��ɜ;Oj�7�pC�x��̨�ɷ�)�����6ʞ"��������Rߵ��b>�P�h3G�j�RMZbS�,�b@��s��~Sk��\V��;U�-��b!u�'�HMQ�<�!	���ONy]���BT����YG���[��9`�Dg30���ɔ�u�ċ�&J���6���)��?��n-���_}!��H��l���m~��L����v)0�+�ٴ��b`c���3�Gxo-��r�#�=���.0w~�H�\�ȃ-�s�Yk��TA��YL����м�볷�ä��>���G̺�"F
�?A�sЯBZ�*z�6��U�)�u�&OZ�M�L�������D��3O�u�ߐ�쭴��d��#m����K�Aco�bE�W)ڷ1d�cS9��h�r3dW\qE��㯶obN]�JLl��c�^Ӵi^� ��F`�)pQ[k�Ǻ�*�d�sU�LsMsAke,΁艁����u����xMPn"��Z���nr3����:Ǚ��eӾ�����nd<��W�WI0�fj�8�X�J| ڴ{��>(^����;�[&XWI�M�%��x,�/r$���x}���:�s��O�2��+�ԫ5�X�C3\Z_i��蜗�;��{�������b��b<�ي@�l���/&ZB���f�$ͼ ��T�9�Ȧb-F�h�;�H��>�,c��q�-��Ti��Ҽ'�{ei��D^kӝ_nk��)>h6\J�Z#�1���1C����8����м�ا35�մm�`�os*����<����.��wl�,]C�M�U�F@���C@J���W@������S�{�إk���y�p��W�s��9+�sz������>ǵC�m�lH蕪L؟s׿ Ŋp�G߻{Mq�e<N:k��;�h�ӝ���,E�m�B�:d���;��/^*�p�7��:�>���r7Q���7�?���n�*�Ts
V��rdBz��'��>��t�@����a���V��,�0�<��\�ȗ=�����(����vt2���[X���M�e�3�����j��Sg�T�ej��b�t2]dWX �W�0�E� ����+��TGku�G����l��-󏿜T&#��2JF�,�+��C��W�o~`��+��?�َ�bg:6h�nb�)�B�uӧv#m���}[���|๨�>:S1Y���hN>�9.ʺr.���p
��1�%�( ��M�eK^=�{� ��
�R�U �fꉩ�~���Ifo�_H��J�WU� 0�z�(��)zڀ2��ƣ���GF��Z�M�ߦo���>`���!���y{��I�r���q}��{����[,F��W�(7Dռ!��B��7�W 12�gPo�M١tGXx���4��(��G>Q����T����ۆ����"M��R%�^a!w�AQ:��sMG������K�꿜�\g��d\\�y/N�\j�����@ q�"��J�DK���Ѯ`1�'�.�F��ir�t�R�,K��{rG�ᙞ�\�Q���O靇���F~O���׼I!��i|����_x�ޤ\�x��ï����H��l�M���P������r��,Y�ۯގ�h��(��:��~mn,�C�6U� ����/n{�(�����[�*����]S��>��q����s.��S�<�"���)o�D>�GsBQS7Kz��ặQ��u�dCPe�_��G}F�#��	�_W��@E��%|�	�Xg�QE�o���]3*�3�}��ח]2}܍�T���&ʘ��K@,7<���������.f�b�e�9�.�@�a�n!�H��"��큘h�̄� �:�K}6`�c�)��G��)Z�H��H��7��D8����pvDdb(zS�s�Q�cQ���E{'n��T�U�ɾ�Ǖ4x�Ml]F�;A�kOO]��֍�����-֤��G	�P�'�C��H���s7��S�c�����g�������ോ���xm)J�#Y���L��(!H{e��.��>�����;���:E�D�{�����gʯ�N2�)\Y�-$q���/0r���*\b���l2��ۘ��q��Co�W&����L.��I�Mg���T�W��O��D0�V�3ḐV�C{��ӈ�А/Z���s�*�]��U1��q�����b֑F���L�z���GZ�����6G]/��}����Ҫ�R����B��i�=�_�5���ҹ{����k��W��h�8xh+�[�p�5���u�����\�l���`uD��O*����'Mr����$\CX�`pl��~<.���f�ᔁ��=��'�=�m�A�-u�M�����k#�yݫ����N�˸��@�Ee'����'�7E�(�|�? ;N�f�Hסu����_����O"�ֽ�J��73H Z����,;l��í$fvG�Ԟ���?�i���#�3��^��H����*t���A)�|x�g��U6�>� 0ҘD&E�wq�Yٷf���g��}hU���D��yO](.�^g�Y
����tV��0Ft��ﭡvM����0|k�y���:�A�� �S��/Y�=Ѳ�f��w�o��5rOD�t�f�F7,Jۈ����ح�[�пʾ�WF�x��q^�d����̞mo�M���mV	�\�Fz4��֟���^4���l0kp�Py�	��?g�T9Tf���h���֯�#ݘ8�p�r�A�JRk4�urb~?=�ή�Q�n��?S��}n��������������v�G����ʾ����h�Υ��:W�>���=����a��]�;|^_�͡>'-zd��o�ZB{?��4��ŸY�ͤ���q�^��$�%K��z�Ă��w�b�R��r�ݜ���f{��ؼ�t4�4ML�l��2l���R6��U�@p�#����Y���X��Sm�-
'����������\|�T�?��$EYKu�\9r�Q�-��K$��u�z�{7��Oh\2��\x&|�h6�S��<C������=�jO,�� ��+:R��}��
u��7�y����"�?����� 9�-Z�5?"��=�Pb��0�8����������xQX*��tg�x����)x�8����t�-����CPI($��8\�ͽ������Xy��~<�M
�����U����.�\<�*��+�4}���m�[T�{�[��/���8'4�֔�*߻+:?_q��=��J���ոY��t�R���<��F��)VOX ���
�ԎlX�U�,1���BI�4������h��֬o��M3�n����U(t1�N�v��XMA,�����K����>�U�5��Mj�Z爫��`T������̒B\�E�C����#3�T�p�	�W�)	��mc���
�ބ�\�x6PNָJ�{������C-'��x�c[C;�GH�6�ߞ�m��b䮸�`S�#3�lU2	:�6{5
�㪐�Y��͸'�/?�۞������U��P��x�l1a4f���uZ8?���x"�:uM}..�mo���'�	��H�37�������Fѥ
�fwj)'#��4�쪿�B��>.w
,zdAG��ײ��f�������0��!gyEg�';`�e��3O]�Hge�w����]0횏�Ye�@OZ�=\e}6��$nd��O�'���c*��ղC��PE�̅�m�hwr�����w��R-����ꍿ�B��.A�~YH9�W3ۗc�Q�
]_|}�ihY�����Uv52*��]�I�]�"_I�z/�;]7��k���=V邘�*W��ڑ�^^�z�&5�#��w��n˲#�6��5h�5��K9A$�3�����gѵf?(~��ȂHNPgo���P�L�U��������S*j�b�8)�'�������2���Xik:-�!��b�a
oyx��?��CA�Ža�Z��1%��g`���8ID-���>�=�C4��ؔ��5�	=�z�{�Q�w�������R��b\����;������)_}��Ξ�|<m�-���X�M��R�y�ޅ�E�����"a��a�j��t���o5���T�蘚�Բ����#��_�6E'z�
������B;���'@tֱ��y��En�h�w�9��G`ⷓ"�ۊ��r���q�fj�9aP�lxކZ�_O2ؙԡ�}�@��2Т#��h8�h�Kt?r쩕����f����N�l�̕�8Ͻ�s守���d�^�L2d��x�ܑ��̥�ݩ�s��'I����# vh-�����ߔn�)tbrқ'��R�?��_I���{v�]�x���Zc���yw��xY�n�bQ^�d]<[��u����J��'A�CJ�����tJ��'�y5��6�Ȟ�ɫm��;U�+D���%V�m�̮��Mǝ�Bij���l�xԃ������Ld��o�RU��h����u�ں�f5궃��3]�a��Q�#�^����s֟�kY���HY/���^y��؂`v�s�&�Ðۙ� �J��� tiL�Ki*W�������Ԇ�g� l�S�t .,N��_���ː�PT�P�f*��O�+�㈨Q��/��E�4��-,�̓$S�z��6zc��G�p"�'�S�A����bp[a�R{~P�������W6#�/8�P׽=�e���D%����5��XE�~�7�Z��q�xm��	�N�+����;�D�X*��<ý�fI�Y�8j�,)�'?�	�umX#ӕ�\,��_gPp������ls[�|b�%	����8pB��<m��6�pg{��� �{�t!���*��^y�>���JAۧ�8��&
u��ik��[��n!D�/E��oR��oF�R��;�7�F�7%�!���k�)��:�n6W6-h���eS�񜝮G�"|��{�"���aפ!Lf����`y���1uB���%���
Qv~5�놂�a��0ت��t�m��nit+҆m$�>
D��k���������(���u9uy��"���+@*B/��l���@�@���T~Ȩ�2��W%�h�FR��|�Ă�B����~��Nd���n��\6���DCLZ���Z؜}M�|�^u�T����w��I�T�LƅQ�8��n�kfQ�T��s�Usg\�;�,O��;i~=�oH�XNl�~`�=�Ca�	����K�	�R���(�A*�,�=[a�/��1�%)���^�ٯ��&�ŕ�L}+���rfr$�dBl��ȅ��l-����|���#y�#�aa�@@���e|��V�G���W���(��V�FD��ĨfZ�+�/v�[�����h��iE�̮��TP�UF�\�j���s�6'� E�_a���R�G ��/$����nK+�uҬ�ѵ�v���y�Uȓ��D���JR)��d��,�sU�w�!��T�4�ktf��/�����GjB����9�6.��O��&U���y��DH��T�yk�fs>��{��'���>�����1� �p
R��//�_�����m*'�@ ��N��ė5�{2N�����t٫�ӝS	MA���Vr�#tԂ1'����q?3��mybҪʘ����x�8?�')T��
)��cu5�� ��B�$gƑ����H�M��?��ȷ�+z"�
���I��z�u��;�1?�@�=���j�d���'?QG;u��nX&:u��%S��a���J����3V,�~��x'�������hO�2r�[}u+Y	H8���9��{qkE�g�H䘌���K^�Ȏeݴ����j�������ߌ$���5����!���c�)Y��з�:�r��0���H���R-Zx)kh������B��i����NS��jqӰ�@����:��l�sQ�4��Q�;E#őȟ),v����ln7c�˻.:v�>�V6�����A>-TL��Nx<���FN�H#7}=�t1�$JB���[X'�M���6ٝ��Z_���ac��\��nl[q��d�^� �nܓA>�2�o���M����� ζb���ހVGn�N��4T�O��P5���4p*�/�{|S�[S�3��~��_�#<cQm]��޿�b���i|����x��8�&3���o���+�qG�/ AsS;�_��ԋN�Z���$M)D#�
I�@x��ʂ��ܬݨ�������Q 2XL�	��=���ОJ�I[�W_�"�w2��狡�Wu!ԉ�} ����T�>���ᒓ����:Z�b��&�>��Z��g5�4�EC��錱�U�[>$�9�P� �����֍���b��yP0��y�a��ۜ@��b}��r/������<��{H��+�m��"J��ئ�V:��������,���b�� ���*T
�4��4�M���o�"�Y���R��7kp�70r�H�y g�W�|��d��h3o8&�ZyپYV,�
�	/�R⛲ ��II*�f4�J���ء�[��刧�F���נ�y�7g�v��x3�[͵�L\5��aӅ�p����n";O�:�)=J[ 0��=����^|=H	���Ю��:��V��?2��m��i��J�,��O`�b!��uT���NTT��U���C0�����?���Ec���V�?(8�j?-����n�V�MS���i�M�mH:2���m�Kٔ�o9@�s��	ȟ����c�87�M@:�A�W�cX�c�����Z���ݐ�7å'�����(v�#�a�VU@��ęEg�x�����a�<���쵯]��������2!GF�e��͔J���Ql�m��{�����Q��V|�epNhk�e�����|���Č���z��C����%�
v���V�2G��3F���;h3�!��zD�f�$E��)؋pȔ���K��{*�uD�_[+M��,2�@1iUj�i̗7VR]����G���zZ��y�k?��wC�<�^xW��]�/th�|��7>*�{�TWϼ�"J�<� �a�M�"h�.�S�O���v�U��>����}&̗:s2��b�}^��MS�Cҿ�V�)뿒��0��.�1�V~%<.��)PJ��h(1ڿ!� }8��HTQ)�3k#���F�ɥh��
����x� }���C"��4WM���4J��;ȷ~g����O!��oyf�乇\O�4� 8²k汷m��Y�;%�ċe�Ș_D���"Emo��,��r��Ya$Lo=�e�wz�/�;S�3����J��f��K�J�_��[��h���T���y�Obc�����%f<~����y�<&��y�5%��	��7�N�17o��]�=��J%H��;���5�����V���&e���V����[����oc�o�Ћ��}]S����=���/��[�=��%XM�4TmЧ�閎!�� ދ�U\�K��8���Y��n~x7X��գ#�B�)�e5�W��=�>�|Ԣ�]jA����>�`+7��Ȭ@oF�$ÆH���օ��j����[cӢ! �=PAl2:pj�ͩ�p�+����h�e��~�����'JS5
��f�6�:��*�U�h��Zv�[����Aժ��3�����ˆ���=��'�P�lf?˔|i��r�$���"f��bi���c��"��X�8���f&U]��ϩoT��p� �������曷�68���n9�eCĮk3�n3��O�T�zu��i5m���du�n�$Y��!��gd�>��Z_Hz1w'�my33`���
�P Ѫ�^�C¦%��m>�I�����*t<"��,i��*��Ԏ5ӷ��������T�2�h���p��K'N�g�0��L<.�}���ͰC
9��Ho�LC<���p��n�Ig;/�O�p)�#1���6�t=��=�69�H�|��۰�,�Sӎ]�2}��֔�.����h�8��m=��4�1�����	��h>d�����j[m�v�J��G.�Ȝ&t$��Wp���u���k���h�zP=��6��'4�
�#��.dT��AV%�c�d��Qj��{H�~��t�zC�&t5�(#�A�7Qƥ�ȩ�jB"H����p�-��j�����v%�x>3J����|q�l���l�J�_��
�"�&�a�u�Ih�b7���p�R5D-|	K���*����L���+����zp�t�R%%"5�]��JqEt�Qe��@�v4�����lJ*���\��
#e]n]���}�iN�S�k"\�� ��պ�A��f�*k�^��i&Nr�T��8�ꒆBE��?�쐪�����o�z���@.�e$X��B6�<̒�ex�����"=��Y�=;�i�2��28��ҥ���۰���gL9�� ���;%��aϤ�nޭ���]+��ኮ8�X�0�+",xl���/��ES���B��|Z��H�0X�-�����z�:�Y���������l1��~Ĉm!]o�Bo������S��`r�&=]�_u^-�'<~dky�yo�����>߬�}L�}&v��x1�҈JX(kEJ��@����(�\0� xK�L�ҬG��И�p���j`�$7eD�w�"I�x�U�V�]�����x�� ;��3���x�}��B��"P��_Ô\��W_���gpȨ� �u*IӶ.�ɭW<D:w�t�(����|���n�qR��HX�ΒqS���X�a����pFE��k�9�����|`%�qb��{jT�;)�u)%(&KOPcJĦa�z��#���[/e�C�UEE�,0��X�,�Բ�#�n)����0L���{��~�5��]qwCK�&�j�X���`���ÝQQQ����-�9�GU51�L�����&�Mwd�X1�z�y�k%��)_���S�}��mWf�Mx��Aiw"��GK��|��}�M�S{���)�|�J���-��BCAR��4����jE^��7�m�맄��E���YU���A?6p[_iŎW��9���_�;���U��C����O�R��k`yv�zn�Һ���]a�Ɗ̮�/g��\{n�_�!�EN�R�o�?=k�E$�Bޱ� �)�V����*�v��Q��cs-�v�0�9��,�M�N�:��knv���b]JE��8��k�g��Yh>/��zMC/.mz���Ƃ%#""Df�9ϯ��Ro^�*�A�l9xt�lX��?������_��Q�.�1���d�{����;^�8��Ε���ެ�Q�F$�dH�$v5*I%27���*��@�3����u�\�#��3�l����{�i�+��M�>)��E��y�(
��8a6�8�|����:�>Gm��>�/I�Kt�'�)�rHH^?e�����Է�e����*q�R,R��1���
~���I�C���8��� �2���뚣UeE��O�~��ʍQ��d�6jxku�/`׍9�(6><R�G��NJ��P��|ᷨg��1P��0��i\~Ŭ�Yi���a{��.,�h]��]ϭ�cx����H�9��9���Rc�Å�~A� ͈�E˸rz���1rN���C���6G�<�=wA�JH����R�g,�"b0�GU�v;��\����o�[���lRFT�"-�������Lk[ ��Ty�ވ&�i�A���Hۿ����+�.?�:���!TUnu�E0��8��tz���6w�F�^�9ڈi�Mx�g��v1�� قm��#����b��nv�N�k�/e���5��L#�D�ҙ���WZ+�c*��1"�K!f���CG�uYO�Ҳ66=��T�^��{��>~�u�G2�'�:��|���r%���k���Δ�P�v�i�)�^?S��o�&m|�,!�����?-%�J�|C*0�kG�2�+����$͛�}��7��K���d�_Y�C�`���[�v)[���|n��%a�=:���y��5�6�*ڔH�_{��&��܏e1{_+�ug7�=�����E��òD����gD�u�d�2���UF�!/"#�5Ƀ�׭�"���Ջ����%�y�K���l0Lgݯ��@��
Dq�XRq��o�3:Ś0X��������dy1�|}��.*	yt��{�ڎ�aU��ӎ��]b��S�۾4�NBȈ؁�\XY/T��<���!I�ܟBe^���_C��""l^�a��͙�M�?QĂ
��BX�(�v� ���4�m1�Ƨ;"2{S`Wx��F�(�\�e�8�LiOlj�B	�];��_��=�'��@o�Z&q�����*��ՙ�&�x��C���!�kd^C�`�;�fU���r,
�hO��������1
 ��� hʊ���;;�t��vµJ��-c�@�+���z�U��C�9B2/�k�+;>�o���椿o��z��@��l��.?�a*�NH�Ӑ�و��8/FGU����G����N0���b�t�̭�7�����&eyie�����<�,z%��-f�%��;	����Ζ�uJU�4�됅�q���#q	^�<�I�XMU�}~"��LGQwO�[LpdM�'>\#��격�KC��+�z���D�߽#!�Z��R�|ݬG�jQ|#�.H�BG� �W}�A�� ����_� )~r�[g<�D�];�aAR�d��nTގ�~~W�gs�3Z��2��IQ��I������Ȳ�͘b��a��.h����f�13��C���\��k���+fQ�0��U�e��N�\���k�>���QM�T�@�^I2n������d}m�YY����?o�N�ЅSI�j�?�PЌ���C����H�wY�)v���rG)ӽ?� �~~��x��v�9�v�L�:�zN%yí�H����B$?���N�'�>�a�36`�����4֓��n�'���0�����Y���9�$�Рgr
��@�̪05���\X������4H����'�w53��Il�e�2���!����M���`��4��Nc��s��K��w�Ө�躛������2z�ݠ�~Wm	��x�������d�k;�n�X�c�dG�y��٫���o�c��;��ٔ3~%���h���fX�VsAm����
 emȕ���15}�T@�	�I��8J΃��p=|�,��A#F�5y�:�Kі����TU0��"���o��i�q���^�j���&��\�ذb����Db��]�!�#��Ջ��K�C�+6�\�h��EA��|4_��u���R+���oL��
;_��&�I�⊂k.Fh���xe��a�!D�L�(]�k�$f�w�������O�E��D�Ş��K��+5��2��{���&^�)�(`��v���nBu����|jgM��K�zPw�;����:�z�j��iYПWm�7���g^i��D�o�L�i�ړ9�Ռ~�}'B��/82����H����۹��jF#E�4�kv�wӖR���]��N564[B?��|M=G7���b��h����B][���\�|x��0:�ӥ�!\�K�	 ����}B;Ԇ|*��1�ʛ���!ǷHVE
�*2J�����Jy����ğ*s����*����'�:���v�gW�u	@/�mu����9vq��e8/2��,]��T��+�	s�����W��`�S�ꌐK?�����!ڲ|��e�W�.핳���_���ZÐ�e=�h�c9}���c�8����.�����@��;^A�3�=�5a��(^6��s��G8����T}��R���!�0:�҈<����܀`�î�(,&��y�~_y<�f�����DB�dK��P3}�� �8�0�9�����'��Ӽ��е@�!�������J�����b�_A<�m�@����GA�l��W������t���k)��I#he����L�G�����/�8�/����e�m�H�ۿ�ltxmct��_����A��/��������DFCU-ƹ��[��WZ�.���I@��a9q����m��+��ca��߃cs���҈�D��k3�^�e~�	{���#��w�S8K���l��xe9��O��Nw����M�F�g\c�ﭭb�K{���_BX�<!�Ja�X�P�]Ն����IJ90=���k$+W}�_�.ي�i�����|
�~؍W�(�h�CX�������J*�c[�V�C��n�[k^?p�ܣ�����\��S�Y�����jy�\��D�A�����]U[�G�@�5}��z���l��oo,eE�*S:�
��,�.W<���Ut����y�7��:~.�<�����+��E��߻����:�њ�q�_3�ԡώGw��b��56.(���9$T���� V}��%{0���M���[fXi���>�G�R
ZW�m8��0���[����G�~6����J���n�v�>k�5;�ٲ���{59�)�1]2%L��z�mӝe2�{���C�f)��y��f�q;�Į��"U	���2�W�N^��}�>��C�o�ݤ��		��`&R-�R����d(~�Ő?�B9!��2���CD� GS����y�2���~�X�t�0��O�m7����I�"C�2�K�J��3'/�pUj�h��@z@��u���B���JO��HB{��f�tA|�����%J�'&Ҩx���D���aI>{[�#Q�_E�Ɂ�֞�#��H>�,zIzC(+�3�q��ŐŅ�±�=8�L�Zi�?f�{|�r�_�����$W�Il����r�V�oA����X��8c�+=���܊Q��R�^��Q��v���n�5pzT�.ƨyd�S~��.k	H�[�ԙ� ���ۄ��kF�1��9PK{���j��0%���IV�����LSZ��R��Q�v�@��9��f�Œ�x���R��ŗ��Lǵ���UT�컿��l���du)g��9n��+0����j�ġ�}�7V�)^�ys�I52j�G��](�N�+�f�ݬKXx*���pW��B�i�
��#ȅ��h22���\U�X1C&޴���vL�V�E�>A���o���&�s��\|դ j{��wZ�v9�1�1���8S���h�l2�P���h���Ɵ��Lb[�h��=(,�u�2���/�D�Ⰶ�?kޡ���e7D#C-0C�sfg�{s��bU|%�$d����
�I�''Ȣ�?�r%�Z�`�~��^���%3�\�|-�Z��(ԙ�d�����H"��S2Z�p���xvZ�>$Ud��Op�1t%���P�i��(f\�]��\ܺ�(���Ө��+��c,J=���w�8e�~����i~���(�G������y��n�G��cDÙ:����b�v���J���ύ��M�_��U(|���`��(�qDin���vJ��Bͫ8[)�.RO�x[e�g�_��1�0���%"=Q#���b~3Mu&,uC8K�Ⱗ5"��Ϛ)�\Ҧ�2�d�X�Z[�
l3\
)�٢S���v��ͬ���Hm�ޕa��@�o*L�4Wp��x:��X����l��#���EM���L���a,;j��;A.ی3 ޳d�����@�Bo�T��-�#v���J��*�=K�&Z��z�g��׉1�	�W�;���$����V�4Z�҄�Ӣ��-�+�K�"�5�{�	t�I�-B�����A���ւ�$��2_j��[�3��۝���tx�1�?X�H��2�UԻ����J�>h<�R��4��7��0^H���S$*��놙�4F!!�1{����7��`��L��}�q輪@�8��M�3�%٭�;?(��@�c����c�F+?���(�% 1XucJ���NR����ڙ�R ���V�`���#�͆ؐkU�uEʳ�;���E�nC�R�Hx��٥]}���" ��wD���@�R�2h.+��p�[�|/��:�	�~���G�qH��N ����� C�]���Tr�v��gig
����ͭ���f���Yq���4�>a ���F�Ic�/��+���uI�_���z�$�)N��ꝡ6�
�Lq���� ]�Rr�It�I�3.�a-!���܇���Κ���t�JT	�*$s�]n�,Oę��.R��o�������<d%ٴ���|&?�*y���!�~;�齟B�8BD�ԡ�Q^� >*�����K��S��[��T�F�@���0�4��|�y�$��ش^��6�R*��n������9�u�Ms�88��/o����b�՚�oȥ���Sby*��4��t��:,����F���H���.`	�g����:���-�H-�\���A�,���������=n�V�ߴ�4r���c�4�E,�_q��%=�k��-y��?���'sw��%5'5�"�����Y��j{�roTf�&�0��:�֬x��̻B��m�n�"�E�2g���!MY�~�=
���/�BS˺�%x���@�f䖘c��S����"̀�g������2�'̖���n���!Ӷ�_Ӄ{ș�D(�q
�8����dA���~
;bkj����';zZ�0D�ٓ]:_�n�0��Q]�tW��r$`i>���c%�	}_!�����O�z;���Ó
p�*�;r:���'�+��p\���g�y��Lx�]�e���!��>M<�$�R�~�S;_#ϚZ��������X���`z��ॉ��OK'<ȅ��Tb���<1�Ë#WUҴU_�]S&�L���U��!gLd�4jl�G쐉�GD��K��1�~�jv����#���.q�`��E�m�V��pY
�$C�\ /bi�U��h9�XWQj�}�2��o?����q��2H����g��7��-�5,ר��Y��s�������~�n��`Yk�(9�# �G�e4."D<N�ͭ�;��2x�>��1��dS�p��F]��Y����ѥ'�� �?M��D����P>o��Y3x��CTR�����û�V��`	��s�Ƹ�K~&My6jT~�Ө`�� �3��~� ��\�55�y��ϔ���ō�A����R���͹]��x�>^��];��P�]�S�+&fyj�z���w��N^�D$;�
δ�K���02�w������~؍�H裏�<2}�H$��$?)ء!� n0u��or�ǎ�89���E�/Т�7s��x�~�Ry�Rر⃮m�F�x���b�(D�~�1��w�:�<�p���o��5</Ü���ez��~.t�F�_��B�~o�m��p"N���p A��Fr7������Q���g8�ɧ%�K:�<��_�>a��y�7�n�ۺb��Pl�Q���ƦQ��{71����^n�w2O*ی�.)�u�YH��0~�Ȇ��=�d�e�Vy۸
�wF��A
� S!�lG2F ؎��\h+�ݟ5�����G��*�Ǥ�Ҏ����<p?�ؐ�j;�.�X|D�pT0�:�6��B��D�W��q5#=U��Ҿ��%��y�P>�}Ӻ�� S{򉈴��|��R�˦|��A���p�U�/\>]�vS]��� �3��l,��gwr��S⋰(��2�	1��PGJ�*�3_��m������!��)��A[�<�ڴ>dKT`�
��=��T خ���BL�"�����'q�i+��*NVqB���c��O���T@���v��F�h��]���q^�_-��f>O1��K��������F��PF�G��p��˦o"髽^������v-ƛ>�
%��_Z�T`q�Ǳ����3��[���r��~٭���0���[���|�<�>���nP��� 1�í<�:�dR�'3�r;�������EO�) ��~��_8�L��N�I�- iԊ�#kf�
��i��%AѤԎ��������ɡ���,���x�SU��c	�fݻ��j�M����W^^/c���Ȱ%J�c�����o�N|��zt��l�ި�xO�����x,{�=�'(g.�/T������LJQ�mT�%��C��m��5��"����p�����p�&���S"�_P��j��u�BkȺ�Er�S���PA�����(\����0��!���{I�i� ��8k��8,Cެ���7B��:'�f��|�4��p?G)V�'s��:�M��t|;BK\`Lx�o�@���Ԑ)�j5��EȄ7���i� �.���1��2��	���/]qF��ٞM=�].��lՆG.<=�ޱ��$N��X�@��Ը1��_�\1X� �~x����Ԏ*'�_i��;�6c&\\=�5ǡ]w�V=�Ǚ>L�;�5�F�z���=�0���Y�	�-��;�4�C��RRnK�;�3U�v&n?[����q#�n��Ѣ���"�"̝���pZ#�?��<�a\����G�3�	m����SD�h	��e�M9V�YYD7�8�"@y��I8@��>��^�.�f��]L��6T3\���&�E��^���QT�O����{�1���L�+�u$����	��1�'��O"I��/�{��������������0`�V{�2��f�N�$�_�g��/��|�����n����m(�f��~��B�8���Y���,!6`)����@Ją�T.{n��GE�H�]NfP`�T6���a�tH�N�=#0y���5��x�.=[H	����gD���ݟ-c�|SP/'z/"�2j0��^ �Hp�x��"����C�`����vÖ-�*cOD����e���d�L���ފq��`�՘����9:�����^�ȑ���^S:����'�_��Q�ܴ�����H|ڒ�F�lU�j�?�,yf��m/퟾{?�S�|D�@a��V9RPex����u~>�"�l���ƫ���}��\��f���_ k��k/�O�4��m���C��U��z��>�%ǏG�R�1jv�C����!ͮ��ucU�NC�B����ц~����� @N*v�v~�ľѠ�M�k�`����8&��XJ�TIh��g��-x"ݤ�47�!h9�:H,��1���:A�q�E�Y?��Ҩ�;�5�r�c�O\LN4��_�v����TPP�7���v�%4Y�&^Wm��	lM'i�U��U�x^�F��C��g��J�3^������8Կ �O���K	h܋��,:��\M �_d�*���q�W!7���e0����:S��,��I�r��������5�a�˱i.
��X����(���7F��;n�%�4W�_?���r���_J_D�9�8t+�q�{΋WeA��E^,�yUJ$>�����l�=<���1v�Ko����i��ᩑ�6�E��~��ym�ENf@�|����ci�Cg?���#�)Dc3��Y�]���=��j�'��!���.˚v*` ��c�,*����[Tm�>,7%%J� � ��H� J;�0� ��A#"H׀t��5�t1tC���x���ó?�/{�k�u��\籮kv}�f�E�?��2�#�MG�q޽t�7f.:w��ɢ��[�����E�b���V�Xٳ�.�6���YM{x���e����?�h��ƶ��6��9��䧘x��m��)R*���g��;��67�G䕸����>x��jɁ�֟�����E��Y�pX��Y�G�f��-	�d4d�[?=xg�R�%����^4f��͓��btV�ys嬱�In ��M؛�~
����`!1E/QB�������?�%� �)���
����y;��d�~��j��E�f�^
E
.8���f���Y̶㽈)*D!��Ʃ��Q>+	�(�%Z�����=��/��ڧ��T/d�f�XG�tV��6Si��,TK���`�~޹\���%H������a���?��̆,�?���f�N20�r�Q��Yj�PX�"@T-�����m/(�g�i�Œfim	��=2��y�n�f^���Ύd|D����ׄ���]�^~�(_����ߴ�m��d����9�O��'f^d+.j���+�|f'�IwS%���Y��f�?��y�3�����-��2�f��n�j���!!���D�]n۶Lץ����1't-�F�10�\p�?5����z���[Y1[)4Q1�fM8�N5�'�u0�FTF���4���[Gٮ�K�٘�`99�3��?n9np�[ɜ��8�ԙlZ�hŹQ}�l����Y�s*Y�z>u������s�6����=~m���Ti��?^Uf�l��BGgJ���C<J�5��^��x98�e�ò���e�u �uf�6z�5�%�A�4��ԅ��^?�.�7��v�}���O[�4�U����t�Sf]��V�Iڻ��X��{T�eͲ؇�Q��b?f�]'Ğv�v�x\ �f���"7��z�6N4�hш��qc�YK$�p��0����u�ġR;�QMV������7s� �?ӓ�!���,�!U��`��"+�CHK��b3�	�4�x���Cm~1��viE)�Bz�'�k�9Qyr�LǇ@=APiz]~���5��� ��E?@�wQzY���΢��zI*<G�=|k��OO����TȖ�H�#��E"h�[������O�r>]���D-9��1
���%�,�6/�^�޳@2xġ�:�!�r�j+�t>�\�l�b?�h��B�f�è�zC���*|�s�Б<=�$���ϼ1��r�,��竟�i�oԚ�.$��I�x	t�ӆ�h/�LT�p�?Y�N&�E9�
4F���Yr��6[Й�O��ŉ6��}����⁆S5�g��^�QŢ��\r�f�d{U�*��}+��������MX�B�w�7�<1��2@�<a:�t��_��
<��)f%�ҬH��:�M��7�h�Bݛ� �:���~�����E� ���1/�}7�+w�p��+m�GfQN�8�!/���=���c ���4�EbcU��|�ɦ�oU!�zr�5U�o�5.Ջ�RA��ɖBأHA�}/�)���
.�sz2Z\�]z�-���8�ёoi'�"�<FB��F{��8�_'��7�<j��"m���1��t���:3�\�ct~|w,A��d\K��ď���_M�~PJy)���풿��W���5����ʳ[EصfOLm髸aG�'����R�/�~��>��S�{v�W#�|$�e��n�:J���cl�ӕ��[��)�1���>�ښ6��{\���N��G���g{�B�)��{�O��aax~�u~ ǲb�����=Xd�q}�c��~Nzr�i�6���[Ӎl���K��q�"Z�$pS�i�r#OF_rR�|Sʞ��V��da� ��r��8\��dU���,��?>�1#�
�>I�ǣ~;�wtX��?�W�-]��o��q�S1W�B�g͙����-���������ۣ�U���l,���쩔�vCvPi�3��4�X�FG�/'�U&�;�;]"�F`w[�_̟ʔ25g�\�BU����tr���,�+}.m��͛�H��W���h�d����	q��5ث�OD�0�h�UZ_�f�y-���/��%�{�0=����V�!�l\7��|���:�J�7�ݕ������\t]T�n�QOy��DT��z����
�cߚ���ߺڜ0ǵ���#��-��3�����j�=F�*G��{���1Ǎ��2�Sf£�����^�#�Y�[!�) �F=�Ky��Qe��v�a#��N�֥�n�tu�x*1"�b�9�̍yh��?�L�8!�j��L��'���/g&i�'��ܪ�tЋ8�vsU��d�K�In~Y���2=u
�4/t�;�f��=s�!bd��zn6X��@g	�=T%�_���,�oSh�����3�l����/�\��ڭ�7��H��U�?}��3N�6Q�e����qL]�|�|�u�����j��2���mQ��.(3O�qږP��V�Il�V���{s^JTC%����&�b��pd�ǥP�΄���D��u�M��O���/r�gB��^+�6\��U��CO7sc��g�r�2�[vV{@�D��̉��i�GV0{�9�{A���*]�����{���$�=�Y�?�"�YU��f�U��<?)[���I��T/�����'E>��훎l�aD������n��t�{�A,R� e_�P�Ҿ�]�<�:�����B�vK��̴���Q�~�q�]��uϰ�W�
ǡG��w1}�;e���lO����`����D�R��'���+��5��N:s�� Q|��F�FBf��(OFO�^����a�FXZ�N���BCH�gQ�0�ʕ ��F�Y�P��4���p$o�fޭ_3Z�ѷ�Uiޙ=  <��Ёth����0�c��<�}������n���p�䇍�.u�5tuj���^_�:��q�s�2]$���x���,o�b�2��X������au���}�({����z�LB��$ڇycs���y1>�:Ʋ��T|�$z��h� ��(���Y��OX%���µ�#��O���u�?��(*�7�"��;��s�.Y��^�mB�;���Fڸ�CR�xp��#`��<�\�䅿��7�\�
(n-�Fe��uy8U4#�q ���D�ű���w��b�1��t�r���.��E֜q�=���QBe��c��?L�0�����8%JD��k�zOr]�n���>����v��H��͸����Ӂ��R;�ȅ̅ۥ\mR�I��rMq5f�����۪��}U]��6�޳��	�k�fQ}�ߊtŬ�@���S�'4#�T�O�Z�EXh���&)*�P�A��?��5����];*���a�R��zS�U�ؙX>��64Q�5,���1_���ٯ�	��ܹh�y^G���v���8��s���#Ջ��:7�Lz[�7�����}�yO�i�m�S=H���^���3�mI,8h�^����68unp��wc��Ǡ���)����"�%�.K[O�K@mHTɿ-�?����\��V�v
����z�۫cZ��~�Ȳ��iފ��l��@D��l��s�V�+������%��C���z�˒�����'o	�l����^`�2a�}�l���w��a��X�t�Sד���hF齄����;eA�Z�BI��0�<=�0�[#|�x�̠ۮ�����'VnS���(�����(`g��dWd�4���ȩ��]�ы�-��\M?�k�~���%��"�ͧ͝2}rz���;��	��D�,w(�qV�!$��~K @-�Y�\����G	��sE��NϠ�\�|N~"����'��N����Cҭ�;A_�Z�+��-� �x~6��L1D��q�eq�|���U�3S*��J��;o�Y�X��r�e7
+ ��ɫ\�$ (l���\(��q�ڬ�ܒ3��_6GthS5�]U5� �$#���n����˰�ih֣{�k����,@����ٹ���?���lx��̲C~�m���g��]TzLP��]��O+�������1uN5Ze�"� �s���gn�is�;��nP��r~�߮�)>�~XJ�8`�0犭�V�ɏ�ɜ��||�������w�y@��/�ĳl�m�G�����K������Fi�g��B�G����Q	��T��F]��Ap�Az�>\C����7�5�W��ͦ�������^ ɐ��ʥ�a-j\�a�+e��o�s�
�E��V��c����>Ԧ�SY�'F�?�ہ_�V���(1<ǈQA����@���L�{���![��d
6)�F׍?i ���
�sx�w�HMn�w��Ū��j��X�#�ہo��lP#�Ol��Zo�Fە�Dc�<���B��ϱ��HC��̒X��e=x�{Bc���A�UO}����ٙ�R��zl�Ƞ�CZ�����Wݖ�SWg�ɞR���K�Ѓ�΍���w�C��ʟn�<�3�~�L&�(�-훶2F�ܜ����\R}�/2P����ۦC��a�����S򛄩�Y������`��;0%`x��_e���.��Ӹ3GmY�GЗ�.�%��"m��P���ee�;��.Sl�x�O��Bw*�}-<����w�p�~%�7���Ǌ���k�n�2��$=�c���?؏�9z<���[�f�GC,\���r��5�R\#�:J��ĉ,#k=Z�-�u�>s�z�\����t���:=���Xx/G"�K�!��X�ڥp�r�DP_�܇o���1����:��O�V+��"��eRS�ꗭt�N�}B���Diy+���N��=oD<j����{ƫIm�8�?)6y�O��mf�ld��hh�YO�}-c�g.�}/5��!�Z��$�w�c�9�+M���S�ؖ�?�K�Q^4�(���0���9 P�����h�D�V�m���ޜO�M�7���T~O6{�JM�__:1CN<yfB����%���-�k�g����ƙ^�����z��#�W��7%b$�qO�ܩr�k���ę(�><,��^6���hu�
7�?�������Ԣ'_{,�_�4�؞m��6˞�UW�4�S���M�>Q�fݼa�ӵe[���C�x ~�L����>��\�� �Z�ny���:	�e>�Kn���d�?
�+Al�H~_�-�7|��Y�I.������(qLߖ����l�\�޺K]O6K��;�ҵ������%O>Es�Vwa�l5_d��5������~d�l�,�7-b��p��{�Ե�Z�㧞܍Q�M�HvHy����5uRp�P/S��%�C��7W�R�m;�c�wo�-�j�-�<Q'��{��j�2�O�<��g�,����*B��&3Iz��<�>Mܦ\Y9�V�� !'j��}f\�����GG��Lĝ�"~U�"�}B_;/?7��#`��]/9$�mJeEf�����u4�W��>�x寠2svG�fU��#��YT{�2�m(��㵓<ʼ��a�8�����J��K��%�u�m˔�ޙ*l�ӽ�p�i7�Յ��b�w-��t�^r�|kn�.��}�u��.�K������35G,��l�>��l^���u��A3.W��ж�ȱ5
<{���aS3Xң�ٽxS��C\��2�ܒ/��6u��1{[�X�Xw�R"*�>��>
��u�Sg��:��%b������@SJ	��'[��7�_���K�ZY�=�%�������ǯ��7|�L͋�YhR�X`Lշ~n�Z��ok��X?d��`
�)o^@n^J��5�]bju��Lq�qo�@b�3�81��^C�i (H{g��!V\8t{��"���3�o�����km� ��a���Ņ7Skw�O�[�S�h"���q,��k���t�ө�d�DP?ݖ>�8H�Ww���ڑ��QF��F��b����5�3���g��������lf]��y�����z`K11���q�S����I�X�\���v�0\x��@��Y�>��cj�1�w�"�m� G���~�>�.�yw����V2{wGmGk���H��*XC+�H������ hr�#q=��������u|��Z�Tl;��2ה&M��� xaĭq~���f���@^H�PX�Q !1�n?�Y6��;~Tg�;��?#�qiQ<m��$*�	uן���f�2�9�ez��"Č�ߖ�T�2��6}�-�=|�܇�?�n/#��n�^��);��9�i�eS�a�e�^�+#��I���}�L��|��^X^��}w_+;YD�������`�-V3VFǋ\��s��A�>n=��e�����uV�q����f�S���H�&��6&��N�$�Y}����i��p��U���"P0�mZ�ի��1�h(p��Al�*�F��XR��r���F�^�G N#�A�t��5����׾U�@�����LD4.@���r�,m��%XH��f�z~���V��x���g��Cޭeŭ�\�v��n�rt��rv	��ƫoy��� 3�?s�0���!�/�D9k��4����Q���}4pBFلWVk�� �_�y��>�tP1ɂ�
U�|��|jI��*��`Z�Pas侟!����E$Yأv�DZ����h5>��\�t"��{cQ@|EY��kHN�O_e9��KZ %˧�ϒ�����U��9�{���� ��Q���� ��?K���#���I��f�
5!� ��Ȥ6��7n�;ͣ�h��oaV��ZT1��R��z�.�:]O�)pz%a�NY&3�'�.��c'1�p�W_p:G>�Z-�B'
�Ų|����l�i�/q7��F�謿��<b�k�v����k+��&�յ	���k�����\
�`�7k	z?�����,�xJ�|�q�(��:vU��K��&��q;�����Κڵ$�p������/����޸{Tu��9]��?z�.�PR� t�I�b�B�]��ȏ�L��/OV¼Y�R�|��;��3dQ�
�U [�Uu)�$����D$�=D�^=_|N�*|��c�s���<�cv�{{���	 ]�]����2�l7Xbq��ۘ��*�"���k�n˪�����0 9����Ӷ�9�����1�qԛ&���k�e���l%�m�lX#ޥr�����i	+�&-�g�����Q�L���B��!*fJ�K��O�pU�m�ّv����R��v�f����mSTy�sՕ7��_��H���k��K�{�+�Ԃc�ߞt3��*��lۿq�"�6�Xg(��5��Y^��YP��a?>j�H��/u�qo�%Z�����+���}�R#��\�<|��.��b��PB�˵���p�E��J�lͬ{M�s��i��3޹���</�ץ������3����u�R*8;b�nPV�َ�R�w��P�`"{�(_���Z<6~^�o,G��Ƭ�Z���o�Ӗ��<]�(��s y� �a?����I�_�5�)B3fb�ڛu��>X�q=:�K��j��☻zc~�AA��	�WI�=}��kb�%�����MX�
���$�[��ky��HY�H�B=|�7�hlH%k�6��QNd��Ʉ�>�a!�Z\Kj��|�1���/�}qQr7���鏺yf ��?�r�BD5�A�]�2�̵�{���܂1M��t&�Om�OA�s�Q���ٔ2HHH�},����w!��՚;0'{��j�d2�#H�^����"XSy#���������gİ�?�K��<�+�I�"��i��gYAGRiq�a���|*
oɮ>h�sX���%$~m�%Ѕ��L������<������fX�TM(a�.;��>5�W]��\�>����Fw����D�geY��r{�tM�j@��26*7m���0_��{s���Ûs��e���P2-��D�Bu��h�(iu���fH��p��1�<���O�Ta�V���I!�ج�9���y��v��h�5$��#���x���Q��Ih(Q
�� �'�Ct'�͉�Gv Ңi.��q!�����c�(�P93��|L�#�RS�~���8�v����q�_�{q��f3"	��y��>4��WD%>?*zC0�K!2,o��[��[��_�ŏ�ݯ >L�y�<��e�M	<=[^���[?x_��g��$D���{�%�E���5c�IF�I�����D�NI��M���b����m=yr ��&����0��q?�zT��ܶ�����l����f���|����gͻu8/�v�?g�j�_��f+G��i�x�ů)r'�G�ٰ� �`8;�{����DZ+���_�=&�
��"�J��³bRY��+fO��<�w�$�Iƫ�,�6����g�=���Go4�#Gj��c��Ol�do۹T}�K�j�$����jK�Y��{�-�;_�Ï�#c�`���V�[�=9S/C:6���;��L�{0���d�&<I{+Y�^���*�g(���W�Cd��u#1�.�QC�((U�|���+�*#`|?Y�
oO�]��.V��J��ޢ��<&tįnVtGn���b�����U�ybJ5-�u�;}��C�ཆ���2�I	{�c�v�d��u��c走�\�2g��W;a��K�������#y�i�G�Gc����h�Q:4or����B�_��z�%��������>ws%�<�����Q�j�:i�F^�sݝ'�I=�=d��bM����s>��iH�ʌD�}}�����N�j����j��Ƿ�����R��|%0(�j�3�����![[KW�b��[�N,��c��P�۔P��pR��-�6�v�5� �s��F��	��D�߾t�M�{,y�8��{�q
�d�7��E<�h�r�ya���3�T��#hJ����m��9w��	�0n�.~ ;�HZ���&r�i̯��W�y�&���:�s�mD�'Я҆��{�
�%��5f��%�H磵~�əv5��J����r�i���6��]���|�F��Ӧ�s�.�/RO��a�#s����,3+k?	qvY@Rƙ�ڞ,�/2Wt�ɯ]���*_��i�8�P`�t+%����|VJ�����و$�"�P�r_#��w���
��')����,��mv�R��x�U��{l `�7ԫ�B4��P��[�2Gzn�8���VZ� �ҹ�0��-ֽ�Po�X�p�jۜA:ULUB��s?��P:�2��nb.C4�Obܐ����� �:��`�wK��R�m��Ҿ������\�yk������$kw$��r�8Psg�)���t���JV^��4l�x	��G��r�Q�@띘�夶Np�e�v�=���Ъl�oKrZɺSBU�v���9S���f����x�FP�Fbl��S@��>fh�	�:ٚ� ��i�{���kg�]S�K���-�-sylW
y�Ҳ��������劺�b\��<�g�x0R����֚6��w��M!�|�GDMZQ�o�����Q�	�@��VT$v��$*r�:u��\��+W��UC�7C)�7�~�IE�1p\�t��;�D��bx������hjv�N�ش�gU7�O��D-�s̫O��&���C��o+(�ܢ9'Zz�籡2R)n��`�Y�|�}��X�v8m����c ��-��� �Xވ���y�|b_��yNK��xe�J���K����W�av�Y�q��V� ?����(k�F�j���7���\�S?*�)a��#S^����9.�@�����3�޲|�꿇{'?��s��7@ᜟ��>��})�MyC�7���y����c�G�h�m�z��ճr�gg!�p	Y�S��)�b� >S���O��������$]��	�Ä#
r����DZ�t=�#h/�������Dtj	�R��>L`��=�ϕN�����F�-?O��U����!8��P�xo[	�&d���uv���~��6��\�t>L+Z.����=����OO�*�_~��ٮ]ƫI�M���0V���,���DX�{8xs}e����??_?+Y�!%�7H�0�	(}� CUZ�X��ႌ4#>�T0��>iˌ�`��0~h���f�1���z�;V���_��m���\������`U�}�˙���/���H��P�V�og`_GǮ�N9��QG1<�5ТYӐ��X�0��7��t#��ڧtwi�D���<"�S�Jl	��nq(S�p���j�N�U��HP�?\#����n0��3���u����-�	 H�U0�~QM�����#Y�/�T��գ�����D[th�A�}}����|P}]�����]�Q��e��#�Bη�3�I��L���1R�[N�{N�P��)-���3�%��T�4�����η����88_��]V�ԟ?Y�nP�i�w����Ap2`���8;�ir��pF�h�m�&�N�k~*Y�}�[���~B��~�E�m"�S��臖�YSTW$��~H�1�;�ǈ�-N����C/��]%��椼7�m���Sz:��)�,�*�,����F��nge�ɮ�媑�:gg�e�oW�:��>��e~�Pu�r���k�GM��b��]�f]�\P�]��n?x�M�y�;FTm�Ehl�T3C�C&A�)аb���h]��EU�4��	}=������>|V�[E���pŀ0��_�	D��
�2ǿ-A
pqm� ���s �������KņJ�.(�pި�^lB��w0'[f�%��c3��|A����^���a�Mi5��ԃ�;<�����=Y`X�-Y\TT��Ϣ�B-�"3"�ٛ�Ɏ!r%�1�ا9��w���9��=,?\�P���]���+Y�����l���I�{��e��(wU�e} ��g�8��]�/H9�^�W����#~�,C���$T���6Wk.��(m����^
XO�97������U^���+�G4\��m����j1|2���pc2��DA��Ͼ��
GT��I�	0@�8W[n�J�C]1
�)��`��*9�,qj�ţ��PA�ʳ�Z��ZzSV��쬓4�j�~��T!a�ls��b=�<��2�o�>��09�Ϡ��7y
`5V"���|~�`�ڣ�9�jW$?%G3���v�ι9<Y?X�ݮ����/j��!L�R��O*g�Fq7]&�Z���� ׿���À��5nj����;��ƚ� �3�����9?����
ظ}9V42 ��˄�}��`�'p4!31��9:�2ԁ2��;�$?_�>�n���:�1C�{����A�O��`�:��	�m��z���J�m�#���=�����.������p����V��} Ő	��'�f]4|��r�-����r%��Ќ�F1�]mA��.a�(o���:�̩�G�ׯlv4ɈX=r�_�.^�A�� �#��zk�[u���-:Q��G�<4�Y^��<�᣸�M����ݪ5o�ȩU�:����Nu}�����<��Yb�z��hJ"�ܜ0U�o���l\_����=Z��2��$ԗ�؀����!g��j��7�!�,���D(�z��Q8���7��B᪭�~�6n�DΞn��}WtmJx!���-�m��]Ξ%�{�C��E�
��	������nYb�� �?��yQ�t�ao������fJ��l>X$�?�~	K����W�ݞ˻8[�p��0�/�Z��k�`��������������婪j,6��@�ֻ�g�����ݤu���X
y�;��ScM���D{��D�dKY�	)���	IF�E�<����?������.ڒuLZ�*�N��$~����d�����[G����zS�k���*z�� ab�Bqݨz,��Er�G[�Od2J��:����d�Ի�|*/�В��kȮ����,YU�k\�^bX��bl8u��5�E�m�&����2n��wP  �WW�n0�4��D݈��Y�Რ[?�o@������|�?:����ʐ:o�#g�x�c���+YYe8$gU'#���809?Y �p>�
�(�}k$x��GVa$9=wW:U{�d��s�������#A���R��:Cx��.
��0��$"�9��QYS�iI�n�	�p��wY3�x�����K��i�G&�h�����W���C���;�q���_-�^�^v����ʳ���x�>\~j���{|�?�C�ݬ]�n'w�&�qv�L�'���
�����\���bf�Ӊn�g�ܤ766�\�v���':�
�>��g~�
DS�yiy@�FV�7�n��7Iɨ�u.Á�"j�E7d��7����\�@�U�p�b��S���:Mt���x3I�D�NP��:�ڄ�����_pn-��?�B8��,#>؇��x�ūB��<�貵>GRL�Mf����	��Z��{i�9Ӝ����dt��9�Ip|�,%C�#8A!oo�L��鿨���A�JI7���Lb.�^��<>| >j��.�5z$s!�6�-���s;�]{j!=q��`��O`DªL0�?�My&/lM��������g�����?��s��C����P���륪�J��m��PK   �cW�[0E  /   images/42df0910-34e4-4e6b-8fa3-2ad2f5724f59.png�yU[\M�4��[p,�Cn!���3�������.!���0��0o�����s�O���յV��RU��D#A���Ô��������?dlq+��FJJUNJ�J�������;'5YU]�(�x���Z(��%��+t�Q��G%��T��~)8�9��J(���,]G��Y�1��R��L�`7�|^��B�n��np�Uh�"���#�~����/�z�;���\3�&䳙D���})��:���s��҆�A{���3&��Ф��'����/�f��T;p;vv�F�[h�iPiֹ'GR�?OF�Ǿ�M�!=����Lǅ_���4"KV����4H6��d*6V�������(�U�(&�4rd���ە?���Ba�G6��������G$��`c��S#�"7��Y��|�!�?�=6�4��! Ix�x`�V�Z=��5�ywߙ�D;㌈s`v�y@W�0�g����F�X���G�=���H@='�W��_m�w�����K��m�[t��9��W�����K��k��M�(h�YI�4��� ��>r�VI'����>�����:��:پ���z�	3;�}4<�y���,<~(�S7�>J�~�Sh
�3]�>Ǌlj�>�/����&|��on'�1�
g���v)#t^���ͅnB��1�9����'.��_?�8Q~��[#���"O��{��A������W Ƨ�cm�hq�e��`yU���w��hY}L��K�J�D��؆�&���8�!�8����Tf�x�ډ��a�;�d?��Le߳E,��V%��ztR`T�2�s�6���[(q�yK���<�K_�9���A�����ʏ]�'p��Cq��_��%@M(��5-�U�d$�A�(JV�6/���L#�V�駠j���<�	>ILqa�5K�� y�aQ�4�d:������3o;�H�[x�q#g�G>"��A��&��M�1�@V±�,S�ڠe~{fObOrO�f\ �Z�Y��3�R��;��Wg�ֳV�ֆV�րuaԚ������+S?�n2�=],��Nu�O�QB\[~Y|Yƚn���k���Ȝ���J�T�8�x��[ɲ��%�� 侌2h$�'R|����ѹ"��Yik.�i�z~�2�p������&�&�#�T�E�^s���&���7�ߊ����,��'�Z��~R>��Y��)<蚢}�}J�ש�j��ꔸ�D��i�G�痋7�zԜ -��D[��M?6�4�7�4�9ʃgՏ���*?�f�g�6��517�ٺ��6���5KL�Q�x#v�D��ޣз�7�����s'O(	I������g>^;�EI;���&���i�g��Wb:��I�L;=�;���
�-q�����D�Ԓ��W�9�HV^I��ȘN�"}v�d�q3w�]�ݻ;�g�Н�"�O4L
R<L�p�p=�5����XKR6�r>_cEK⒏N��oƦ�xf���V����>O5n�&����U��,�X�YvϽ#��'��Y���5�7�9o<͊�<Tn�<a�'Xc^*�,_�2!750ް���oZ�(EL��1����7c�}?>E;�=�\�[�9�8��W%{%�h���lt� x�z��S`�S2x��2�s��-|d���]�@3�fVef�9���Z�*r�<2��6tV�ft�yns���?ŕK��䤙�<e���r��ݶ�~��b����������8�A}%b������(����:??�O����;7�<@- 5@��5
�F��AHC�A�����sha��c}�*��@�o;r{t����z6qq��`%�J,�LXF�D�C��_�(7�ڋ��qy��m��ٟ��/�4��d�ޔ��m��&?t~����
���F|�ʨ��S�t�l���5�[�����uX��G|7�e��tL�^�:���}yKs �)=�ǁʉ���})��ә��q7���hDO��6�2���(c���(�,�RD������(����)?��?�Ƕ)�y��5�%�$F%f(���,v<LD��%K3�:���Ê��h)��^��z$k�n`I�"����K}qq��5S����od[��},�ڜ�{[M��uuz!�R�G��:T`hT�La��f�
:�9!5#Y ],���a�gg?}�ގx��Mc3��tnW�c|�kX.�^��I�,|[���e�<B����T� )�^�Λ�v��E�f�5Jȣ�G�G�y�6���~��uT�42y��l~]�_��A)�^ql�߻gOeJ���+'�`ܼ2)1Wlv��{�+T�]����ז��*�c�t:ߴz����:��V�Y��x	�
x
�|w���@n�v,��X܅DR��,?8+�h��}�jv����s��ǝSt�3֣r��ꊜ��A>����R���uZkZu�Úʫ-��\R�\����]|9����@��dȿ�ӛ���<:s[bo��7���Z�HW1p�p�f�����픖r��'�[�s's����ݻVVy* �l5z`���n� xuC�����x>��p�{+ܓ �YG.¾�4�H.�~Bz�l�L^�uuw-��_� >��S=���ba΋��l�A��1>��F��Xвkp��eM<� �t����4�d�ص�����hN�Mb���L`|*}��eX,����G�J��/{�}k�ӻl�1#63����7�V��@i)��Κ�j2���1�9��2߻��cw�����2P�	��WB�x�*�q��+�s�E��x/X�M�3�!������U��xq�V�~O��O�����[� '�E⻷�iR���
����hf�V?M�w��������_s�eX�4����B}�K���e������9,7 N*Ϳ�ae���j��b\�f�{�	{�����m[��%�	�������SfAp[��~��.�?�>9y�����U�R��7�LW1�Yܡ�k�U@��������;�٦��I��/A�g�m"���^����cq���A��D���T-�,-[����%��S-�1����fHR�F2$<��a��\�5��E����o%q��8?������FRbR/�j'�Rў��sLR���n���`���ߖ���K�nV�@^[�v�9�>�'{��5����9ު��db��-�Oხ/�[���Ɩ�t����/�������#��m�{c��o#/��bڽ^G0d�'���mc7�+�)-��G������Ϸ���6�
[ʣ>qc��P!�Pl ��ϩ;Z��*))�_]�--o�d��~�>>[�{e�ySӱ���l&���c����ylO���Xo��2
l�r�޿b�MH�x���n���{�ߡ����^dX�l#�a@Eܑ��I���[v#��7.���B�^pie��G�z��*����.]���H�	&ލ�CĂ"�ʾ�������x��I�t,/��#�x��|--Ws<�6�-ܠ��϶'9"k,�Ge���GD+
~���`�Rk�.�g�#�l}��y��ݘ��#��G>d �ˣ�-�%�9�b�Nx���OJ�@����!��-�<�g��S%.��ۚ|�h�}}�S.�iIc3{�Hc�77���S¡,uK�nl^�~����1v�N�	�r�3�F/WkF���*���A�x����P���(�p�AT4;�J�'���J62ƅ驚�}-L���L>����p>���`O~�j�C�`r�압ԭB�[�!:]����*)+�⢸o�C�M�v��� ��#������;��ۥ��6�lfa���4�>���-p,)���5���nt��v��B����bѵ�|�k��֨`a:��9�6l��K߀��:c�V�f	EQY�V��Æxf��y?����'�����L�j̶-t�~?�����zs��Ƈλ��^^�CJJ���/�r���@gw Z��,��l��SK��:G��\��b)�c:,��{y@Ŋ������CCl�[��S/8d�Gq1	/�&j}D��jХ�D����?؝�`������"��������n��W[���&�rɫM��/���Ss���G%�б����'�f������OW��L=[��Xɹ��n��v�u�[VO*7��<��$�F}�.#��V�茴l'��r��H/����U:G����7z}�r�m���mw��HJw�笾g�hj>'��MF�0��^XX��\A���S�8r/��E�..�˄hk��;R���~�ӗ�����_fS�����e��Ф���Z\<��Pco�X�?s�t=z<7D-���&T�O�<���]����cO��Ǧ�k�On�X��|��UM��}|�������M"�|$���1�X�))�*���>\0��y��u�j����������QM���*���ᚘ?�o���$Վۋl�p:90�j�ޗ?^x�
XU���/�T�W�[q���#�n\�ɉ13^$mt��`#(o)~����1��^�����QA���������G%W�jug3h��j�Mtis��tό|p ���R��S����β�h b�����A�������/!����~�b�\:~��Y
rʞ�aH >�9i���u_��Z�A�*�bQ�KU_�#�E��.��W z�jb�}i�������EQrr|JX�k�)V�f[�џ�7�����_��B�	[�Xka��|y�>�F��D����"�9s+ʫ\�l��wb��DY���WĞ�{��� ���Y�X�2�\Z�.[,ƾ�q)��>G�������%���}�`5���O��Ɉ���'� "X{
��y���s�%���5M�#4dB�MLvG��
l�x�_�R��ջ�u9B5z�� I=_�`�Z���?9$�w9�~lv����_n��4��Ȼ0:�qz�b�lx��^��K��8:��R�Y�~�J �k8:���`0�-������y�{�{��؞q�Off�Gxf._�O%��h�E���f[ �������� `�~ r���ˍ0#�x��8��\���sw���POv�*�������7��tp�,�0@6��v�Ch�g���`����x.�4n%
��:�"dծ��~�^�R�m��*�
�=��iDN\���_�@��`���s�ǭ΃��Ɗ�J���8wj��B1?S���X��Ň�Ksk�Az}{Ia�:�N //2�� ����[!5i	�Mb{�{n!ǑT��ה����s�1po|�'���X��E
\��P��1�W��v2�~�� /�a�s�%}�d�L��� ���'��mK[U�8��K`+�\Nl��Ǔ���� ��*��G9'/$�!���xUH���)�����y�M���@��e��\����)�F��P�5�2�()1o��pX\i��5�]ű�pKU�'���4Gֹ��.'f�bu&�E5%�>\{i%�Ob����Y���#�s�p(<m�w7�ҽ��Dn�G�Ͱ)��Pdf��9�z�3�P��UM���&����Q����./�z��7@�����E02rX#�B`��w��ە9��F+�5�3*
���D_�Ք�Ϸ��h�%��~MlqY�&�RRf����{ ��<33}E�Ѕj̯ZB$[��o>����&�X1�|֓"4d�&Y}o���u]�t�����r}�q��~�YB���R�IՕ���C��݈;����Y���H�ʷ���|f�3�H��oG̴��������u�u}�4-7�N5�T���ĉƌʝ��l��VG[w��,k�TD��_.`wY��D����7�*����|l}���JĴ}��e��f��@NVBCt��D����6������g�u������\#�����7�E=g�=TJ�(ܕ��|��Yؙ]��� Ԣ�9�QCqq���!�E�D���M�����2J[���Hu�.���XX6�K'�����4'2�"c��ߗ���a�"��-w��nn<�5и�{�����
��^
����\=ga��0�n�7��\ �����W�����y*o#���&���67��~��4��nE-NCJ<����~�f�p����q��twu�
f��ߎc��Ā``b����qRsR���9Ϩ��g�����T88'�6�,�4���ӏ�RgAаf�[�3Ħ&�����/-��
�8^2^鐳3dW�F�ݟ&�2�aۯRĿI�*7c�"��=��u�����Q>�~on#�	D�[���L����12;F�3*+�cUJ�q�?��d���S�M��y>f��E���� �GB�(]�E�e|�ǵ���
��'���$�E��.���L9Y�]�\r�_��v�o����p�x�t�ڑ�n�Qjo�lr^����XXY��2�����B6D^����2���$v:a��Y��3u��ꚺ'�Z��X��sS�h_��zq��xܫ��i�P��[9>F�-���y��ŷ�m������a&���߷�T=��=��MwD:7?M��,�U�M6L����"�]λHq��u�����W_�ڭ�)x������Xϗ&X��:���9d�f���^���.�*A�ks�w�L�H3�$/~+k��y+�� ��;�����)��ş,���}j��Kx����V���\���6뾟PJؾ���z��a}oj�]{)�Uex͞�٘�Y��M����8����CAr�K;<����o�H���P�{j$�bVa���{�Y�=CQ��Ed�*d���n��W�f9� �t)ʢ�8�����?�F�b���^f_���A�����X�_+p-�(�i�kz��r9/{�0�͜
��!�~�`�j2g�q٩G���{�0i���O�����n��4L��3���ݴ�7sto��j���ɡ��޸�3����y��b{V�-��2p��Ǫ�Y�`W-
d����-n,�.gpx�g�o߾m���m-�[��I5�
Ǡ��k~aI��=�dh�կv�c���0���)^�B�QSU�QUU�A�V\'-�9og�V��h2��j�qb�$���\�w"Ƌ�ۯ����_���gQ�Y4�>ez�2��@�*��N�'�e<8 oT���s;t�_x���)�n^{���9i�B5�6l�{�W�����P���H�ۘ_��V����f�4��:=B�}����	����e+���-7f���Z��Q��� �b�z�Y��1���%5l=O>,�h����ݠ��;P�T�&O��GK_���p܍�m
tp��a��G4��씔�s�þ�,������t���������1:AKG�Lg�U�.ӋJtny����#��w��W�XBbb[t����>��ϟ�|n��Bv��8��$\�+��"���h;'�ӑә�)�����d��2A�j9Y\MNI܁[FP3��4ҵ�66#��3B�[9{j/*���񺡯�@\�ވu�/D�F�NAb�ذ�����0�W�5sm)�b�jIdI�� �Y�Řұ�1^�'��u������4�}T�9�l`�&�����G
#�٘�	��X�X���"�}bcb�i��⽊j�\�]�]+M:�m��!⻣V5D�b����u�iVx	o�Vw���0�ϴ�ܼ��C�p�Td��~fv�yY��1?��M9��v��]��_q�q�1�������D��:�Y�C�F�\ݲ�\�wz����]`( `��gJ�x�=f���"�J\������y�K����'hG$3�)`m��7�e
&��_N_��mXEP<]5���iu��dQ>^�)8L5�ii���+H�M��ii;Yy���|ZȽ�����|�,L��_���������FJ]�7�_)a[�JH�O,LJ���ۓ�z�/�(=e(j�}G���(�gM�d�.(���>:�$�����V�(#�SiSmsr�J=��EM3﮷b�L#b{��;"�_Rm����Z�ڕ�cG�aI��'�]~)�>6���*�����6�'������L���mA_��a�fCSg��eצM��#�D�2rR'eye��i�m��S5=����Q�R?�14ŻMg[F����O�m�AF��`����ܬ�k?���,�����|�ir�س�i?_�A�Iw��� =$��|��b%n��6�)[>�?3����#%"낔2�x�E)pO&�S?rr���/�)����ƒp	[ �sU���7�<x旇�������]�2J?��&q�{/]7�rg�*<�gK��y�6��Ƣ5o%�vk��L��UV������y�loW_α[AI��{�Y����ݐA��ZP���ҭG�(NY3���(0�Ş#6|x<64<������h��u��r�F<�����Z�yV��ϧ��[o��[��D�X2ܢ?��\BBvҒ�w����~�+�ޝ��`m8m�*��4	Df�h��P�Ua��$Gy=�7c�JN��b��ߟNڻ�����M��LNL:D��)�Ơ�hm��e�.j>|�e����v�%09��}s���x驽KYM;yDMh�G�`�0&�Crg�W�^\�R��SC�F.��:�>���ʀ�����H�pI��<�L�Js� F�J�z]M]�bb���M�c�x�b�8�^��0F��&ō��N���Ȅ��#B�v���!�,��-͖�Q�`�	6����Y���1
x���?8 �=���tk�> �t�մQ�Һ��8B��}�/_���-��n����ȑ:K?݄�0s�T]��<س�����n/"�b��uU�j2��/k|�y�	x���i�u	�j,#��`����S�����lG�5�� �����Da[[��ءȅ�E��6�)$ՊY����� �����B�ھ����Y��pm;3j-��A2�w=�����%���؄_mBeH�C�O���B-(P~5ܷ��ld�����~��L��V
�f��JLk����Y����2�������=���rA9'PB��ܕ%[ˇ���P�i��"��pi�a֥l��$�e��/?t�3$aH���B�>L�O�*v�d[�����PL�@���Mw 6��x���jc���Pڕ����L\���#��f;�D�T4�v�ϛ��:�m��\���)�h���.,�/FFB�x(:1Źٶ\���JXkg�˃����8k�j���L�_9
���L���6^�טih���z��j|˟���uY-�W�ܯ���鵐a��0t����gs<Fy�ĽIU�2<���[�W��	��i�E����g�o,����l�����H���T��) bz�w���r{>�TlNx>j��(��R�c��j�wu�\��X�.�)M���c�qD������Z�7���
*��+o��[�]ԉ)��A9�J�:�z�σs�tw�0&��l��6��1z���o�y~�����h^�]?)�AU��y����C�*ĖZz���&����a�êad�T�i�j�A�?�5����Q��U������ˋ��W#�P=,*6@�n�%�}����g<	%@�T��ƪ�+Z����̎xn(.@����5�s��c��Ŗ��S�[E�E9%%d23��jO��z_g�cs>���K����H�������h��b5/���ތ����$O� *"|R!�	8W���iՄd2s�9$�ާ���6⓳��#� ��L��?�!�>���G(}�ҎjXG��8}3�Z�X`��m�#���RO�!l��0�mjs�����^�{C�(=i��o�o�9N7�u���pG"!a*��MR��㇟��h��k������/" �H��N������Ѵ�s
UR��:$y����k`�E�^I���r�O�#�C�B3�(��<�Q�����gĥ)P[؝9\@γ�p�W�oX�{;��6F��c�
����w;pT�Ūo�\#ѻ��$-����ד��V���[7D����G�s�P��\���|.�q:��"�%{ޜ[b�w��^zO�@���^���S���~����b��;Q>�Yh���V�A��0����	����+��&/��<G�+~0S0B��d��1ݣb��({{<��l�r��'���=�v)��y����V���Đ⦪��n�����ꑸiADc����	C�o��6{1�["N�j�!S���|�?��W�-�R���S���Y"=C��S�zE�f��yAo���b�M�mP(��Y�@�촣��P'n`�pZ���ra[�/�Am�}T�!���� .7��],�	؎��s�^_KzN�m@�ߑ��캍�
�5���5������%1���w�Dd�t�6"���X�V!�)�D		��q�d�w�e�u�5j�?n�dk�W�_ 6���L){mMǹ =��c���� O�7&â9yar;�7S�����\0fN��؆�/�'��qq����U������4x�NUO�Ȉ�W�'YPoƥ�7��&�/���'G��#rc��?
��P�y��.k�<��K�?��*϶)S,�N2=��Ī��r�G�aϸQ���7�ƍ�*_ve{�_P �f�'7�2�R�T���D�ٞ�N�>�_$�X�#�.?
Rm��XYX`�&#~�/7��H�-�S��[ it?�ϒ���KJ�.�8OAN^&p�dx�T(�r|� }���'{�5�6��S�	7B4�����{����*]�՗ÑW��<k���Q�D���%��yc�,�Ե�R��I�1��Is�{g�"�$;�]�i��(��f�&�y59�w�)E��!$�D<'��h�ٞ�j�3*yk�S?|��@������Z�3��)G얃�Y��j�3'}�໦q}t�N,.�J�����=
��w��wW��B�¹ܗt�'��8�̰��4�����*"A\�Q������`b��u) ˉ+��,�z��`th�)> 	�B��#H����W/�\�fs��iB�9אn��򐵼��5�޷��	Q
,�X5�q��o��<
��.�>X
vU4@��t�6a����_�N��	k���:��R=��]�� ]��\���`�^o�D^FW��:��5����u'��O�� ����r��z�����
'�k��(���2R�	e��ٿj�YS�O3y�H)�z
g�&�������#��NV���Z�37�� w=QwV���H��������08����=ݍ�-��1��vc�E��U�!��Z2�I`ܦ�����r�Y(���ZB�[�*m�B�H@�q �WVV(Ik�F-���g$ܑ	�QW�.�Ϸ'~v�.��8iY�����cZiX w�8`��8)��پ?q
i�9��4��"\�W��w �kC���8��5h~��ʻ� �[tr\iL���u�Lч=�Gh,q�@4����6�T�:�
<�^�0�O�H���}� �?������ ��v31��Ҫ������_4^LC���<��xz>���4Uj���k+�֔��ۮ��&��ep��+���_ ��\���lj$| "���ΤUco��	�B/~_B�� �a�
��-w��?�#|b�A��z騪BE^;}�5+u���;���x�U|�Q�C�Wi�-���w7���3��X�G�0P�=�绥\��p,M��5�7���3:Kc�A�cE�`�K�-'h�;(���6g)��΂��6��N�W��#"l%�[:�|�[o��(N`��2�=���e���?-������.�$q�<�I���2!e#6�����.���;��1#_htR~�n �����vIiC�����D���oh��;�3)d�Ka�>0����]��V�3&J_�����롛ǃ�k����c�EF� ���� rt��C%?8E9��Gi�֡{N�JrS�̦<[���Z�1Q?5��9f����{E{�6s���R�|���`46��};3�̚��;8D�9��mj+��GEX@ ���y�
�N����p|F.I��o�ߕ��13�ϥ5�Oݟ�L���S/�o��DB�L_?i-ve(%O���'{��&:V���=��u{\��)���_��#(-��t�ːw��4d��^����v��)wb�$�t%zOlʘ�G+�=n�X��q�[���`n+�)͙�V�Ky��F����xj��\�A9{�
��,�LMw\LP�lW�Fe|�]�g6r�q	��&O�ִ�.��Z�-��|L䢔��0�X��=Q�c%tի�����~K���CHK[���^������K�����ȕs��>:0��W�͠a�Ɂ��5W��|�x�uaqZ޷v��␕yw?5a����Ε/φ�	'����s㕖�X�}���u6zp��_�٦WV��W68�e�]��`�)�0k3��f�Y��Q_<�����x�ܜM��o����O��J�뿴W�G�KpT|>��߳n��pgv�w��]�Sc\[��o�<�H���0���}��2�g&�5� ��G�i|�"�ߏ�O�ԟ#�.�s:��k����fA�v�b����*o���"�3��ӷ�����,�;.�s��#���<�x��Q�:J���S
�K��|ӧ��BEV�L'K~�O?�؄(��~dy��o��h��%�^GO/�B�k��Q�Uj��?�:��4|�Pf�Ūm=Z�����Ѯ/�'O�{��u��Ũ�/���T)��N�����������|=��W4e�܉��q�X�R�m�v:���1�\�9��:ǎ�UǾW����	�e"B� 9��(���=l������D�$�[LG���l��E���6fL˰�n�;��	JS���	�����t�q����@y˜>�K �3}�9��*]��X�ݙ�sl.�x���]֚�..��3�PEx��?��>����Q�1R�^�l�������X\��������{z)��..��^6ah��E	��'�K����3v�hJ�+�)��TsS�9a��
m�%*��[� Wױ�Q�&9)�c"։�7o��VZ3`B�t�`�߷-�����PWR���|6.�D+�D�����owv6�'�3�	G˶EB.��3�{v����kt�z�˜��T�&�t��_�T�`oy[�I�ո:���V3 q­�23��eO��8V�vIE�U)��q�7VE��g��^*֏LG��D�B(�i �$�ʉ3�yv	h2��)ŭ�&�%�Ky�t�<�r#�y���/���j�j��ͩ���d(�H��lH����$�y{�=�(�U�ss��4��� �}�#��l!tÿ�~$9Ax��mn,� QN�!c�cf�{��S�3�m"�{����t��8����_��׶�#^Fdː#d$v�]l�F�Q6��p���~��2V~2|8L�I��{�8=�=t_�}��<�K�]�𺳵�׽9	���������s{��6��ޟA�d �yo�OW�������+}�b=ю���-M�P�ޅ�+L"'��}�bA��
9O����9����4�k��1�>g��H�O�㣦�ժ������`�NuY��0qT���&��g P7fJ��W7A�Ǭ�)�=ƺ���9����Eu���'���@<�T��%������Ԓ���)������!>�7���"���罛!�w�[hR��0�8vA	�t/�?	����Њ�3Se���~��/����]{/r|����p��'=۩��^|9�
��N^6A==�H���+Ag(���B�����)���#����!7�o�	&&z��wV7ͨ;8�?6&�9��>��A�攔0��I��V��P�r~bl��,)����:������G��֘��74�;��j��)���z.���d[}�槧�nG�f2��=���;`���T&i�jMR��TG�"�<�)���,�����n�І��ٲ�l��w x̻О����b����\_����!��;<`�z�pq�f�%)l̨�6����'�hG��:dcʦ�2e�h�S8�:��eyEo��T���h�z�s�9�毇+'���:���i�L$�"a��������_R��X���=]��S��!c�Qm�K��,s2nx�y �u��KT:���,���i��8���(�O��e���f}?AQw��	O8�6�#Q�e��X
��-�D� ��Mp���.��"%����dg�\�ۗ�\ր<�ƭ`�>Ƀ��C ���$�w�u�GG�1�'��m��v���&��d����r�-��gna.�.v��IIH��pq��rS�.n.��A�S���C��#G�-����R��0�����9���\	��_��4��:��p�N�����&&����9e��Z��M�KNcn[c�z�ig*����ͅ����������'Z�c%�W�Y�vT�/j����*wq�L�<�ClW�{�"N��O�[�DU4 ��mj����Y�a0�� |ۚ���.�f���(�q��>�6�w�[�������eQ=���O�U�'�k߯
�6K�d��^9"�W��� W��˒N[S.��X�%�壛0ˈ�/�0D@��5壳 �Q��W�8�E��i>�ӯ�%�UF��hr��������\#dm�0]*P�h�U7��ob0��OJ�:/o����>����`�j���*(�X�y��Ô�X� ��u������u�����ױID�q(+`��� *h���� � �`�.:���F[�eB�ށ��j�(@�;	ͼ|]I���vyLd#���-ͥ����𸭷�-��ϔ��7��ż���HY�֎�v=W�Y7��<=Ξ��F �G\u5�X�Xv+�jkr��q��/-:���Ĕ$}ȑqO�_$x�KK�V\���@�(�7�z�q����@S�fo�ꈮ-o�_ONQvǡ�����1N����FZUB����G�� c�n3����E-���l���C|�K>.5�?w��c��`a����̨"t���<�9"	e�&sb�qo�<۬Q\�����^������'����zp��jkDgEW,���w+�v�$���p�@D��;O�wm�҉%8~#��R鎝�k��7�D5n�Q�9�ȹ
՚ݚ��ۘ[%N�}�
Эz9�I�� �����SyWs�ԔW�(_�,�}Ԗ��&Tl�T4>��DTs��2=$�?�x��h{��3��m�{:n��ٵocbc;��i�����X��=�k�yl��鉈2勇rn�
:����ȉ��8QB/�3��9�׈�n��73_�e����c��q�?qt.��0�"x�����и��!��h�A�Z�!Zkc'�l�+X)��7M�����SU��mf`�*�fE�ׁ끥��EiEq�ZIɃ_�k�M��+�Yg��@cIÓ�9�|�� � ��[#7��< !�%L'ĖK�m��ģ��U�Mv!���?�8��D\�L�s2�Hj���B��a���CE{$��A�ƴ��T��؉ΰ6�:ϛqr��������X%���M�ʤ�����D(}7�n�?��&����g�&�P����g�܋���jҶ��CB�A �#�	����׍[+��%��e��V|l6N<��{H��FRBihfWf���Ǣ�'S˴�'�)��d��
W�'���{d8���O忰
Si}���q�O�ſlp[!�)URa�g-��Px��l���~31	���ܭ��*��b\P��i�}�~�ꁍ��A/�ٰ����@j��,_�G���~�
��q�ӹ�af׻���9���[���4���koߡ�����=z����(�M]������̋���g>���r�tSz�#)��	�b0����ג�"�2��X
����r��̢$B~���R�$��>
/.|�н��W��J�ҽW`{B�K���9�ƾF��z�u*JU�ߗ[�6x�	�1�$��Oԓ��e,�,���-�hR���fn�	��cj\C�q��F<wIe�aAд�C�BH� �ƔY���/֮�9�|5�����a�s��{����t��)D�x�i?o��/��Y�Oi&�v����U�ȝ�5*e��Xy��o �4l�Gu)��|��|e�^ͨ�6��t˭�N�d2���l8�~Ϟ[���+v=�ע��}}��!��̀k�o8n^8	��7wN|���W���B0_�]���Y��Ҿ�W����1��O䍽�� ��z���^���kd��@����/^�'4���CZ��i)���/�O�.^G�Av���?:=��������US$���5j6@�'NO�7���WR�yޯ}U��Ҋꛇ�yf܌�����]4���hZ��`�s��ml�j(�Ǐ�z�Y};������K5g��u!�uR.��<����Ӷ�SJ >�!� v�0EZ>����? $@ۿI~z���5���<zw��82�^�ژL�hO����6�'��٨��ظ8Zu`&Y::7��O�N�zU1�6�vsgf�Pc�&А��ǭ�h�z��}�4�tFf���%��=>L{٘��	�VF���U���[XP;jw���`�1j�Ȣ�l!8�HƸfdf��Ht��<߆����R��9�Ѯ�Z�'�2|�Ӕ����������i`-��+X�e�۸X� �_iY�[�zHI4�|h������]����2|���˴�9�T���C�F��Vn��I�B���5y���9/q
B�o�r���t�G"8h	�x��Wz0x]��ׁ`e��0�<�ٚ���*/,,�lE��{3������'��Z���֞����-��;?��O��5:4,�V��P@@����X[Yi�o�uu��6O6���Dw͵׸¢�g���fd�'~��J%s���cc����i
k��216�$2�L�"�dE5�̦xq���j݁�D~��և>��9g�c�oڹ);/;�-����h��qz�k��u�\m[�Sc��E.-�֯�A��6`�p4ERD�ېL$N1��8�X���ӑ+0���0����;pȝ>s��>Z�b �E�uǡ2W���f��$�s�;91��G�P۟��+vA9o�Oˡ�ѐYN0 FNWp�9U�b-fqdƂ�5�eNvU�~N<�,Z����7�C��f6��$�q//;�k���'��^< 	Ƌ?�!� �:��Y뙸#�8�ΜtٹY��|˂9~^i�KGծBa�q��5�U
sb짦������p?h�MGK���ITG���Meн0�a:��W "��s�
�L��k��h��t��s�s5u9w#��{X	I(��䂳gN�USu�ӛ��7q����)�|	�/�S��{�����-P[S��L�DS7�[���}��E��Ѩ��o�Ϋ��G��S��m���j��L���3���į���r��;������G~S8:2��ˆ�Ϟږ���xnA�&����&�����>\Ssz�%�\.D)/����������hoa���y����>����6�c��]W~�_��p���n^>8�z�q �EeԆS\}�i����R\~y��
�v=�3�r�T��G�LM�� D:�҇�Ml'L�>��ݽs1R���*�U�.Hw�wH�z��J�&!���ؠ;t�(�y��(-5�#�w^V�A�����#��p�3d��D##ل�dWRXD�\A���������6��b.�2Qe�����
��9t~�.�VM��F�v�}�:Y�}��enA�<s�r���/[��=���f���#�c�ڐq�Iy�.̀D�w���LH0T! m�����&P�"*?�ڪW]������*w��Ѝ>�	進p8���T�}�]qq��������r�ߖ��&������e�6���"�y��,w>�/�I�_BB\W��������<p�=��WQ�Ҋ%��ܟC�����!�����g�L,p�Ȟ'���b� U�{Q7���r�L��,n�^��?�{���8�����K�̔�h"�c��f�qM�5�m���I���?������}�?���G��믾����ퟭ�>�����a��y����v[�l&ks���6�&0�$_N+�Lq�zyii���ʫ�Q�lΞ�(�H6t�ά� ��u�s��U^}c�;r���Fs �	8W��\^^�+c�zJJ�D�LS]��㐼N���&�G��08�pZ��b�c�0S־ �9���t=�2l��n���GqML~�k���Ю��b	 4 E�>�e���(�ǩj�Y|b*܃H�kW+f����������"����N��X�[*q�I:
Į���]m�:W\�k�2�HN�)��Z:MZVTJpbѧ��c�R�>%�[��(�p�o$@i��#�Q�2���ĺ�N�>�~�߸�!��1�$KJb0�x	����z�rw�Ռ��%�h���Մl$�'�-ߐ{�����=v���{P����t�jd;�R�67�]�C_����JJ�>�|���^&�Ë�4}����<����x��_�����	�8bOjTr�dR����m�����9G� ����1����'DdԎ�{���cL�-ѕ`�i!�͊���n���Ҥ��g�>��/��{����G���?����mo}��<���H�L��b3�P9;����f]88��ڒ������Ѵ�	V�&�rf�[��5((��9e�h��+����8��g���-O�N��	�P��3R�h��L �x���L*[�c/��Ocwg�;r�����Z��	2�@���z��g�Yl|��pNI�7�c��YG��(CX-�)t�����ОB���z��3���d��a�����6�Eu�\� _-a�\��;w�*DzR8���h�s��YU�$������+.we̛�@5���Z,f��ca")0�@B�l8нq!�?:ӑ��r'*�PitC*�9?q'��/��$E��1�����#��/��%�C�tL�S�=�9VSd=����-��K�� �!�y�q�Ήᯌ}�^����1�*��\��L�u�*�Y���p">3)N�@_�3A��ٜ����BwWzFn�_�s�ϳ���w�o,������;����J9���6FsV�T�J�d=Ǟ����4��Jd�?�80su#5�����ÛV+j�1Qn�2�h�BV���bv���������}Zݦ::[����|�'���ߍ��G��I5���������N@j��(�ED���0�s���Y��l�ё��1��Oh�8�n�ZyY�dUG�z;� ��"��*=%�^�L2Hj���mh�@�&�:�ٙ��6r��*�����xߎ�fWB&�,Zc\��L]�!�^?h�49�P�� N,���3���`F���M�d��[��8A��4�8��{�E��3�h��U�����	gMY��ԁ���4���w}]uՕ��:��2��ȹF������"Ļ@�e�������!X\A���1�9�I�t�V����mB�i[� �k�vw�G�&���?��j�������8\���E0��g�6"�]~�en����u�f^�"�!�֎6l��Qvн%M( �U��m5
��,[b<&�����w
:g9p��R!�g{�1߽�W��C�޸$��tI}��V����O��vI��c��򗵀���e���Ef��s��nh���v��C{!=)[�@�,2<��ہ���&2�P���Р�U�J����M�L婶��Ի���zM&�ԧ>��͛��.��X$ufM�\�`����Kɐ��Z���23����y��GJ�D�5d̮L�W���;����ￕ�姎9z����T��eY��)������Ʀ�!p0H����v�� A8��~G�o�ځ�i�w1�8�b$����Q�q��m|���>��t4t�c�~�KX���g��***l0�����&��nr֚�f�L��� �
��T4�����ٽ�g���C���������+�=��p�Cn��ݮ
}�MEcʧ���@���{�JX�WSz�S���Q>�a��0����� M�b�4�$��:�Hb�K���5ҫJYe�F֜ŹG��	��}�췡��=x�C�����s�H������t�ū^u�+�D�[d�)��AWUYõ�!��6tĺ '\ټr�WPd����N�>��O:*OH�u:��T�TP�E�dgg�+P9�1��=N�jG��ʽ�=��n��J
v]�U�KL�;����֬��E���.�w�/�K���f�;7�����o��.c�S]Y�Xt�-��5�`�z���骫oxp�::Z��V�yw�ɓ�3[�C���%�ޱh����=���C��_�ѱɩ<�@\�x�B�a��q�9�����G�Z[;�1j��ţa?��!�Jk�m�81 ^e�}l��z�i�&CNMJt��D�
R�W�o9.���F{�R*���LN9�Vj�8p4AG�1=����_���潫��=BM���fJh�ț��A�8���+j� �"��MTC􅒅��ɹl�?�zg�0�igi�aB�2[�d��=

����ƈ����K/cZ�u\�[C�kr'��1kT*����1y�@����U<�s	vgN��:K=YK�'��r�jT�$��M��9�p�*!��wxם D���g������h�K��ݏu��{�U�EN�k���@u��6;�]�7�p�A�챽�$X}�"��OiL��!�`JR��8�B`菧�����A�WA'��!a�"���V���6F���.`���W��yf:�����Ȑ6�]�ExJ~^-_�GA�Y�9_�W���̬�����w�?�|������.�v��]p���ON��1mҞK���uH��?�񏺺�jw�M7��;?���wj���'�C�#���B�-��ҕ�����nX��Pu�%8�Hz����m0��� �ue;ba�C�
���y-Fʵ�Y*� ��je���c�B��C�Z��l�RVRl�5��2�Hv�z�q�cd����� ��Ǘ�ob��BG��>��)�N��`���줺&b�\�=��?�L�g$h�4.dC[GS��`--�8b~��F9gsI#8��'v��� �wq��`��߻�@�kӗl���`Q<�`���Ƞ|?D���\#z�d���3�r�y�D�]S�&O��;?qQv��	t-�y���j��̗ ��!�}=��'6uw�(�Ӂj!��m$4�Ё1z�Cq��^z��Ʌ�O���z�>|�U�;G�=��� �̈́S�<B	&6�B#Y�/�?�

���Nguz��Ex4�����6C�����O���6��v	Ƭ�����D�����`�(��x�?��&����m�2w+q���.���-��}�WB���l �Mx�����5�!����y�\Z����2.�e�5��r���c,�e�����P��U�z���S8:���U3_�d�+*.q���7]Z��O�zׇp��{H6��bk����ɓ�ܷgW��ߎ��ы�,]��0��(`R^1�2)�2�}��{�W��F��{a�'@܊1����"��̤3J۶n��c�O4p��u��%8�������PN���ׇ�Y�:�9����a�Է��a���
ǉ��AJ5-ޓt���z�U!e�!+QJkd���Cq�攽�nO�}��nHz'��+ c&��ߔ�k��]�p�[��ju ,o=Az����4%M*{��A��i�����A��H���ؽ�. -���d%R\����ڦ�=-=�r�Ҵ�	<���������<���O'��%����9�;��s�pꓒ��.]��U|�}�oh�$���.�����v<��%�^�����|�ꍣ�-!��v8e�ʊU�F:������_�ꪣG������csߛ�Ăǌ�>胑	�Z�]��3��b�|yq�.
��h�`<�*P�����ޥ�x~�]7��;�����Uܽ��wa��ޗ�����_wvo�=?���a�v����P�?fS{�k��OhL��^�ظuc���������*��w����n���U�g>�o��뭅�-'��0j��~׻pZ1Gv�>����юm���T-0�PEk{��e�`|B�af��C~���Df�j��;�w]��4L�({�,;;;�����;�36*����;���w�����gF��y���~z�{�����.4h:�U,Xh��dTqt�싙\�Đ�����$51������C����(�	���lzF|``���%`YS���Ⱥ!Շ#s��_��/m��IW�b��2��I�h�B]�(UgO�(L�|&����b���aN~�,����sW��6���(�W˕}e�s-�OP�rڴ���L�ԜФ�k�����l�~J�O�r����DhÁ�IzUkQ�>���E���Xߺޜ<~�=�{�! 1�BB�g#���j��38�Z��=ˈq���HO�k�V���O�C��w{e�C����.���1<(2��7�k�L�4�W���BP ���}�nۓ���N[������a���mr�sɆ���i�R|��%��^���������p�&<��|����/s����g�vv�Y�����Q�?�/��
�_�;ȅ�2?C�0����?�?�Ž���;��K]���S�f��.|WSm���W��K{�j�w��U����П���cC)[6=�o:��e-8�a��_ϖ���]eir�R�m���`���ⲭ8���;�^��?��o������9��<��Ɠ�O|����4��l��Z�nYX"����e�'���Yk��xܕ"8&%3�0e��_��a�C�q��dor63���G�U�K]8���b����\Mu�Pb2�Hl���2sݢ���,g�E� VQVn�Ʀf�������|� �,-�6�e���3��-+T�"��إKM�]]�}}�獀.h�)D<x�(��ĵY��\�&�#��L�Dl���3-��Æ�����݃�wee%Η�t���v%� "B^���t��Q���X��|A���a�x�����iYkoc|-��B���O��>�4�����lw!�h���Wp%H�G�j�����N�x�ɉ)2�0�hI$M��t�g�Z��ꮹ&����'�����^�u�vU�c��	V,�w\7H��'�	PLf}�0�����&��0e�؈�ך �E#Bc��~^>������S�`x�6�]�k;�&�y��*�Z��P_���������J���U���e�R?CY_������x��_�¿uw�$˹O|��������:�����[������	X��:�x��7�&'�\��3�EyIGk�u��m�C)��z�:z�����ǝc�y#ҝm-�M���kߐð�d6q���amn�k�_��������D^|ѲC�UOnݿ����O���J���x���~$g��6�R�$s�`tmԏ�:��Gv��xK���6+���.
�M���8!e�p�=��ln	���D�����w��N�y��d}r����i����u�蹧"n��@��X[�z������޳�� /�I���\G�����<������T��[�����Q�L_�1��7�i�Nr@��;=qq��fk��4��';岀��3�%���H��q��2;���Ν�� 	eY�t~
dgu(�X��­\��kQԓU���C���	���P���5�%���#�E��z]S�;[y��>�������@R��<� %��^mxB�)S���?GϠ��8:�/-1f���C	�B(a�Z��]~�Œ�a��S�����C٥�db^8�<*,�&���=�2�'����{��ѱ�W*�PI�?+'�e�C����o6��&���,�=Թ0����87{3k6���I�0�g�']ѽ"ҟ�|9}!e�k�������5k6ly��P�3���֞���-PWw6���}w�x�S����ܵ-}d����Y(5��.���g�x��;z�g$1�u�#j�t��4��U�#C��^������ҿj��w]q�u?~�i��?�M��c�֬X�J������L��7��6��ׯ_������~��g����)����z"[nKY,ޓ��)���&��E�ŬM�sA�Lo��4���AX6'�C�L�u:�`Q18yj�8�� �æ���ܙ��]?ah�X�K�Y5�$ms��c#c:"� Ǆa�A������O�v�l�Z���x�NU�-�W�O�{����6Ǌ���4��6� �e�rdZ���yj�67L���z�/h�U���O�^�n��b�C���������--x9u����G�mg2f��y�~��yY*�s�F�y�thH�E�Jҭ�>���`ܟ8qҝ<��A�[щS��� ᫣0������旆�����m�V�mN�=
�Lr�<�q"R�n�_{�+-G�Fw�v7\�����I#�U���|�����k����UP�<�����(O(��#G.�_��1��;����B@�t��>[4���s��3��C�O����b���2�
���?�w�����$,�y�#ܱ}�;I��4�S���kݚe��60eLrdѴW%�lr�A��2���%�͙��V�,`v73�C27^U$!6F���Z*?�<�����������^Mc@��,q�+=N��уw�e��{�SQ^��z��Ñ�=t�Z����yٚ�4�#!K�XPƌF����ڈK�F!�I}x��"3N����]`Opu���9�;���
2$�T:W�G�M��N�)s����}�������;-�71�����s��ĺ�+��Ed��M�����"v��[�=	�L��sH�JW�����r���{s�2]��
������N�~�j���rgSh��O�;" v�2�G��� n���eԑ�t�Nj�}h��e Y\II��E�Jv�sCj��=M�@����ĸ�L���o�6w��{�!ڙp�9��)z�A'��mm*��5��~��Y2�p�ᢵ�Y,S��>��_y�6��j�����"���z�S�PС�D�"f��*��~�g���UQ��u��}�90����F�k��8��鶫��}#b� �����ں/^�9n�����g�v��2'%k���k���y�ޗ��&�b#�MO���U�U]S��_���Λ����-����>�ݿ7.h��ٵ�[u���A��������"4&���es���HJ��U��'C;p�;���c<{�\��j��[�V�\aҭ����6�@w���Ė������g�����7������ ��(�̣O{պ5����LH���6�����1H���o���359H�mñ�l�Z�.ں�O�vey�KHbl�(�cW֦;ǣ�6���5-o2VA�C�����V���.B��(�MA݈������y5���Q��^��]@��bW��>z�$Vhs�	���ѳ��b�P�����rB"e���j��9V���i���^�S�k����oAҽL�۶m��'\?/!��iJZ$:������n	����Ŧ��L3g�6�3��u��n��P�x��tp���E2�=R��l,x�S�n��s9<��Y*;��ds�d���vp��)S��;���c8�P�b��q)��W7�ˠ�_R��Up�	��I��R���Z7��zW�Y�V�Zf2£��U��}�����U?C��t�Yw
[t�>(���_D�Et�x�kA�:�&�/zz��@��8	|��(����υ<�Hr������9�D���2�W���C���U]-�^f.�j���9sU�=$�cD�A���]��sǎ��]�ߗ_T�yJHHz6C����4��!�?��w�+X����E��&�"m�N1�C3�{�dU���,�s��&��T{��т�٬w�݇C�v����B��w۶�W��7.�Y[M8���W]�ޕ���a�0Ǚ�8q�uu����ƛ��M����W��.� ������]D0����;�;8:�f�]O ��k��X�������'�gp�qӓc�SӚ�&?f��ԋ�QS��Ix��ZQ^��x��J��
>e���&�?��)�ͨ��׺��n���B���2t%��%-ŉ�>eb ��Ȼ@��1��o0���M�^�-mZ������%o;H=x�>11�Y�����{�5�ed3�(u�}8J~!��~�2l� υa���\B�c�'��O ��,m����!�NA8�@�U,�x�_��Ō�i�d3�?.YW�^F��q8H�R��o
R����6�ܰ��t72lO�)�q�)�C��嗺2����|���vw��qWMP��wo�G>ε1���W��\���S~��uT>!�����I�ūi�3���A�Ķ����]vf�kk����r�kvn�[�l�˂P*��S�DGO&�l"�S��S�S�>�{�(���q�ꕮ��ȍit�q �g���4lxe�B,�-	`�3��:���s3z�l߻@$���Y�oì����T�|��ˌz�u󚠠Y�ߛ�`�������EyHߡ�(/����g��gN���������E}=�%B��Fw������L<�կ~��]�H�"���n���V�
6LJ�^]O����߾���MI�|��;rx��߾�����t�E�"+.�soy˛��,��$<wC�sG�u�����2IV���b1CH$Df}�^�p5�^ùx��3dn��L/^�8y�T��Q�ݶ�)J8�C�mE�b�	Yւ�rZ��K-��Z�ʱ8�����P�F-S��q�Qn�(��J׾�0�d\NL�����y\˿�mL5y�o=���hy�&}�S��d��e��JB7�l^��cH����\f�k`��������}�=LS���px���V�x1���Hli��U+/BI�1�VmVFM��* �����|� �N��Q 1E�D5���j[�f]��{�u*m�� 1vqz8���>�=���ѫ�[�8%�B�5n�2c(�-vW_z�e��\?�m&@z�_W�����(B����(ЈONEfV����/�ءu���c�r>8<� �%�Q �n	�ʑNO�_���D���h��t�+a�G���y��Z�L6�:W_��r��Y���!�.�<T
��z����'��t��D������}UkW�,$ ��H�7�@$H����EQp�e��~xٺ��uy\=<&��m�9v�ϴ&���c��</01��~F�v4gf�=����	ɋ����?��/���w�/��}�l��#��N�|Oo�5�I&�f� �y���S��m�@�^��џ����{��>uǑ#���U6Ć�u�57,��.�o�w�7��M_{����YnKJ[qL[w�j��� ՠ5aJ��F�!臨)m�����K=M�-S���/X�$T��kΝu�}�@��睐M=4��ޅ��4��U���z�=�p�d��E5q���FN@�Ld�X!٬j�Kp*�a��I6��7����O�`�d��-_���4�H$P�xF��$� 	��|�Q�L�"����ܫ`m���1U��z�L�M�.)A׽d��Y���!H�*�imm2vv	�=���a��<p���mFVSH#�59���2��]�b��~�!63+3����.A�^��0Ú�,#���Y�qfϻ}�V�̇��6�G��*�L eŶ���k��k����쎟<ʐR@y�6`�G�=0�,����Y�0S�&���F�&��J�/��f�41ڽ��;̲N����CG���:��9>��s|	�H�'��r&�	�	U4.f��#��S;�fv<-���C)���կt�>�j+�t�������9�B��sf�2�$�P��0H�IbA�S;am\���(�tT@h�`�a%�����6���>D�3�s6��w>��q�S�[���|g�5�34���%7���j�GN��t�k>���vGx|��/����_v���;�����>{����3�W2�Ġp+��!��/�䲉�G����+���c�-_�|]���]?�v"%�ڠ�q��[���/yF�]����?���c#L�D���un�*�F!?�@�&0e	� �p �i �$���j�j��Hە��.FO=���h7����=z���!^���$�
�w��e��z�=j����V�s���V���`��=��S?չP�]�l)��r���&�A��������LL��U��d>�TɌ�{U�nE\�~�@���Ȩ��e��^QVFm8ivK"��0�E��5Sgnnn�ib����S�`�Ӄ�3oiit��Ȝ�2~i�+@Pvh�md�r���S#OOa/;x��b�������3�<)�2x�o���'զ��Q�\Ty�'<g>+g+��ٶ���v� ��/sk׮�ռ	����[њ�7�Ҁ�K�\N�6�l;�]>�p�r��摫E]��HjjSvnt=�S	���ѿ8��İ���vw�T%�}(�E$بO��9��Ț�}F\�b�����M�Κ�h��g�\[7S�h�� �����Z��A�·t�"Ȏ���T�D�
���Ϲ��Lunc�s�C2��֊X�6o�L�֋�U���.^P���b�E_�*`ƫ,������Z֌�,��케ܽ�Z��MN�|��C4�xf�E�4�6q�͈�Fq�+`���8J��+�NI���)˫/��'Žp����X�;?��/�+�L�.z�?���M �euT���S�RI�&B�XO������Ӄ{�\�י�G�����KK�~:?��S��NKI��֛p\�6$�MJY���f6�! �n��Q6[�r�ȡ�'��0|����|���K�b���T2�L�䷾��W-_�ᤎ����_��O~��iHJCc�ı#��rW^qZ�Y4�2�0��Ç�Z]�Fsj-l�a�,�p��T�&u��Y���T��`U�gSMT���Ū����8�����,�?��v��	������q�	�LRcmhl����i���V�I.=tO�E��;;�1�EX��~z��;!�u ���ƹq��
�Ӄ�� qmEj�[>��˙XJ��HX"H̀L����F2�JWS]e����D��'q���X7ώG.Ul�19r!	��z�u��I�U�0B�( ���Z����-P2#�!X�_%*!*���|��i�Y�A)��M�gPw�ܯ�w��e'#�#�`� ���(�u�+0p�j��ӫ|b���>*�\�̅3�W��pFr���o������� �q(�]k?��h���7�������Uy$�a7*����6D��W۟��k��J@b_B�}C�x8	��ض�e��B�L~6��{�N��ƶ�0��Y���N��pY$ĺ�C���AIj��WF���
gJ��.�hRx;QK�{������>����S)�7("~�?��%�/���w������G��D������G?�a�i��-�ooo-
��+�3�����=�y����۞����_�|g===���Uvv��l�":��PƐnf�m�qDs^0��ߪV����HO��<۽g���!�1}߿���o��Ω9W��ʪ���fE�ݓȞ`s��>�^��;.]�dݶ��=�}�w�����nI	D&��*�p�r��%x����^�T;y���8r�rr�0��4���������9�[�#C�L`@D5jʉqlxd\ʄ�{�1@y�ԡc��n`�iz�+�F)6*�e�pӑ��;�?`�jnH��{cA��Q9{����)'2}-Hv�`WW���J��'uX�4v�xW9ۈ,+��u�n:����LAXK0kj:�嗚Sn�=��U�ػ�v�{�U0�� ��Hx�e�#�|mB�E�.2B@D�S�$�����W\fus*%B�zX&)�cm�d�B0���3�S�,r.�NDuz58��[��Yu�Xt�d�˖.q�)̂�!�L���=�i�qCԦӰ�xB@ 'r��"�P�),�q���F�� j]�5g�����U#7����5��F�
)�b���]���+�Xi��,�:;J���[^q�$Z��n��Oп_ñ�~� !���m�탮�CA�7�«�{� =����:��f�B�6PPD�v�XwXh+��9�P�=�$�P8m�}�������,	��s@	��s�kY�gD#u�@����U_ON[�hDL�Ѕ�+��+��K��^�����}�_��o|���ʞn���ڻ\{���oٿg�w�~#���Wٕ��DK�ˎ�����Y--����O��ƹʳ�DȗԾٓu���0,�M%�����L[���%$���M7��2�7�u�'?���gEIٱ-�����ݣ��f��[��E�P���"�P������
�H|�^_Ss6�o����l�������_�l'��e	��5��m��Ͻ�9o��u���M[ϝ�o�q�*6D��� �3j�}�n���~� q���/w�q(�@0�s'�wO=�X,�Q��^�� j���H|��ѣ�l�R���U��62�,<*�%�
�VVj�X�K���xZ��/NBpuCc+�׏2>�s�Rv�d�L�&�'fе�AJ_�M�KNJ�l��e�89��E�<u��~°l�jP�"���\�6��VF�� �(;�#�೨1�= �;'��ah��ѡ0d�lD
��X�6؇�I�m�6Kaٺm�khaƼ�����)��є:�Q�Z������j�Yd�c�N�u�n�9����
��#�_�f)a(W�_��8B_"��0�t���1�|��ʟ��Z�<��}:DԌ{�?�R�yL`��._hB�������>�	Z��$3,�A�"PŎ��/sKiy�,��%��U~`��8' ,"���8+!��/��t�
�v�^BLt�KI����yF~�;zx��D��XS��!��X_j�0��p�m9��ܼP)���D�EfmdĲ����IRڊ�|����C�/�+z��Ϧ�W�������~��W��aT������������T���gz�U�-��Mk��];�߿w��ݸ���������{��bv�h������s�N����+./ݕ��rZyͩ�'�ߺm���C�ҘO�y�,`�fP��˾0gޮ��$���k���i����S8q��{vl���Ij�� �>t𷣃7�GǘS�6��w��(/����۠y<�$ل��nd*�ύS���іc�R�(�Pd�OA��	]{C�A<���d$%��kN���W�4=Q��Qo�)\J�S�{(p�r��ʽ}]dnGM�#�2X{6e��@�i0���G�Kf֜�:����3���ڬ-�U�ehԧ�Ed��ՠ7.iX��V{���`)3Wߺ&�͇`����1t�{DF�0>�a��L�Z��	6��A*x2��L{�x�t��
.Lڗ�CB5%��vΦt�9��-X٢$�*6�Fe�qw��!k���:��[h#�(C�eѼ�6^H/�f�Qq@�C.	x]SІ����G�~�+([AFٱ)���\�\>�)o.���^;2��PA��(�n���y��pi�]�;y���A�5��+�@�ʊKq�I��`D� �����	���]�p�א�-M~)��2�6h_3�e�8����^� ��n�n��E�Iidʔi��ԝ�u��aG�W(�KG�WAJ�B�� `�t!"��ɕ�W�2N�v�΍nX���Y��� ��H�˥������z2���.�K��}�#���;Ae�	݇=غ'|��c5u�>r`�G�ON��#yy�����g��g�/�+y��ǁ��o<y�Ȼ��f�hc��ڕy���A��)`F���xN���������������j�֧,$���fQ�@��i"���i*��tv,���xz�*v<���ί|�0#;�YY�Lx镗U3���k�rE���{^6�x�ͷ͋�O�޴-;]w�2��w����]y�C�fz4��\叟ھ�uA���mh6�0|*==�`tt���΅ugW����m�.V6fᣜ{kG+�]��5�aibP/��(!�M����S���h��{衇JV@ˠ�D��Gf�݊y��O�v`ݰ�WXt%�"�hI��
�2���A`h�{V�ǩƨՊ=x_�uSES;��/�����U
�V�iЯ������܃�h0�;1���#�H^1d��m�G�^�d��@� ����G�{�;xu���JK��-1�~�$v}V�P?�Ƴ
�W.���}��C_��əN>����=y�xOR>p䘧P�c�@GW�c�Wx�}���殾�*WZ����ܗ�(��߿�@e�8���,�77����W._�A��>�EyF�/96��M6U�1�\)��8�(� ���v?�8��y���G�##k]�d��n���ޏҁ��n�Ν�ȑ#n�7�F���!=��h~�E�V1���zD��-��j��
��E���x��b�ww�����j�X�%�X���K�r˰CQ^>��*�HfX��}��:�7��� ��n�~˴'���֭�]Jj�w���n��2�NK��'�]a���  @߿�B}F��!hW���%*&�{4$"���ޝ��+��K�N(�zO/Ї��/�w�/���:n���?����0A��T��������J3��Q�"��lJ-G�Da�������W�8�fG�����Q5S�u��� k+ڹ{���Ԯ�'+ηamcC�g>��;��ͯ���ˤ�yˍ70�Բm���9���|�W���'����]4����K�-=3�^dL����7�߳��L�Z��g�W`���P��àPe�8m�<�IO�F��<����pok������&��@�j?��\q��Re롿����3��j���)�TlaY�����걓1dfYlj��HdŃ|U����=M�V�j*?�:����Gɨ;q�'O� K��f������K�G֢SOqS�֧v-�|}��u�h�J8ZҨ:��ܐ�~�$@J$��Lu�_wǓκ����+��n��s4B�x���de�ktd�s,� �C W][o#Z�H �I)-7�:1���<��R�N������?$?�������r�^V��S����z�#�_�R�o�׊�}|�Lq���W�ZB�\O9QO���q�?J���7d�@zz2?w{����T7�nȔ�C��H��u�ϸ�%�+�C�cp�M�i����"ݭ�ތ�q���gM�n��#ǎ?ӡ`cZ�B������a����=�^s3T��ư.	�&L��?�A����O=� �� !n�QgZ��Oٹa4C7I"B���2<����u����Vx"ߍ��6� ''܉���b7�U�G\N�|����P{��E���H\��S:��k,����˹����G�8�Zyg^���O-��Xr���������'�������j��5��Cg1�Ӂ\�dd��#�iȔFG�ќ�>�ki�"؏����T�X8YS����C�����d�z�����3���&��w~�}���4��-W��]��)�z^9�Іfhw�6�ѡ�Y8�Zij������������wR�m����HWL�Hk�xj�;y��Qj�!O�;�NU�-r�� ��,y�9E�V+�9I���h�#[�9}�M��2"2������B��#��˼z�jہ�w����9�S��L91.�@�z�i�Vz�kQ1b��mJr&}�T�S����6��	e��d%M]S�!�l�R�&�C�����q]([�}�uғ��b��*����`��4P�>u��5nɢl�d`�W�����v?����=���!�CN_�Z�


-�6iR�/r�r��L��ȨTg��@1F�Ծ&u9e�3t0$�w�!$�d��tH~W}�����{}�e6�T�VBy�(+*q����D��09{�	������N� '�u؈U����H-�Y�9.]�����i{| S���[$;��'\����']]}�A�Bu��R�@Or�Y�n-�5�mA��hD��،p}U���8!r�
b�Kq���tP�WYG��*�(@�!+�a��M�#8���k-�K���Š:��P�hήAD�q�</�%�媭���2�~�M��a?"9 K�M+��N2v�R&��;Tݱ��ݪe\8�8
�D&��A����)[�!f��N";�j�1�L��tՕG\*vH&�(_��AѮ�q��#��+���bZ��	�e���9&HL����VH�Y.� ,<�!�����oWV=���;?yOz���f]�s^�[����X��Kt]�g��z�Ё��̋M��l$3����Ļ�x�3E����<pA����چZ�ȣս���K.������ԏ}��{x���r��D���A�;�a�E0��k�hj�z�ߋ�)2��3�	N�R:�4q㰈��Ş�|�wݵ׸�`XmX+��ջ�/#r�8�iph�Z�	8����1T�B�?�yE��7�������)j���}߽�7�G��b��BOZݑ7JM�8z�U�]u��5������0x�,���b9�~�ƂiE�Z�z����,�oY4� �ndb� ����A�&��7�� �q�L{Z��!���|֔4�ީ&䚂J�x���2�P�	��_����vMԟ�����x�l�0꽚���ژP�3��Ԍ����o�^WU]M %��#1�R?/++u�����~���"�i���t���}��ǫŊ�&�7DI�?��F����Is�Aj���Z���@��ʫL�F�Ri����}���#�{�Ș��gK���1'�_�箸�
;7�� ;�=��u���i[@��D��u�`br!�z�ew�~�cCtFP\EVv��@i�w13�rOk��z�%{��ej�v\�_�5w-E��'3����e�u4b��{��:���GJ�^���� �nGGa2۔A��[�t������pݔq�HW�z���捛Ȉk98@�hČю(��M@�Y����v�u�O�w[��xJr&4��B�f(�θ~M�k���]��p�Ϝt����[_��Zu_�c��S������h��f������d�%�T�-�`+����e��ɿ�����h�Ż9���{m^2+;~�����M���׳��HS����p=�ƺ7ɦ�1��V��4�"���sB���o�a��ؤ�~@=�f�k^{�k�_����������[�J��0r�������n��"Z��8��C�t"���O9��9��yN"�O����c�v�������Ae}lrL�IMY���<���U
�����[������W��~��|��w��?M�lo&S�s(۹|�k0�?ԿՉ�h"e�@��+�Īv��j�y����[����f.b���y�6}�xPe�ڨM6S�f޵6������g��y;ɰ�)j�c�����^�`�[��4bD��xx�n��ݦ���������-G�ߥO�"y��n�2�\�3AA��T�(	���Y�9�Y�2�Z�<�X�q������.y\�$��.�2ӳ����|qO��띮<u��ع��2~O�tJ������E���\�y��VV�eΎ�#�����l|���H�xi����I���`G�nd�Z����f׀�� zO9c���l�kÐ� ܣa���4'\$�1j�
B���L��;^٭XW�f <�4��,3�;!�)��B��2Ā$	�P���<G$�0!2��<��pͥ��`H�zg���VQЖ�6�m'>C0������ A#QK����6��Sqg� �U�9q�$����裐Ԃ�%�����rl���j�'�brZ��\�Q�#	*��d+���@��q^?��J}�͠|�{��u�@��r��sӅ4賯π^'�@+V��Ǯ�P�t�Y��kz�v^����td�Z�?�9�~��^nz/Ƈ��_�W�%������?r��c#W���{r��j+B)G�������nժ�<�m�sO�䑃�{���AH�$�]� �F**�ݰdՆ'�ܙ񦸡���w�l�ehP[k/�4�ߴ۲��ŧ_�k9� Q7��Ƣ��%�(<�`jrȆeȉJ�R���u���k��������U�ʳ�ÌM��L�a�QÖJ�I�	ZI�f{�׾f��+V���uo|zhh$n��-E��FEz�!dRx���W�F��1�����ʜ��v��)s�0� �d�a {ۓ���B��q�A��(p2l�UCV,�B&Se e)bW�;����y-I��w-�.���Ò���Ð���k�������G"+[){�۷�,�t�3�BۡZ�T+NgS]O��r�1���=�P�g�0��?�9� -x��D]ăg��9w��e/�sX����+�[]!@�c�afؘ�,^N�|�3�#�M�o�mƹ���hT��g�8�p�ƪ��enz�g�³_��/�*-�tMI�G�|l��p�koo�?�r���.D`��A�*b���Ũ��3�L����`�nCrNrn�o�,�K5�����&�$H�~��57�x�[�p��Q��s�JR�Y�*U�i~<P�'B,DʔC?[UM��i��K�������'E�S�-~A��+B�߷g�{�)J<���GQM�8���٤:�$���n�����OW�� ����ޞ~����?*b����8�l�l4bcc��7���s/F'��P��O0�/R�q�.:y��a�È�Oҋ��P�,�����);�c�2�fx����6^I�2y�LIvuD����΀�ҟ�g��za�%���Cq]���j���Ohjb�����������Ju�˯��pumC̵�^Y#}���7���������G�n�9�Ͱ�颀����t�²_����t?��]�ӻ;��B�2	H����%�}�5�:����"�'0'm��󥆥�Φ@�gc��Mn�����Cn��ml���y�kr�W����ӫ?�����_�`�u��\0��P�e��̌$t�}��s8"�[�M�U��@�$6`��]z�%��k�'�	�Z��W�76 9�8�ћnH�l��ᔭ1�F��v��>�XH7�̂�u@���"6�,H�4m������'݁SG� Mpp�9��Uʀ���̃q�JB%f�v���[k���&l�� �Z��I�U�B�&6�j�R!����I��'c��u���>�
�Od5�`�.M�3F�j��};�MA
U+�W�"��%�z7]�%��oW_s=mqT�V&:bC{�ңބ��z��I,�HF?�5�S�O��,���!���atXZ�F)V��?�d[!6�Eې��͛6�]O?m�N�b!n�I�����J�K�-qW]u׫+O��P�k`L���!�fj+�*^���hXͼ�2▻p�9ј)��%	̽Ú�X�x)�Q����Z)4�(��������:]�Ϯk��� cW �^�g��Q�
69�o�;}��A�e�㱅�����2t=Ki��2�@b�ܣϕ�Wq�#�-�ϠP7�L�r�����o��z�4Kޕ��nيu��/uQ�t/ ���S��>s�	�E)O_�S���l�b 7x�:_f�� ��̪KD���J��ʲt#�!�Ęߞ1��.>%�����3�&F�MHX����ՏGD�8�������}��g?������������7�qG���p�����WvF=ĩ�[��?��Iff��s�:+���f$؂�`QB\�&Uk{��\;6�����֘�JO+$��z�xϜ���<���������Z{{�s���Ī3S��%��Gv�v%�l7�lݽ�n떍dq�_��7^�撫�8�)-i�?���]��#^+V���v��j�26�Ԓy��]�k?P�d_���%��c�&[Ԧ�t�|�r�:d!���b��m��(�
bCGS�Rc9e��!秮�� {����P�>��E�s���y	ph	 �h�`鬬`Wz��ƕ\�:�$b��!���S�l�	�l��2Cm���X�1T$Ƌ韖�څ�˙��^��ANE���8B Q�Za�s\=�i+*R�a�zW�W�Ӧ^� K��8F
p'�1M���d/��� ����b�Bglk���2\M%���/)(2�^�ƪ,!���h2I�_v���u��h�?Eϻ`ꭇ�ϻ�">S����c[P�Ҿ��[�)�q�"x*��nΜ�yl
�|�����R��{�Z���X�T�4�g�JR
*4I/����1� ��H��Y�&jFW}����4R7!YX��+ �2O]o)�I:7���[�w���M]:θ!'(äӞ�V��Z�j5�q��L�F��!��Œe3���*���q���7¹�2g=>	Z��>	C��w����
��?w��꬛��B�]��4����9�q.�S��v]Cb��R�����ɑT�󓮮+-�����#�Z2�5��π$�c5�R�1�X���͊����dK�͡a�(���e0wa�%�G���rd��;��ul��<Z\t��ӳJ��;������	�_�ܻ��o�[_GKڕ����׽mm[K�MO<��W����#^r��Ȼ�?ւ�r��C�N�^kt��\�Z��Ԏ�F+|)��9��t������tD�I�u)�ֶj�U�s(J-(r�E����=��_��~>�^��;f\��{����]}N�BcK�}(����!��O~���3��#������#׆��I�dM�.Y�A�d,�5Ļk���}%B(�&٪~����Z���W&��BܥG?DF��޲&AӼW$�(�2���E̳�Ȯ��>�R�Vk��ӷ�x5�abS&��|���sn�۹( �I�>�c���W����R��(H^����©�kZ�%.Aa.�6U���(.]0����q�lCD6�Z�WWS�ڝXk5����4�T6�eb*8|��d~�	WR.����*�l�	g�����ۥ���[��*�=*i�$k�8���8�p��-(Z0�9Ml�_$���B?�9{���
�>�i`�^��C_�Aj<k=�����C\g��u��&�U�.ް�6�&��v�IfwT��ƪ�R�H��_��j�֞�o�ץK#�򁂭(~���j�k<yz����@@��������!�q�J�]HN;�zߢ�bw�5׀�@��|w�P8\yi��8������n�"��ġs�)����kv�cfKP���l�05�-Z!sZhF;���fj9�A����MF����}<A��W���+]&���4�\@^$�H&�:4�(��)Z�rE��-��X����W�v��V��(���|),ٽɀ`��K�=�u�$r�<���P��>o��mYϔ�
X�u,�,�97w�!�T�hN������u�A�����Vf)���슅���;���͏|sOn�ү��������}��װ�K�uU�?���_�7�����r/����A���������l��k�����C��N�_.(������m��M���O��g�P+�nF�;>>&�<6g�^&1My{D�Y�2>�Yٱ.1=�54t�};�����W$��OV����ܚ�7��h�������l�޺e�#�K�E����%��w��ߛ���uw=������S�-?��Tu�0�Y�d5TBY�Rpն����q�&�&!��Nً�8/$Ҍ|)�#�y��-]������y�z�\M��,!`X���90�i�+�b��j��@�׫,b��P�#��\�1��^�"�R
k�zrs������_�
�k�6'�ř�W�Q��.�,VNxȻ���Zl�+1Ȋ%��Y�4���l�	��^���Ń y7�=MvdY�`utQ����N�C��KC�:����S]dE��HLA���2P�
M[���/--;�S�`\��gq����@A�\��T�D��6R����@��U��m[ATM�fFӾ@:�70��J2�+b����W�x\���o�t���o4Q�S��p\�2cq���?�g"&.ړ���Δ*�ʞA��K����=u��r�:�~�Z��]@$�_��Q��҃J�{457Z�~%�yS|T�؂�w���TA�܊��,��Dw��h?-{Ed�)^p��b��8`O:R����oS����� w�J�,���>�[�9�6����`�:2|e�.� �R��LpL���a��5�< 2�n��IF�N���x�(M���s(�h
��� l��"IٚQ���vô.�
$0f8.��^��6J"��&@��m:�J��Ir�ӱ�"Rs��·"� rtq� H�=J��郝.�h�-ʋr�9��c���7����>�-'}�73�?������_��;����_�ٴ遫������y�<�{wf,��v�"�R�̆�'n����"����8>oɩ)��ko���p�̑R>�-lYSC�݋�:ko��,��rmVJi��͖�.Y��'��c�Y3dG�;l���#T-7cl��d%��8�ĝ=���>y�嗥��V��S����͋MX������]|�{��G��O
N�ӑY���ӝ��Hn�����`~\B�+�.����e� gɊ�!bQI:�qj��c.�9`9m\��l��K�cM8�Ѧ����^�_�d��T�p*�vtt���^ޱm;�Ӡ[�v�9[e���-���,��u��ɬ]���%B2�Lr ��l���L���l'��MX+�� �ƀ*�QW���FU_5o�Y]���F���B�|&7,�V)e��m]�|����5��1xDY0G�XS��{a��!��H{j�Jh��6�@ "�0��$�bR�!ed���:��M b�=]���|wwo��h' ��^x8��9�Q�K�D����<���d�aԨ�V��/2F�NA�j���#�`�r/��4��NLc�VvJF��ꫯ��}���."�P	�D�iF�8�m� G���0D��Hsk�&ƥ�|���~^f�B]W�$�9�dXY�z��Y`H��Eف:�$�%s߉"܂�r�t8�CA��ŋ\�T�oe,���F��ѓ�kωd�ɐ�4+]Nۺ��m��M�(�m��Pao��#@R4�ƨd����P{�^z��L,�]��@B�t�"4W���mߺ���G�Z�2�U]���a�@�(�aD���� ]
�En��H�����'=(�8����p4����^4(z��G�RK2��i��H�;�3@:�鎜�sM��n���(F�Yh"8#+�N.!�����&]W[�kjtK�ʸ6��8ǰ�Adz�6vo���ޣ�7�}I麯d�>k9?��h\r���;�J"(۾f��z!^�'Ž���_�e�c�2���|�
ϝ=���|:/ RJ ���|�&ah�����}����Ry�&��C�`>A��ԪlSP�^���Ѐ���y)�ͅ		�@�8��(ǡC�C֐���N��CU�hm��⢺�e�H���bm&�����[iCr%�.%#�M:e�˛�F�w�8���M �N��}�i{rr�7f��>�pdth:|������Ύ�\�5o2�j�M(�Փ}h�GO���<U�l��e���Ȉ�c�!Xjc}����[޶h�����^d�q_��W�<���e�-Mlʌ3e"�j��V�Z5��z���Fe�p-l��l�<�"�[�r-2��l�"�!E:9v�4Y�2�X6d��ώ!�E�7��I}zH���櫹�#Ԯ}z���Ӭ��3��DLnŭ.ָm.RI{�^�Ong���F$I�k��N,�x)�ȔU���C���Y�7�Mo,�X
s���`N0�������Yg�i�[t��T�%�&��+�%_b|1��OA�z��F��'��7�L]6B�n�F ����ס����(����N�֤���X5�z��)�`������!w@�ȁ�x��8)x(X�Y}��M(*̵Z�A�|^jkι�ɀ{�V�*m��J3_�	|��D��w�k_��'����&�&���yb��1�F�5+�)l�P�骫��41Ba �3��_L@���02w�aB�p�;�ow��nős!Gk=򳁬5Uσh?����׾��:�OT�R �{�v�|�*(��x��/B���M�k��3�	.���������`?�'�[��@�z="3��DGO���:t��H�}1M�ƖA:���p�������Eb���ݮ�R_O�\��k�9�B������~���X)/)�`'�s����8՜���++W_��纏��'�����}�����q��u��5_�C]����P���������G�|���+�"DP�&6����P�K5G��Q�
%rG�305+e"�T����  ��|��lSTW���6Ć���z �u;t�]WC7N<��2�Y-�(���j#�5O0B[�7~�ы�1��LS�;r:b'KM+fu(}�ͼl��\�h��ajwm��&�t�U<�(��	�����g��Ǩ��#xiZ��
)��t�v�s� Si���i�bA۹����5/�d=5X�aC2��'Ds�m�Z���sh�C5�+_�~}߲v�V'Po�0��/�����Y��,��-��9�Zo���ih۱^16��M��YԎg�d�^|�!�M9�{1��i�z�+��H��$%5�������Z��y^�q�4��z3r��`t��֮,D���D�eV�TǺ`s�� �xMY+ELFٓ1�Ն%8����Ҩ�Z�m&�vFf60)Y�J�z�^�ޘ��)��L�Z=A� �ehp���v`@ !�E�3]s�զWn'��Cޫ�;i����� ��:K�^�'	Y���|+�%��'�igj1S	@��Ns�5%MP�6jc��r�L�s���O��qWn@DDɤ�� �T�U4��W�
��#��ɡ�\�Z[p<ǁ~{���9�æu���^�4��׬^E0G��^��J���2F@��{��L�G$J/��z�,��������G�@�+�P����&u��_����y�,%p���t��w ն��Q.\�W몘��7����b�|w��K,�P�!4/LL~��Q����L� �Y�dEz�G��8�v�ޅCU���S�BCb�Q�%�N��.��r�,Pv1��X�a��.Z��8>�񴴍���"&2_|�<h׳�r��5�.��b��P����<:f�A��H�],ǈOF�&���a�P��Y��u���??�\Չ�ttt����L|����u����r�C-�2}��#��ط�.6�
1��9�#� r��"�)-�[�����I�ˠU��G���'F�qb�b92�Qw�m�n�"k8���}�Lc{�2�1�:1�����
D���b�Y,+��W*j��٬s����+֪T�T�D�"չ�o��Kأ�,�Õ�C������#��D]�Q���tC]>#>9JB!$83��bg�Fp�2���ػ� |�[��]i������`�md-�1����%���p{�S�~pނeV�OMI�ԧ?2���z��Da���Heg�״-i�J�K����q]���ST}Z�����^��[��C[����L��H��uZ@�q��8����箼��Z+�^�@��tΫW�pgO�5�Ia�L�@Ȧip��x\kl�` �9��P0�m�K' �'����Y�V�b�
��]%�����ud��:��M|�zҥ2�|�[�Q�e�7	������VZ�$$8�)@$Hm`�@��#d��7F���r�x���Ycb���.�+�̆i�m-G(B�r&Pb��!>�s�;
����.j�\W������Ok\z
ҭ:O���	*ĝ��Y��ZE�T�,��	��q.�4� �d�B��Ń���閸"#�@;F{63���M.�,X�s��� ��ӕ�6�G�3j�SO���Cױt^�u�3�9�0��5�}����"����P����P���[�d�j��M5�n��͊J��'�F6���%�S�r���Ud�#--�&��Z8E�f��}�u�A�k�s#H"�R-"���N�Ռ�Û�+n��1�Es�&�P)E	�r�@$��x:�@ú+R�u���>��!;�f��I��F�����������J:f\EI�4��k?�Za�G��X�/.y���4N�\�ڸ�g'��X?:>r=���i$�� N�op^��w�/�h/��<����l`�4�g��Ѻ���t��#�DJ���D�X➓�%!�2�G�رk�k���{����+$<d�_��ށ�����nɊ�]�;�OC&���a�t�y�|xn���&����â�a�e��$'qp��H��F�t���A�`���~��s�u�(wQj1L�^��S��h�a�f)�',�Κ��#[�6�|nh���t6�Pv9����'��1�#	��f�cLhyw�ӻiGj�}�YS�~+�	���ڹ�����G����k�A�}�{��V� �HTe�%���צ��A
h=L�2���Ym�Rg����1͆a�;N���a��0��y�^�}'��4����æ�I�L��� TЛ��7�	ў-d�2]}�EȽr����Q&�9�HU�~�CLi�ŇPcך�� nal����1��>��j!�8QL_���bc2��TcV*��U�����L�׽G�6%9�l�>������'$�`0NJp"R)�V3p��5��M�,Ip���`�^B�<���0����@':�}�W�(��P��������|z|���<�N>��R��V��;in�e����ct{O��#�v��S\cu����n�2N�z�R 0�(�}��E�$�X5v-S득�\�d�GA�юVGy�Sy��/���~�{��]y�e6o^���/�>���.v۷<iA��7��;(�P0/1�q�Fdf������%O���!(�+��2~!B-D�����@�']�)*���
4�m%�p ���¸>E9��V�1�`�9ڽD�	"�֣�PdL�Cc���z}��iv�MOŹ4�G�xCA� �����Gۂ�g���#�E}��CT`�����A���2�P�3��w�wԻ^_������z�b��|�Y>4�����Lb5oB�4�(m�Q��^��������5g��ml�Ogg�-G(�b�6A��44�P��P����%�C��8�{-ā^��A������k��|��7���>��k��������񋂃z݉�Ud˽0�3]v.-=8����q�/�Ť��*(��X��M��Q'���t��)�G�=�Ç6��jg�I5D9?1�ɸ��!���Z.�:��};]��Z|J+�)����3��3U�c���^��]�N|(^R�t���Vy�x����T4db�[���ڠ� ��!�b���ɩkMV� C�����.�{5
m�0�Q��އ�>d�����z��R��\��>���.��K�a��:z����M������h�"����G�G�����ՀEn���Y�(����[��C��Ѡ:��8�d��	aBi���NW�s�t8�!:�@ϴ�t�2A��Q������_-�ƨt�{x��1cVOr����-���s8�t^-�-z!1�3��q�Eϱ�(�5Y_x$�\�dʥ��k������j
���Q����---�8:����V��(u�fF�K��3\�6J��"	�P���l�q�l��/]�i;,]�r[4�ROcY�{i�JB����ئ�®��P�@h��� I��>7H	A⼺�:(� I�O`��:��8Ъ�=q�du���Rr�v�8���@2"�?�8�f�+���R��	���Ms	$�j���1�p�lK�(�ϩ��Ck6�$�m���fy��}�ƍ�h���G�BB7����u���$U�U�"H���P"MG\�p�Aa{�Be�ϟZ�/�GQH�Ę�Gr�iv���j1�>�lU@E�È:*���K�D#�v;#���T�����Xj|}���]�I���(Pf�D2f����#��]��t�L7ܳ�+�?�28�~z6L4�|�#Z��Л��#/�����X�%��]�6]s���ޱy�q�d��3P�c�c5��(�v���`w���������=��vn����c�0��z��0 �T}��_�m������ѳ�j�����ޫzz�]nz2p�<`|M����#QC�b�Ȧ��!F[�e��=�:�|�wW�[���60�1�B�]�*�h�9S�����}���d�{����Yj_l�S�ZLsy��ʝ���#'����=��������Vl��M�m2���|��׼f�FW[uh����]�B"#)/[�V���a�P,���g�5٫�b�#b��q6N�����шo�������C� ��MRcD�^������t�
AWf�"���"p��զ�nٲRW�/L*Vb.�P�e��׭�����o���-g��´*y8�+Y����X����v;w�v;r҅��!��X����fC���L�(��X�A�>��K��CQ��QT�"�S�Aui�U��I��l�&:k�+V4'��	�������	-K�$#(ٜ��Ky�~r�G�rO��7 |;e�^(_$���/�����lqW��)�Q$5��U�
f�~

�Ⲏ!��xg�I�:����Rz�.�J�2�����6x��z�ʹsE�zzc�I�J�A�dhf���CGЗo��U������a#^	2����n�����OX��O1�OQޤ�#��E�W��AY��"��!J���O_�
mF�? �fbR2:�٬�%ߪ�K�􂮈jd���� ɚ�Z���= @�����������`�Dk�A�)$*���.�mt`�=�c�+V��G3�ǤУUk]n�BW�l�:Zd�Z6�wB�A���������S��ߛ��J!��R���;�MPd4sBR?� �v�-rsk���bHw����Oq���&�)�t�_��mގ:!�م����ǪeSbM�([��F�[��i~��]�����/��<S}|!/�_�Ҳ����OO���}&?`VeJ*Y��=de�X�b�=�����程��؇�������V8th߂cލ���`dǧǫ/����Ȍg���wtuly���9W}���8WQ����F+����K;��PנvI�GBd�cHI������+��c�k��׭���i,�������R�Y)��4����"���=9ed m* f~��a�:�zZp�c�t��u�Ό�)���͇2�Zڸ{�7�������2�N���G�6e�8ߞ�6ڦZ�����6)��	6<�)s�G�G�i ^����ѕ�&�ҥ���E�d.�$�g�u����Fft��6#��"�Ik[�0�g�X��;��u�����FIz��x��wt����N�T*QK�{�ٗ-_�©�[Ϻ��T6��(J�u��''�Aˮ����a�+��N箻fZ濾gmF��=��Dn2S�n��Z�x��U:1>� �Vj���Q�U�*�^WiA"<��?��C��o����\�4,��j�R��n
�]�-�Ps/��i�f�'��m��:&Y9 �L=�r`r������_�Ap1A�}��� 2�@[d$���>�P�!��/(q�q�Q�g*�$�yM��CJ������f.8ރ�{��mۆ@�*���,���c��ٰ�R��Ǜ���mLw�HtSj���=��F���{3�L��c�v�N����u,Gie
V'�:��뺌�%�c�Nw�H%�|�TSk�����ƶU�R� � \�z�s�=A	B$F�L��C;lT�JK�+b��^w���&H�^xoR��p{�Q�!!U��zz�e��l~�@k�����ܘ\��k2̵��c6{l�}?O� �����w��y�[�����_�����w�zw�5]r4o�>4�}90Jko�/	���u ���ƪ@���~�%Eѱ�Y�������{�>�m��_0Qi��%ԏb�����ar���+֬{CRbZK}u�'�S�W^q�����t���w��[;����7R���?�Ɛ)jw��p^�}�K΢�#�H=��6F'Me��Ad���d�oi9�
sť�8�f�X�͆��N�J<p�Ť,��V��_���s}e.�*��p���Q8�j�idZ6��8{�M~��8���`���cd�!��dZ-<.>�-[:��mF���-�p��O���I��Gf���ڧMQ� �����%f�`긖=k�V�-g�=��b�۹/-V���� �z��b ��8P��T���%��T�ΦmY]�H'����$�"u�0��P6���FǓI��M��C��Y	�z0�µd4-^ʴ3��U��lq�qz=`\kzo��G��t4xE&A�%�-^� ��،��չ��A�
bнA�^��*��ګ�z�i��,A
W�W��1A��D�G;S'��>��r]�ԅ(�B�JHN'HR���\��{b1�#� �I\gI�fge�Ƹ�肓�D�.Ț����z�"��~�C���x������J���hW1��Z6�ü�@ټy�^����Yٹz����i=��Π��?$9i$�Jr��A�*�������KN�=�$�3@p�Ut&���ߕs�	m�s4^��U3r��}�Aw��K�Vx|�|�*������^���j���$�o��q��*��W�ln�U��	zҶ��\-�[���-?/��5��߷=���x�iGH�(7�@�R�V˘ȳ�(ȵ�>� @뿖�Z��m6S���h���A0gkj��Iz�H+��aݺ�t9� h����'C�����"<���=�S�:m<k��|�ݫs?[�2�wi\(k�������~2��L�fĒmÔ��u�..s�|F�j+Q����pjZ�B ���.e>
�|>GF��ID�:
���4��y��p�^�3ך}��R���y]s��<����+/o{ϻ�}IMM�ͻw���n0�l G�>QQ���+�х����[�ӹ��Q�G�b"&��ָ8�Ђ�z]�iX�r�2ܚK4R��#�%x�����������yFٺFrN��M©7Rk�qk�Ż{�ww���+�1}k&ޝ�샼���6H�#�b�I�1*��!�Q+k�k��IF�Af:b�iu�T"Q����"D8�N��O�X�jv� ��S�z]�0�W�!# �)�wfp���>��m�\g�F�m�Sn�a�`p��om8���7��c��"��t��s�]�47��O�~��#8.T�x�`h���ę䨮��AF���q$v�Z���E6T��i�pA�V���s�j�i�1>�Iw��1��S��qΫ4&u��=����ޏ��97�}�
�?g����b��	^�L,|68��ջ�l�X�&��Rٜu0���g�M-�l���M�d=��N� ����n�� ����+'����@{<��hÆ˸w
9Q+�PV!!ѐ�:@�q�gN]Y���j�HBb�i���~�D/���B�0d�j�|�tb��m޸�˭Ϙ{{g{�;t�4]�Aފ>a�;�x��I�Ku�� @�o1��K%O���©���B$/�`G?�V�/[��~@�WkJ��u��=�� IF=��"�$�0)��T�Ѐ�2N�(��fɫD!�9����1���mu��0�N�1<A�I��(e�x�)~"�f$*��@�(�1��}Q~N~�yNN�{�ow���%~��
8C�RSS�v��d��M?�u�^˪�xv-�Š�;/��M�2s�ۻ����~���ύ^�	J4�wA�,O��p���<�`�G�2��H�	��t���>l�OI��>�~3��G\:�f��xh�>�8o���g=�w�/�r/�ם8u0�3���}էO]�����P�Q�./_xO[K�?�WWU�C���|��G�8����<,,ZX��>�|�{�65~�5��uFF63ʴ��JT�B��3��D��P�2�`�~F�t-s�$-�07�0c��e�3@��탮 7��vS3�r�H����x����Ϲ�E�0�sȜ%��#cs�Լe޻���՝�&k
��]Fm�l m� �8=����,uR4�3�IQ�h	pv�m(������������Ǫܹ�4>�r8�lL��-��[��$M�lWcA�V�66J�NR���(��%q�L�Ӯe�2���?pn����uk)C���F`0�����]�k��<:�8l3✆!�L�tD#�:<D��,[ٿ`�AI��1mmj���s8��;ȶX�7���g��I���A�|���ʽ��]���,V-[�@���M��=c�� �U��p� �I�����B�v��>U{��΢v:����\e~�Z(�R�"���sǀ���=�/|[����$c�?��	���>�%WوX�w�K7\w3�7�6�=`K�:j��l"ύ���%�H�f���Vo�܁���?e���=(��T�+�U�pO2}Ӧ-�7y�Ɠ ������+���ǎA�Z��2��j�ش���]�~=�L�PoG�L�1����H7_�����P�u`�s���n-n\Ljx$��H���:!ds3�1�$�L\��v젃c��y���l[��G�s����]A~��":�Y��'2��U݁�+��8���P]w��`���~SˡM�#�b��}�ŕHM�0)a"l��H|^��=]WI�c^H�lV��3�^�V̃����s�޽��]�~��7��u���ɦqT_jS�C�������n�\<-z�.$�
ؽ�e�`列B�\�vLp��K6��e?��@,D���S��P�@2��}/Խ���Z��o�g�G>�/�tU�b�&8�-��R{��R��҇�#��4�qF������\�����d���E%�>�g�\�ظ�}1�^�֌�c�;��5�K������a
R$S�(�㩍���E�l�Fǲ���aġB�k��<m�s.��rw�|jSdN���n�a���{z\WK�;=8��Z����-ES�	�禁��ج��y)d��:�&
��C߶'�.V�v*�h!跧e����cbX/����>�梿�I��Ը�p͝��`v�B�Kc(o��&�<
z���]�� ���fu����2yo	�dh���]Q� ��l�~��C��!U]J���j����ƍ��R�FJv��t���;{ص�4�]�nCУtJg:m@��_ɏ����WU��lg,m%S޳&d�sgTFɢ���}套{��m~������0�0�C�i=���Q'1^UٗA�,i�zŗcUǐm�V���,ra
t�h�, ��&�yB�Ab(hp��(*oj荵[Q��8Nl� N��
�/�2�"�`Y9���l���k4�[0vTC/�ؚe.��i�cux�i�/�C"���Z�g-_������D #Mt���G��kF}�H�8�9�}9��y��������i��u�"�]D}<��3g\5���2�O �_�6ɐ�.����n�Ok�
Lx�0��CN4�6@���AK�2���[����MH����P&���,���}��}����3m���������<8&������G]���&�� G3('�,�-\��eej��d�
�<[ ����h�x
Q0g텳�YDDv��l/Ӷ��>�^h.7�m�}nF��6ϔ��+��Ӻ0H����eWH��F����W�L+]{�V�/��E0�}���~���Ƶ����v� 9�N5ŵ��vO�CW�0r���;��?������/x�۷m�'�]�u�㯭�<�����BZ��pt8ؽ���s��ˮ��m�?61)�L�)��`�JF3�h�fm�wD��<H�չ�����������S5��zse�k�끬D�V!#*!�x\�W��o�q���W�Li61p������ձ<�� E��&;Ipg22����1�&`ͪn�J���K6�B&�  ̽�-��:��#�v�sf�KQQ�#I���Mde��yG74Ny�������[��D�Vw�Y ��N��4$&K\[w��ٽg���]�������Rw���Y�^�e���� ��;vj(�9z�� eͥE���/s98��m�� BeB��j#�V���8ۂU��N�N0v=y�;u��������s��n��6�����2������J��v1����N05˜�A�F�K#2-�!`�u���S��[�z���%H�LT��R�"�*�����I��|Wq���#�"�y�n����dL��f/��r���`�Ϩ���6EFy��	����7r�9Qs쪩�!���|����Y����)���OD/e�se #�)P������!�شy��BDDm��{L,H
;�F�.[�����JH��&�i���<l�Aj4�@��j�*C&�::�.~7�|3�+�!"B��Q��
0I��Z��L[!A��爺`�AP���&�$FJ�{퍥��kt�j�vO#��|�f�3o���LKa�([%"OH*�s~��@���� �����6o�P͞�7���Ь7�y�#�)GO�ρ4��T)��(X��$*h�_A��\�s��x�Kd�Y��]+��+��e�s-�s�U�>�g?��M%���軵(�}n��׈��{SB�OAz�3u/�u���<H{d �݂Z	:+�/��)`��n�B,��O{�p|��Y��Tp���1�v�O�Y��������;�?�Z�sw�����'���0�`!G��5�k]�`�z6�^�����Η�S��W��(�Sd��ԞՊ��&�@���F��IkX��`K\��0��-�#o�C����� v_׵�ff��Y�زe�l�h�ph^�~��5ezm��5Imp�1�$˖,f�i�33}��Ͻ��8m��׾�7U-�\���?g��k��bS����Ǔ�"��Q��M7;�Z'����h&��%����eE�� ��I�U=�6&���R�&	\��֛#کk�{*@���깑���>�1W��o���ظ�,�c_�+�ִDj�v��"�\.?�\3��ñX\R����r��]��"Y�N}e���<�����=���5C�is��O� �ÇZ���9�H\b�>���b��Q�X��u� ��K��5��Z��3�ZKJ�]O�j�'�|�H]=8���b0���4�q�`��h�n^�������Ы����U\�vW.�}���.��`+�Z���ߋ��<���r6g�Q�x�!������؄�j9�(�Ht"��E�3�]вT�T�V��[
N�ى���φ�C��.w#Cj6��"}��k)�ҝ�&x&n��.2�����p��x�����0Ї�O_���XS���o���"9>1��E�=��5�eH�E٫j�-��.�8�w��7d���{qY�d���}⩟C��0�\�\�Kv"��N��S	t6�u+����rB"D2��^qg51M�K�c�e��t0!��?w��c��Co( 	[���I/�2���mE���hO����	� Z[���Ip��	��p�չ�{"��h�ǣ��µV�;�^E׾W����8t��� *+�yyW=��o�#\���G�&�Ǔu�u���vD�+��B���Qj���6�/�D�51}9�'}�xH��V��b6�or��"52��^nA�b��:�_�����l���v���z ��]K�k@v7��ժ�xt/�@*zIx&�����=�b�Ϣr�Fi��z���]��'�C<��[���9@�ޡ� &f���9������w���r��_Wy�<u��7��mD=��v��h�rІr��2�IB�h���Z��3(���ԏ㨫"��j���cD���*/'�Mʏt�&���D�BR�pgN�3�0���b�R�4p���[jd�����Dr��n� ���,�O�7����nR�WB�800G�S,;.��?R���!QV!m�=��9w�]3����O�l��6��Ux6F]�� �PF�R����g��Q/�"-p�eY�9�3�P��� l�>���L��biq�c.�0��"����k�%n���o��|��m�T�V����3.6A�7��W[�&]X�#á�%�a�8�ԙ\-ףo-��>dK%/z��	c�+�52��d` qx���c�ӓS,;�g��%WVrUm��S�����^�^
�qd�Y�Dc���Gy����F�9E�S���uw0�^(	�x�eҒڴѨ�cr�+�k?I��C]#X3`�+�Q��r��*x��"b�PWW�6m~� 1	�
�<r��W�ENǌ�꽬��R�n��j�/ˠ�@ 	Ƚ�J��iZg�iB\2�*�eC䚠v�5���y�koF��_���{/p��P'�VE`����h����^|���S���y�qIJJ��h���f�� ��ӧ�|��IIP~�#���ា��AMٟ�¥�F�/*at��r��fh�sH�|�Z?�����А�1��ם��#�ﶿ���j����`IA�EV�������2͏�Q_T���lonqG!=V�c�T����"��b�����@���?V��㑢$�R���H�_׮���8f~����n���0�����&���㝫2o��1�cp%,I�Fb_��!Ï8qC�<��~oA����{_���g��ɫjiq�l��V7B������oS)єp�[�^$J D�e�m���S.-��/j�6hh�$�b_��)�b/�=��T��x7������E��y���K.�����U��ܵmm_��y�ې�[/�!'�Yr�m�2ѡ�T��椞F]��7vmq�[��\p|������[�^{��M��\:��O�u����Ij�m=nΌ<j��@%��1ň�q�9��4R�!�� 14Ĺ�A�6� �\�;��z���|U.�,#(�:.-�u)E�Բ)(��L�B�;y��e4��Q^�L01AV˟�g�X�F�����Ec������+���
�r���+���
tp��/�]*o��V�ZfZ�wJ�]ii�K�A�Q���N���8c��0�|���\2�E�-3мf}�7 6r��XmT:�&�*UB4���*��_$�����7�v�,^Y� ��/e2!�1z�\7�XoG��x�Fm�GX�����Of���� �I�;�f�{�|\8ʥ+���5Ü�~9���`L2%�RAD�#��ڼ�
o2�bEo۾��c�lPI||�� 1R�b���n��un�2Doа���Pc1O�<�ʘKe��cFZٞ��*��(�dT����6���?e�:���ŧ��Yf.aZe��E׍������g�~��E����@��P�J��sѯ_Af�Y岻Z9�Bƛ9|�&���]e&�Q�.�ѰҞ�"6Q���-VZte��n�̩n&d@��u_UҲ����p|�p���K�ٽ{�B�Í&��祿7�u�O0�vG9[�A�@���]�/O�Z��J��R�%']}�[�C��?.�.�����{���p�*�(��ԯP'�)T)b����A9:U������T���,b=%rd] �?j�����H�+��'��6v�-HZ�.�^x��C/ ]��N:�=����v�yqn|Xۛև=lk#���B"�Z�\HE|"âط�@�Ӯ��}aDN�XJ���(�Gib��&�A*AF�,i�BP�B���շ���=�u��<�/x���1��念�W??0ؗe�_z��5����Dm:�Qj�"����6mP�0��-�n��i�j.��om����sŹ��*�<����K�a�m@�U���Q�̟d��aj�ʪ��~��^\��P�V�u�e�r�4�	�����Z��ܔ���>����@�I��1�����Q�ط�>��6cN�{�*�;�.��펖0t��eO�Cd*
l
Z��$?�r���Bzȩ�FXw8���!W�8�ju�p�����;1E���g:F�kx4��=Hgf���}2\?"8�-�h@��dd���QAC.�y5=��m-d���5�3�L���-���Lf�<��VA;�)2E��8e��Mp�D��QX�ci�<O߄�H��ǥ��e�����p5�WI��F���[��'M)3�[��9u1|1�R�Ӕ<M�SmYs��T�L{x���W"E��#>�0��j��t��iڋhH(�+7��� ��=�����\�7�.]�$�*�+�~U� g}�;�f�T/�ae���mJٻ�FU�U�1f�	�ԇ/Ov��W����(_{�UZ��]�<�aJ�8e�� %�ܩ��vk7�I;Y����2��&w��	���͚�����ꂼ��P�3�-fmJ�Z���c��!���'_b��H��j�[[������s�n֞�LV!;Q0�ɣǎ �s�҇��V-���f��[�݁�C��'e�H�,"r����/�?���l!6�\'�u�ED(AJ��F���묈2�ϕ�$;w�a��Z0JGI��'|�m۶�u�ns�i�Sߟ�Q�����n�C�q�"��os
I��N� $RB���_+ �����7������ٹᏈ�
�2�sL�9�+U��fڐ%&q�Y	���5Q9��%q	���(�7����[�Ї�8t_����=?s����u���g|��};?��_z�s�qN�i��v���WT��*�8�N�c�۾��_�Dll\���HJsG����G�ĕ1��6)����P�j����xɂe�u�sG�v7l.l�o�a+i��X1�,�� �Q��a�z���$�t���D5�%�&��YEL�qO��Pf�[B�<=��E+�㼍�g����u���ъx���u�|����.B����v�[rK��N@��#S)"��Z�:���Pv�=k[��)��:�[A���C��u/���!����ő�3���#�X9�Nb���K�qќR����c]s[A�cD�>FH����J����+W�(J��
!\�L_jr�gMw���JR4��T-[M�<Z�_�G`26�~�_����dcqƙ�����9Y����TI�xj��3}	�'Bv#�#v�g��!RS�d�>H s��^k-R��EޓCW���ٳݴ�L����I�������t�[%z��]�<B��E��{��H{!�i�O����tOo��[I�=c�G��[Y�e�2���d�3�LE���
�`��Rx	��}�|����W�v@}m��.�DZ��|�P[J]8�sǎ�B.�Ե�����6�9�V�K^�c��(R\s�c���
]&0���c�|qI��+�=�b7��ȌR�7!��yL��l�\omc��#/"VQ��h�!^R�ܳQH��̵��Q�ˣ�K�x"�	�^�b5��ɔlЌg�z�(m��Ok���,[J���������#	�DN�]�t7��/ں�z�񽒎�@wx�~[*=		�6H�|ݛ�e�W;ڰ�>��INKv�<���t��;r� ����~_����Ө�ϵ9�F��Y���88Ahݔ���u�}�g�w
�� ��`O�:��r�#϶Ѵ�ؾ�sf�E�#��Tf�����?K@�C)9����@�g]BK}a��,>�������������}�w_��}Ο;9�ȡ�ߡ��R���98j�	��?F�O=�2t�
�E����O���~�o���-�p8w��O���\3�E'�h��7{ɝ��y�>=������[����̒ʳq �n�L2ϴ��f�����Q��G��]@ԌMc�`Yk���8k�c�����aH׮�� ���9 &Q��DФ��N�k�k�	aN!5���ӧ�܂(7yj�+��Ϝm�+��]���&i ��1��Quld�w�|9s�c@lM]���@��A����CP|#u�D2�FWy�����l��F@�Ƀћ�{ �
R1�#U�;�v#-j?y�q�:�!f�2h�D<�a	0~�)����*����W�{�� Sa�4]�(�/�/�E60eR����.��{��!W����#}p���l�Ξ�`���G��-Tb�;d�W6or'��]<��:���1�,l1�\��,_���F�u?y�Ǵ�]42��Y�m�~쨜�ڧ��&�����܋�0E�"��k�t4��M����*7R�,��Ã}�̝t��ȶ
y�e����f�ʖ>|)���k\:Y�r�X�^�h��Z����o�-�L[�.u��b���I�l3�ii<φ��"T
��]�2l�3n�C-�dA�v5�D��-���ׄ
ym�(���Q�[fA����Hr�cd���Ʒ`_4����cyM��-л�6��z��"��cwS�Y<��n�A����c�����	����m��W�k���m�����i�T]H�T��9����p1�y�Z�Ͽ�,�I�@�+�O�8�Z%%	�)���~��Q�ڣaBM�</��q8�4m��7]~X��� D�Z8�N��R�Y�u�{ ���J�)����*�G�C<��>s�&�͙7O�/6Y�6B�{�0�E�����{T��� i������W�����]B�T~_�mǦX`�*���|�N�]��vW������|WGۇ�'��k��[I�9yʁ��#=�i�Y}����:�.�L�	�������'N�/<v��A*d��A�ݵtŢ���Ew���|W���*�r�A��C����#5��1�#`��LdÂF��O�n�cg����T���2�M+�w�u��{]3��[;a470)m8�w�d�8`�wc(J��F�SN�
�>���!T�T�D��NRCW��UÔ�gO���O��>WA�^�Ft���c; �L�6[�e� �C�%��4&��BC�hq�O]"�rK���Hs��������-_��,2G(���3i�Ё���5'3����������[d|KT2��/���[�XY�"��+k�������j]-uW������ԒR7���DD;Y3���*	�dH!�!-@�d'~�C�Z}��Q���Y�#Ǐ�<�C��V�C=�RS6�+9Xԅ��<��{̙�@�,LFx�޽n��&k��r�=1��,��a^C]z>����e����ӂ����k��3xR�e?PF�Z�ϝB��%��5���8��FUk3
c�(�˱��>�[n��J���b�A�A+`϶].'��g�\�aԓ4��q!d�q���-���>��sף����������~f5w�/�ۣ7m��Zo��Z_)��l)�<� p��ň0-���`�/�M�s{��?u�d%2�[��*9$������М���jZ�P}����f�:rr�U����&Ё� �Ӆ�����&�I�#��$`�	m���15��㢉�5Nr!����;!�A��ǳg���i �J=���W���5Y���?���l���@
��)u�k-��m0�@]��ݘL<�'Nĵ��ϩ���q�P���k�Y���|���Ϝ����J�����g�l�̪I�`pP2���>>VN�w}�� s�.#5fJU#}L \��)f��^���)>��M����绐�/�d��_����ٯ�_��HzJJ�-��]	��*�L^�9%5夜������FV05떳o����y�_����u%��e�FBFJiK��>��ZD1�K|�|����U0�iMw� �-������Ϛa� ����Q��sw��B[U;��]ͥX�5�=O��a�\��QaKH�mM٣z���m���A�2���k�2��$�š��By���Aئ}�c���Z�A��im��0K�h+[K�D!8�s݆�dS�� Z�\nN�1����T�\$�"MsA����>]�0K��6��� �x�B�����ֽd$��#C��N���w�z44���ӡ�0�H@b̬��@�d�h,�nY=>AD_�1���ʹ���IW���RƗ��n�3�65�F(I��?T:c�5� 8D��j�yWQW	' ��*���Gc �y���[o��:���G�yje5VV-|f�����
�j�cHq},\MU���ʢM�#*�|��3�c-cq��8��qX1����Y_�Q}QA�%��)zܹ�g,���W`�{�я��J����B��,~��@��	�1 �#��a�X�&BR,":�$u�Q_+�%=$���!n񊕐�'P隩�����=R3���r����JJ쉊
�s������^�J�k�H���N���բ��=��p�9�ʐ��j�nL�C[_H��g����}L�K�;/b$�}&AzV���'>��>�4D���9.��C���(J�F�ޠ�t��H�Pn�g����N���>m�S]+���] �P�@k����L��"���o9�G�}��o-�r��9��pΞg*�yz-XQ��5�0s�L�|�
���KcA��DVw+X����K/��5�g�ÃY�Y�� �2 ��{[� ����dbҀ�3�=h`Ź��tR	hG��V#��4�ؖd}M"78��"ֽ�@ɡIi)G��e�!A�sCⱕQ}a���srr��N8s}�w��y��K]��w�����[)�7?��?Z�����ؾ�{]�-��5H�[��с���w~����S�)����ҋ?��1���9�	-�iw �a��g���`��XW��kf��o]�q)nߩN������ԵD��ȡ���:�Fs����vB*`��0���S?ه�E�[�2�L6#���!�K�H���2W/��f{E���(���!�����d��"U�ydHiv�I�Auq��|�V.�a�k[��*ejiJ`�a��Ry�uB�)+AtFY0�8�N-�#f��2ܪ��Ȩ�ܿ}����f�mr��G�܁Ih�x���O���w��V���pSi%�ȯ��{�ٟ"DRm�F4~3�{�HF�N�4�7n��C�Ěȁz�%0��e�Ȟ	�B5�s�~j��w��Ɔ��b��z��[�it��|.Yh]}��ڔ�2 ���V�6�.�f�O��|���3~��a^������#KeNB4zCX���*�_�����1.Ck�ez]d��t=��K6����yeek�\������� XL_�\��yh��T)�xZj���L��^�� ��D�H��ǁ"hx����c��tF���m�cv_�N�#��I��)L�S�ۃ"*@PɁ�G?S�5�}�8{�?rNC��B(�{!ڛj��>p/]�o4,V9�LN�ҥ+�E�$��&[�WL4���@T��uR�aUk�,U0o(����w��3�ׯ���	�A���*�I������]t?8pȕ#~�'���Q����͞5Ӥ����BP ��-PW��-C��>^VID�`|F4�{;��
�4K�JZ<YS�,Z�f3���/~�j�Qj�C!P��zS��xm�D���F@g�D�4��@-�1콊ۍ&A�:?dG�v���Wf=�;{�V�!��(!H"KfA`Mf�F�YZ�,��PPeJv�at5h��IX��CQ|�PGK0��\597/�u��.&��O�g<�1<"���o�����������w�;������������g>�F&����H�-�_S[��[6����佝m��my��+�7�ı������0��']����'�'1pq�#��3�w���R'OB��� ������R�V�Fu��Ң��f�rT5�`�f���Aw�]��D��'�=7���fI�HA�"}ԧ��ե���#ٹh4b)w�^%�h+�E*����z�U�0��Ԡ�"ۨ��U/(���4����h�t8,cj�8�q�����qW^U�>4e�N=p���p�+-��@������wgN\��`�tԝ���#m�_?��/��9!�o���@i�6���Ϙ=v�(���AHUY�s����gX��I-��^�����F_�bPd|Fq�$��"L�T�r:9��fM<��K�C�����.w��k�k���bÛ���]]ϨkB�eT��u�P�ZAg�{�+��p���h���я}��\�9�t%�9R��e"�b�� &�r�
&d���ʀ��F���8�8�ku�>d\��ʂ��`(+�S�CY����8B?D�/�U�:���݇!���������nh��9����Q���nɊ�$Y����3r�}����h�����4���SJ�Ai��2Eu��T��IeSm����^������c�Ĝ`l�iDv��$ݩ�-C��2^������o z��m��.:���:�n�a��I�rD${q�0j�&�B�ƼpTm���y�m����'z�4YQ�$�E�k�p\�D�<r�`��������	�ĕ�G
]`/�A`���B`r�l!x!e`�dh�u/	�}�v��Tf�9k��g(p`�ʐ��Լ �W����f������KIH��>oaʆ��P�8�₪l����f���3e�D�kd�G�m�řp��E��̶H�Ɠ����$pu
�	(TJ�&0͂@��=L��Eo�bI���m���H]Y ʹ7�,$���>,hP=��H������A[�H߰K�]-����\�|tEjz��S���c�\��C������G�>}$�k���G��^!�%�r�D�;wl�kld����ΑV���J�2Jm-�9�W�?���6����5E��s��������h��攰�W}���]DM���џ�^��!�I��GEe35�`���8Ǻ�Sc�K���O����|$CG"����x7�1�?ɽ�b�!q(�Ÿ{Β�r���L��2A'?��7��e�z3�0��q!֗>>N_;3�U��"�Q�v��>��2 i�g�Z �E&cDi���n�B���Uz��i�F�q�Z+�BԲ�S�<��/A�YB� �`��Sjh��qSf��M��|�������=J�2�1��M�l�� |/��d4g͜m�[�Ԃ�u�M�� ��S�R���r ![�����94�5ͬ�/頫�/�һ�	�W]�O�mN_����"��h�7��	{a�KO�F�BG�B%+2V���U�6�e��<)9t����!��y�V�L��
A�"z�HNu~^[
���l�Uu{�Z�]1�9�\����j�V��re׎�@e`�2�{>1�V .S��Z��_[[��#�"��z�մY�!Nf|e��Yh���K=$9�uXٞ�h�`�SК4ÿ�fO��%RS"���ݫ�k*_�bj��{IPr��1.w��䍗��aȩ�B^�~�����Y���:�rr����Y�4 �s�v��\&Ǣ��Xe�
�B�,��0���{	���s��B=Wn���� G�釅��������Sj��AJK�p~�D�Q���� 0;�y��o>dFEm��#�R@�鬍[��Ӟ�L�`'��~
�3f����V���8.r��.rY�j�~~�r����ۑ	��7���@�&�6S�N�Y��Jj�&f��n��M%PAl ���F�&�Z�/&{�'�6G#��F��=�{�@Z�d���{-�=VVQ)F�RWh�Q�T����yY�,0�E4I �ĸ��<�v}�ͯס��+����c�s I�����ۻwۧ���>�:2*$M��+A�0�TN۹}��#c�wFS땬�q��GbW�a��'%2���'����r@:#&z�j��ྫྷ����V��D�*�n��ݻ�����d�dڣbӒ���B`c�YzFme�ݷ�y��h���������*\ӕ�Tt�����¢�1]�
=�"�	��\�k��TF��9:
�Ʀ.��Q&�]��R��4ո�24�!����3�6}/P��×Q����wq�!�����LX������9��*�\Gw�����IF�Dg|Db n�T��ūn/8/�ij�$���k_s�t|:Jk��r̲��+��k%��`��XQ�ĩN�Q}����"sb�f��˘���Ր�P�2C�,#�\��kӦ- �=a~�2����F�j
֏j�f��rw;3�� E�0ż[Dm&�����}��U}�Z�wr;
���-Yj��z�e ���$<$��گ@k���������A$Yt?ulA��P%�x��Z��۳�|=�8X�z�ٔVQ;M�� �I]1�x�f`�2㙔����"���Q��zn׫��Ո/B�/�2�>q=GW�|I�a�,k~�J�>��ή��tT`����[���DQ_�İ�8�����F��E ����\�	�p��:w#�mx{H>�kL��45Fq�+ �!uv�1����k�4�P�jspJ%�H��H��!Բ��!����z��a���1�v�x�o��/pI߇��T��ʪ:TG���F�&%��L���/����"��'�l�q�!�{����ʀ���ט_�įy�"ኹ>b� ��� ��u�Y#!n6u� ���N���A�4�U�<�������}���׉n�qAG|��wԵ�nK���7�~>]�<''�&�9w��s�#�# $�@�<z�A�^?�΍@`��TH\��y_���)mJ�}��G�%I�'���}EJr*c�߹G���ν��������O?��޾���Q��hQG�=}���ŦT�+�$F�7�luΩ.���	�h��Бډp*������Z�;��x]LX�xLl[hzv/�R/�&�ݙc�.n��"�H��&����"��p�;���)�CbG��z�{y�e�6l�M��T�ˮ���<̠�
��l�HV!�RP�a���Gp�H��p���Aj�q		Mv�[A�f�3�$#)�ԭ��b�L�a1{w�CG}��V���dס��F�D4�����7�.\lCNt
G8�]bP���DWRD/o��qꡥO���Z��6�0TC�]Id��t0!i�lSJ���:fn71������v��5
4��2Iª5L�c;$�VHz2:�˖�ȆȔ���S��n-]"ֈ��D8ƍ~���񑕵� 
�X7�)XR��"b�o����eNW�1��Տ:��ګ� d�S�/��n���r��C�Z4,�t��0� @��&q�:��؆pP#"�YϷ:t=�;�[�Qk�����Ѷ�l2�#<gH�W�p��S�D�B��d�w�(�8�K9z��w�
\�#��+�S�:k�tk?+Ejt$n��y}���ɩ8�G\ʖ�k���5��+�Ift��o����)%	���,��X�3�K!x�şD������vOp#�UA�@p���W\ũӐ�#���e�v����^6��g@�����ؿ�ҙ'v���9[W�����D7�7A�ᔘN�:�Ҧ��tf�L[�6�Fk�=���k���LHrXDK�ܦ�q?�_N �3W��<�K����E�d�@�D�'�{��k8��͓2m��yz���y@j��3I`�&r�/]p;��`���q��yQ 7߱� gsV�^eR�J�����͌��Y�7?�JG7<,�@�:/�3ec�X�!��lF��Lĉ@%@��R3��P!��i��<�{����A8�%��_Y|$k9��˶N�x#5}ٵա��Xh����U�1g)�e{��\{bB�j�$%�0���?�u�o��;��V��ݳ� �| HT��fHUc�lC��,��iQS,�R�#E-�+X��]�+��>[Y5]</;1jJQ�[6/�6j:)��̌�JFv�ysK�R���U��y�����~��zIC������s=m<9���k#r��%n���v���aV���ch��I�p�2��"bU#'�����"��Mm1�YKN��l��m�67��IK�2��{K�GڤS����;B}��F#-"��&�g긍"��h8���w�%��C>jf�GzF�k?5�,��Z�YG3�����M�R�I����8l�p���y�dPb�z�ZP��1��0�Tp�1ԍ���*�`T笀��i�0�U���YAC-;+�-v�ޥT/�*�.Ģ���}��_3�z���|Rmlj��YvVF���g?C�B���s��x�# :��Gp��Dr|b��J��j�Vַ� ���]����o�9�r "q�
J�����3��Pk֘k�~��?1 ��I�zwՒ���ؕ�'a���Nއy�F>S˒���&�w:�=�8HڡxO�&-�D!�?˔�^i۴~�&��eP�3hpF9�Y�.O���������J����q�����`(ӍT�9����׏`]t�Z���Y��̥�:�!3߽�U��.�f/e�2I��!���M�=��9FA�r�*M��R��u��h[22��&����
�W��~�#WGPӏ��&���*ˢ]��%z�̿���3�\�̆�h̟!�8A�\m}=��Ahw�4��xK�.�w��X�C@�?���7i��Ç�4��rt�B?��r��/Xk�� �N���΅������i8����=LS��;̛��})!JFd�ğiQ�)ÿ�'�cYULvP�"#��#�����;ٙ9P�7;	��^�*ئ�	��%p��*w*�2�:)��N2����NH����ɤ���ޓ��ga���:�-Z��m;[�w�GW���1��׶���ѱQ�QI�6�خj
��$)~9so�e�"\7�� ��a�+�Np9�i����?5�d��֚ƥ/��˿{ۆ��%+5�y�t��Uֹ�e9ԸSA�i��6�)   IDAT]�&�t��v���n��)."��=�](�b���dHb�ҶF�z��!�����j+�����n�AyR���NFeL�(�:�L&C��B�|(� �f0}�¨w'�ToA-�J���������{��))O}J-nj���]mV�Y�|BS� �/}8��%�lZ���nv��h���&���N�uid�3�)�Nq� ����ӏD�,Qd8CHpJ��jC����q�p�������+�u#��K/�I��xe3�`��b-)�}�C�'k`��1�4�:��ڳ���/�І��|�NY�j�2�������E�b�8�������!H@"v��M������A+���Z�i�;y�;u��r����hc�K˺�z���f�m0���_�v����ϓ��Z����ߵ�Idr��?�������}�cCNT'���	��ڭ���JD����n}��
�}dh�ٵw����3
���˽��E�8/˭aRY��eV
�x����;�$J���=5)��U(�$�b�D����M�)�=��LegOKl�8�ӯ{t&�j�b����2�=γ��}��#mz�2Ee䑰��:�@���En洩^�U� ��ٲe�;A=^�� �]���T�ƫ2�bFy�v��{7��\��Ja�{�z^R�&WJ��:�������za��O�p�������x�-+�=k.��BC\F)ˈq�@�)w� *�-#�iN!�4nu655P��!>�� ����@}�g���3�����;�����{�dHc�U�Ѽ���R�#��~��Ȑ}P��]�	�����[)��yP�&�_�6��Zw�����܄aU�J����Ҏ��C���Г���J��0}����/�]g��C�+�6^���uǎ�}�HQ"�(KЌki3뀉��zSP��G�fR���m��;{�[ۆg��zX���wϼz�NF�����@���Sh�ʧ>�C��9�d_]=���zKG�,�^l68lM��A��@�A�!�e1�*��fp`�G%����\}}��9/�z����@�E�������G�kD��H�[u��]�1� ˹J-<�H!iH[/��H��m��d��0�킼D�t�/?؜t	�Z�rv��ц<�q�&l��$�$�g�L^r���Š�~�:���;�6��L���Мd��ƣ2���KP1DK�Ut�[��,��jqJq�axq\�2�2�"\����ՠveQ"=��Ts�Y�g9f���0f�N3�b����q�@ڒ��&s�tu��Q����O���N�m�h�j�ᓔ'���aP�cDB�@Ǒ���	݈jԬ��Y�$��^z��V+��N�32�Δ�T����3���>����iH�k���ڽ���L��ʠMOF�O��KI��6�\�`�E,��h�p����B����+ʙ{q�B=�� �8$N��2���ǭɀ�]�H���^�p�[�~�����V04L�O?���%��1�ƺd�k
ua���u�R�B����C�ɯ�</B����8&��ePf>D��ݽ��3��u�Q��18�H��qV�ݱ��}��֯[k�i��Ņz����J�C!x9;R�2_���>����P��9yV��ޣ흪M����,?����T^�$H��3�r>[�o���x9}렰��X�ܒ��`��������(j�.���o�������>�PI�|�Ϗ�}y������o6�����k�מTn|ݍY�(�K�V���#�Y�v��ϝőO"�L3Èm,������q��䭂�k�������,O�?���6�^��Q������5�}�I"2�g�̉�ad���Rz��p'��w��]�_��WkZW{�c��蝫��vE�gϝG��*b(x��O~�_�6s�NBRo�
����q�ja4�4���������}�յ�����Ё���5׾������T
$6N��ȢF��Jh��4��ɞQQ�#���vlk�MŸ[i+�1=������ð�H�u�U�'���%�n��'���5DK��P`���	E"��Ġ�D+Rt*�m;5�ک�����xa^,Ѫ�T_�F6cN{O����4z9�\�`X����̑$Sn%�6f7��b8U�a����/!�9c?^�Z��l�1�����ʹ[P����Y�J]���M�^ ��d�]jJ�bL���r�R���ǚF:r�  ��[��g�C�]Su�}���r�._6c��AxrJ��?1��!G��=���n�us�F]�z���f����ɑԧ����+�&k�@�k�D���O��@���p�mV0|2S�&PV3\����3�Q�%�a����{i�5��7�թ	$������ *?R��5]����a�
}�58^������r�jU�A0��P�L��A�.���.=�-f��D�c���\g�����D���g�w���k��B�#��h��� y��>�я�J)�pg�bd�Y�����\�(�8�[�H� �%�gÖW�]������zȔ���	"le�I����~n-f��?	%�����Rg>{{�.�#��#8��z�5X�I���}Ͻ�G$��EP+?☻��L<��'��Vf�w���eR�j89�,��s%���T[�셆���t�
��A�����^�Q��Ͽ�:b�0�Q�B�P�����ut�=��E��P�[lg_5��f�0H�ҥ����r��c=�>���,�R`�\�� �����F�ۍLx�u7y0�he���]ǅTP�ɤ%-��9�zT�.:���8`�-�8�>��P�L	�j��(5���|С��r@2WL�ѱ�ǰk�(�V:��&�-�>�s��=2��D?Rcd���yڴ鹩��onS�%}˻�WX�_�%͵WC��~�_���7�O��y��$赹��bMM�����g�7\tɣ=n�������~��=rh��ǟ�Bug�%��ο~�}퟾�rGF'�r[[�����]U����6�V�j��]�0��6яJ��(�I���u��d|�`:�0�n��*�2��l2]aF��qiU]��T���e���2�I&V�:ab���lҩ�������W�f�Ah��l�0/�ƊR��X҇�)mp(ؼ�A"e�}��oqSˊL<cT�u���Y1��N��x�8�Q����J��70vR.��P�~{{�;y/��yἩ��i��#x9�q��u�h�I�P|���K'W���ׯ,�C�"��M,a$������B����L9����������{ߣ&]o�A�jk�(C���\�-Kw�q��1��*d��m�J�~���V��V
H۶6]b�����L�(�c�ջ�#-.|�{I�F��%����V��mcL�5P3׌��W#��Y�4ξ[?�W��YC��C=d�=��e��׬�13Z�ɤ�L�@F4��`J�����}��[a��{z�Ҧ�/�IA~10�\�p��<$n"��4A��sO�����	?$�tޅb����v��.+|�7~�?�FBS����HS
F�Jߘ4��n�+ؐ��`�p�#d{�N�A	�(�n�ƿ����|��aN�:��q����!2���U�W{� %��'��������)U+'x�DmT��{ ����AJ4��6S^�%��rJ�-��J�[�O����萐��ŋ�k	x�̱yZ��Dz
�̹k�)d���/��;���Ŀ�c ��8)���JD�?��l<�¼�0�P1��wQ��"� (a����f���`���Սz0c����x�G�=͂e�0>o�;J�P�ӚVW_��/*�ľW���0��-N�����f����@�g �gP/�K莻ؑ����"M�-4��rK�2���G�v�fsm�R�.:*ޭ��������ؾuvcM��G��o������������~��¢Ү�����S��%��?��?�}��t�?���s'n��-���]�x���������!�L�*B��df<Y]�J ���<u��m{��͆��|E:�P9_�6)�vJ�n������fys�QNE�>��q��c���V�&�#S��t&x�d99W}�3�p R '��*5�z��a�fP��Z���[q���EI��\����l���x���&�N��T{T�7�p5�ݴ�T�]�0���!� ���F�t��-^4ɥ�'���8��^�I��t�c����M�s/��<ƻ��+���*��&c)��eE_�e%���������NYC��T�N!�q�������F�nnA6�_�)#䚳S�f�G�B�[A�Ԣ����%%��2Aȉ��@����Fw��+���̀�f���p`��r��Eҳ5�/�x샏���a�b��7m�*�X�b(��V��k���e:Y�JڤV�$X��ն>k�$8��ȉ�7��RG���2z
�,�?ד�:� �$�~:�M�j����k��;�� kW���1�u&7�zM�n/mr=�#d`0��ֵ�ʲ�z��ښ�n$��(�jv��<�]GK�b�� ����)`R;ؠ۱�uw�)`Q���z�'��T��\˩F�6� �����[��|���vZ�16�R���/�a����GݑF���ܜ9���[:%�K��>��4V����wUx����В+��^�uw��KЦ}$ƶ�#Ո@4p'�aI�bIw�������x�'X��|�M���y�{�H��"��(UC���nX�8?�n9Asx^��כ}YE#�%�$�>��ov���./�o�#�( �%��# T�	�A�]rs	��p������	��N��j���� �1r��(���
���M DIe�)��~�MJd��e{�T�*�Ze������y����;�ޅ�߉U�w��/����x���Om���)9�kɂd8U7�f�1c��߾Uo�v���}5�feD��l*�/�yo�����	|��WZ\QoZ]'ΉCU@�c��L	Jř��@�ead�����*JpuUνN��O���ue��dpm� �iqX��z�ͽ�|�{��i�q�~��u+��&��xXZ�*�?��8���K��}���8��.��jޒ�T�fк�1 [��>��D���k72M��m��q��v�s�l��o��ZSlʠ�6����`���A�V N2����R7�N�@z�����cݾc�nˎ*�M��6D3��/r�f �{M6�n`�#�Q>��2en���qP�� p!�͌�Fa�e��c�>d�(����͒�SiBD1E�!�ŢEZV���y�-����4��}�c�6�AX�j+Rv<o�,kҔ�1:�"4����}�@ƷԪ �������ɶiב��F�������ní��}�$o(��>�h�)�tR�W@���" �\�1U�7���h9iD���{\[{�[j�$���⹆��c<�	��%���3�T���K
#K��"#㹖X��m���o������B�Z�����mhh���ڨ�hr��+���iC�̢KA=�r���>�y�9Iۙz�Ǯ�s�������ot2b>�zx������n\���g_��yn'򭪮�`FN5
'"2��>�a2�0/e��8��h�#c��:e�r��y��� "1�	f��J|U�{!55�4��U|�H�sw 8����Eʤ�-��Qj�gΜt��i����u+�3=a#�eSW��}А
x�1������8B+Nj����l��ip�֮c|.�i�A�K��=��M��ʃ�Sqe�68����Z9=7��	iz��/>(�j�G%�٥�OAG��&�s���$h�����+���΢�0�`�MUN�gT\��M��u�u;��Vy¦�����GIb.[)'33De��[��ѳ`�ˡg�R{B�MI�}��<�N��w�eމU�9��O����{��d>��G�s���0��XۋV���8�w_ί�x�^zA~�+��w���k��		�Ԅ�Qw����ʹ(�8�azU>R���R��~W�dpg+�1�&f"͊I$r�����΂A��m�H[K�[���e��JٰKό7�r'*aq��Z� �1�(����G���9N*aYld2�3��Q�N�:�jQ�GF�`�H�a ьY�GP$rZ'���K�88��&�Om�>����g����I��+&7e$a�,״4z�G�����n�-_=�ŧǺ�j���q�4���V�pT�d(�T�y�B��}ne�^`e��h����]����
�iY�9tB+�w��j�z�C�V������g�{�k�R8Yд΅�ȉr�UKmd�Ȏ�{�	�V��}Cj��̘�|Yy���?w�{���(�@+h �%k��-�D�iZ�Ð�੃K�,BلJ5\����fz�4��08c-QJr�A�Z��g�q/���?��*�W��2D��K崹5�^&��.�C�d�?�����Zv4.Ǯ��a����80�$Y�ù�8Ig�O��/Z0�����4G"������W�q�eCp"�¡kgZ�m3�3��KF����L��Y�@�C����J(���t㒁���y�W,#3�XZ_8ҽN��q6W'-jVn��8�e7���|��Fj�ju�d�ަf�l ��{���Ϟ���R�Γb��e�EI'\�HdH��h�L2�+�������2���	���5���l*��9&�$�X��Q��	 �A����_!0��G��WR/筽�?�i� M�#��^~9���ukܚu�(� tuQ2��"�|�/��+�@F������b�K�V�_���o:AL�����7ڼ�|��2ͯ�B���ȑ+Ȍ��[JzBu�ίgO.X����Us$kk:�v�C�������� ����ŮA�{���͡�4���:{�gׇR	�42��d� -�6h�ֈ}}��rC�:�wj%oz����?��?~��5ғ�yĹPQP46�tr�%�16��{ZSu�OO�?��w�WߡG6I�WщI>�����x)����8-�aFr��m���JWy��A�d�d�(�i\����y�v�D6m�E��>b�Г0�%%�n�\՘�܂��nʂ4���:��C))��$57���
�5#��!�e�K�\򙾧����� �00�8Tb�"�ʠ����NV� v3������(WY�r[됛��
���1�P������ՠ���^D�$�Sh����t�K�ݱ#	8z]gG�E�lR���Ip�/��]��v�+��N ���e��U��N�CH�>���I�Vk�"륉`#�FRH��ĂuwMsGQ�J6&�,�婇�����&[.,��/Gc#NɆ11����Z1��������XD���Q�� �X�k;a�:|�C��a)`R]W�B�D٘���7L�����P�w	M.[�rY:�83vc�2�\W��0���ܮ�s=e����+>�06�8\#�LMCZ\mT��2_i?�RY�FK���$A"e�?3?$wO�#)_T�BV"��8�^����1���m��;?�D�"Lw���g�ZUDL��=�:�DQ�=�<eh�_���]��HZ}����G�)�v�+�#��\�s`p��Ww��/�7^{�=��G���8h�%=7����*T� ��:�7���N�}�K�$��@LJ)S&r�5�Wwǘ�.jI碣�!���p��"G��t^��l� gb˖-��~�6�l���r�v_�s��^u�/tk�l&Q8|�N]F�O����18i!���Z����c��J@3Pɓ��^�9"�Z�ω�A�K߀���h}a�yA��jS���w�VH�mt�� �!�_��6�a_�^�w��n�ޭ�W��D�X�=�DT +�~P�J�ԇ�x;k;տ�/^mi�a.8X�d��������2z�X�mO| L�:��I�����܅Q��i���ʡ�G)�b4�D9��f[����]����ܿ�:�������ۇ	�S���;�#�����|��"�(Z%{���ރ��� 뱚q�Q	������[~������4/��Kg�y�Ys��}���tPňVmW�z�A��N���<��`�n�Tw���M�遂J˒��ىn�I0eKL�g;��+�]F.w��2'f	�5"J��:u�TǏ���,9ä@�kbx$5�f4s��O=��m�l���L�ٮ0�)��t�������e�[dd�yMŒa	3]y9�f=5�\;����uBT���"��m���2�^n�s5?����zYG`�Ą'�z���8�he����R�2�:x��6:�ad�L��թeS���$�>%��f�ˉ��N�2`1��r���)Wq���^j1Rv)Q��ӧ@�Z�s�A�����o!���6YT��*�3�eU��u�,�b�!�;��4��QP���h�k�ɏ I7s�����^H��+Նg�jV�J@�"0vI�	OERZ�@�%���z$���7`2�
��n�n�a$+���Ai'�}�O{�����dR
��%���(�?�f��i&��N�$�5$��������X�.��yHU=��*�v��s,CNz!��b������H��� ����������?�s� p	�<bP� �P�����'����O�A9EՊ(*g���!�?�N�9Ѭ�m}��?��f2?=��=���!�� )�q���2��b�D9�b�r�Q����"J�@��qƛ6o&����CPТ���' 8w��������~.�:N��o��^�RO��O�#x�s4@�jAq�[G�E��z���������c������6�:��ZZ-\,��fd8�X��m(?�Us�U�P���m�������{җ��l/�G�,�7�g/��,=��z�o�ҵw�XL�s}���]S��ϼ�wsM߿N��@�2�Vc9t-� ZE��ڭ���	G�dÁ�Z��Sg%2r���L�޼��ؿ�u��:�B�z��-��׿���v�#{��K�C������}�F�]e��$?����1Ť5kow��6�P4��~�o��"+������o�j���ڭ`j�>R��2b������Y��Z\H,�"mb�M�~�^�d*�~jS3�����"��G]\�rW4�����	��sG`���O2ѭ^��.;�o��4���$�-���.0S��>�����Ғ6o�b�x�l2�JHf3����lWb�^�il�s5�DF%1��M.�ݽr�"�i�
G�iE�"~)(	w�N�R/����(ϓ@��@��M�h!�b�8�5�q�~�˦��ٕ��+R��f�3`����'I��3�_�ץR6F�]^6��s�xp0���0�� ���":iD�j��#����1����j�W]7�'��8�a�)�]�Q�nE3�|�Y�k�{�Y2O��0M����h=�R�8����� O2������5�c��U&�b�4��2Q�?L�<M��������T*�\�h(A�7��S�� �A�egϝ��p���6#g-���qn��%n
qb�ېX��P�\ځZ(�Ș����d{�L
�u�A��U'-�Z���C�ي��%�;�����7�@�[��� '(L���d�!��w��n�k��t	t1�g`(�t����c��\�ߕF�4��+�lM3��g�񔜍w!Vx����OI��er`�	�.	�DXx����p�ǭ�{#t��d�p���k������/��쥯{Ls�K�?=�L:HH�"T�u����T����D�b�� �0h����1ic�!]q;���H? 0��� ͘3�͜����vA�0�����t��p��������t9��V���H ͐>F��*$[��D�3y�e���A�nYu�����^[�g��Gr��mot�b�ap�uѐ���*o��p����僠ؓZ<-���۠u? ��ϼ� t�ל=Ͻ�u���+��B�(�q{�Dhj��VŻ��a�W;��j�җ���9�_�I7�S���}D���{����`_�\���{������2nWt(�u������;���3�d�+�2Yc����it8�j�q��b�FM �b$B"��E��&������Fwxg5#1;��2���bq:#(��?����bNI�����#��2ط�="f����;��G�;V���+\L�b�WF\��u4-0�Bx��R��[[��@�2�ݝ�0]S0��x8�^�.2ܥ�Ѡ11D�����%��|�L�֩����fR���H��҂Z����U�N�������F���N�:[���٬��K�N%X�u����f���sYh}�8�A@I��!f�/b�g`��d���Lhz�c��n�c-!�e�Y��Pp��M_ �G ʔ7n�z��X�T`���z�5�A0�MS������ګ�D!�u�0���)vW��c|�n��������[�)��e���tȯп�����z�E�y�J�<�,�;7����HHFz�
@d4c��7���_�k�l��Ɏ#��U�V �:������괴b U��u�} d������
�9���m����u��o7����^�xgJ#�^��h��~���.���##�#h�\)���b,�v&���r|"�y��O�4A6�K�H��X���̑G���)���3[`���w �$�p�/g�SSYH�?�y�H Uq�4�g.cN����)8��`4��s�C AI@�����dY�u�\���c�s�A�*ݨ��PŽ����C���sA��؇��hڹV�Z�N�b�V5��A�{a�BBb�����;�d�)�ः�9��C����Ӳm�YB3<!P�mZ���4ƴ�ѥ����У��M�J�8�X�Z��|��%]<w�|�Yo3"��5�	ԃ����h�s]� uA����GV�6ݛ!��3t��������UΛH&�F��I�Nb������e�yƲ7����h�`÷��]�oU
���<Dφ�w	9�Z�w��md�p��r�K�o|�$>m:�<��L�T"��Â3��\���\���ƈ�'O�YeU����
��2�Y���MMl�P,��TDJv���t(cgzP�ajF�XjF�7v�=0�ߝ�9��0���q2H�6xn�dj��[0�����{�>Fe΂Hم
�k�����g7_u{�5����r�W��Yc�Ca�Ҷ69�1
I�'/�����}�7�|�8I���Z��m<�Y��(�����I�]oi ##+�pO�/<��w+
W��� ��]��ZC�����j���L;��rBɶ/���� �*�6�/����o���ҥ�})�����������ц�t'ڒԎ6����@[C4��8T��oZ_�å-d�ڷȇ�753]��׀劔x2L�� L�Z���4�aNW Jr��F�N=�da8V�bm[>p/�\�x�����4�%��E���$����AWq���w ���7���������z��P�sh0N"2YCc���)��K$��X�7�l��v%�f�����7��n���XNU#��d����1���;�����t�qX�jS``�[�'�觯!L�{�ͫ���/|�{�J�eJ&��t�.�b!s��8�88UA��p>�?��M���h�H���؛D��7�8���a=�ʈ�0�aȲJR4��w�Q�9�x�.ڰ`�'����k�!�C�;r����>�ֺ[A	�,���%í���*(�y����d�R�S=Xu�$2�|ڝ��c��7]��	�)��%� H��*QY�K��5
��qس��I��щ?L�(V�m����pC|�w�M��|k�CE��g���J76zW���A�^����h�\�z����c߆�Õ�����f����up1��� [�鍒I}�OYϺ��h�L�z�5��T]]��>���l�ȣ����L�i���k1��+ֱ�8r�Z(k)��Ss�ϖ=���]��A�-Ru{���A��+';���N��{�TTU��q:Kφ|)P3�ͣiV1��*n�%{(s�um�F��Ե� (�-06��{�=�]�5���6>o?HS�ko��+� ��hsX�L^5��I�44��ٞ��W�Xa?��x������X��u���?ȬBn��P(""2nܶ`�IԤ���U�)���Hmik^t���S?������ц~��h�W���_����mA|�~�a|R=�d�3�������).�Q�ƀ��v�D��Z��t���!��l���~F���B�G����[\w�n��r��TL�gj�!�H6`�B�uM����� R�	�$�Y���tV�z���ɦKJ3q�dtʺ0���>W]��25���uȫb��\6N&��9��������d�C#q0�ϸ�)�pԳ��Z(H��yF/;9��%����������h�
t�{��dU �b�53[Y������{��U&��J���Lb�R��_�m���|�$Z`r��[�+T><��^~�Uw��I����:NV�Jq���:%��a��H;D��;A CUZ"���2Χ�}���s��2 2rM;������Τ�4��hR2�e�>����Y���(��^���\���e��A��/�yk�j���i�����,��t�TO ��k̷�Lm=���K>�Fh��+e:�9 `bL�f,�����exh�H�_򹚓�5�Z�N*�:ApC7bd��T�'ʸ�#S!:ηLX"3�0&��� � �N�?~�t䀵WK�R9If��i���7���rK�̳��_1@t�!�	�����͖�N�R톬K$��z�]����6�����{�<��X��M������ی{�#��Jd��L���>*�j$�kNO�����p�l�9�	ڞb)�-�?�Ђ��{acG+1�=��4�/�eP79ܫ����o���>u�͢��2�����rPF�n�.��
b��e��!��!:*5)����0�Ϝ9��2���RaJ�nT�����[�`@�)�DE�������ϰvV��uڗ��7걟���=�F)Z��q�߯��
<�c&��e3����2n��X�1FG��6�g?	 �
��fZk�!���T�陴I���Rυ��3!
4	�,�|W	_��;��u��f迠Com���g��t�w���b�����db4Gbԇ��њ0�X�^����T��e]8{�mټubƬ��<��+����K��=><0ú[�+Ô�����(y��7��Z�vo?�f��^����!��,�˵1�_�~�͛��������V6N�r��)
oϾ��vl�r_��B��#ȝ�B\K�ŅmlDy�
�si�R��~^_�L�N�1Э��,�?ť%qhB�ho#"nnw5W%2lu�9�g#�z�U@�;�C�at��J��bQ�J,u�g��	%���iO֯���LOP��S�6~s�<�f"ㆶ, q���-��?��,&^
��߫� ~���Fvb��Fɶ�/���m�]��P� �R�M�7��m�v��RmW*��r�'�+�������`X�!;��F��x� �V��N�gdā5q�cd4����@�+� ��	왽bTG�1�
��A��YXThN�Gs��k�oH�f�=B٢7}�
�ަ��z�"���#��c6���4𷽾��!��]ʘ�,��䘔E�U������>@+�T3^�SJj
�<\.�0�~̀B���+��|��^�}���r'VC� �'�BM���8��H��kS�QvN;��l<�щ.���@���������k��8D�>`�V�~�|܁#\yR����,��z��{��}�^��$}�C;z� #L	���Y���>ao ] i�k���x'�U��Lx��B}p�M��C�X�^Yz?�]z���+$��6s�w'S����ȉ�W��
�����p_G�l�!1�������^@���E'�1���G%�$
u?��f��7[���J8�{�����81|�l� '�^N��T�����Z�hN0 s�X�6�]����5�Y����>C7Gk%���^��@�4"���-�07� �boqa�M���}?�Ն����M� ��˽p��&��c���Z�^�(�Q���t+���l�����H��J�$S�đB���ek�F���v�{�E�2x�F���-K�|�tA��������e����w���omy�_�0��`��1��os�UX��ܴv2���٩щ���8�,���#U09sm����A+.*}����.e��w�����9�K/����8,�9Q����]���7{Z�ۿ�������k'�i�S���q��g�ǟ<���;�{6΀��(X�7�h`�q���������?#dO�:�^r?�J�D;cjۢ&����.Ћ�t�$Z�hA�ޏ���uXq�Jw}
5�!7u�t$U/���뚹���3�!��1�"���8����F�述  @�h�r}�#��aLJc�ʡ}(l1=m��9.!�!*���.��9��A�2��1������ ��4h(�Hgb�r���gϜ����s/���ftb(y���a R4�PO2�����^�1��;��Z���-)�!���Xt��s\Ru�+��{ ^i�-�, �`paQ�z��;�`t�k�����ɺ2R��Fb�2�Vs�e�l�:T'${ii�q��ϰ�:	����ÐH�>��"C#����|��*7�q�"y	�hx���4O�����v�s�,S9n�̙콅�*�M淌I��Z��Q����(`v::!���9!bCc�3J#c[i�C �}<z L�b�	vpv�9�fK P��F�7DHZ��8{����x`t��"]�
*k�j��BW��� F���k��NI��8�h��څkH�wG^S�}i���C0�-���T
���3@���$A�F�?�36��"J�'�A}h��<�_Pb��<s$��C����X�Ps>�d���Ԝ�!�p���9s[2$��觱y�������Q��=��m�l�d�5���w�@�N/�Ơ����Ar\M�۵7�r�j-ZD���~�a�0�j��"����̦���;���hoeN-x� �� ��X;>c�����aH� ׯyړ��C�}.]m��j�����RK�v6�]����+�7�BA%%�e(A �d	 z������6Ic���\w��6s�Į��-շ������8�5d(Qh}k[/{M]%ٖ�����J{�֨�S����%���C��jj�M8���4����ږW�`B،����{�=|p^eŉiI�UFp㗮z�ɻx��=��@?]��y�Ϟ~f`��,�x4h������Y��-o�ԩ�qBǑ�m����AMJ�cCd��WЦ6��w:ܷ��Wɮ�0,��ݱz�[0����Ĺ׶_v���!��2K�3jmC=�!��G��i�:ه�����r���׶6�S�Ƒ�a�e'��x�~�D�_��$y
 �)��&p9X���V���d����"�*"L�L��Ă�.]8�6�q��5�u���lz�qcc��\u��:��Y� �־w�*@kBM]� A��qj������3��68&G,(�^s݈�Ξ�`��k��,X�^�K�^��2y:l���L�Z�"��<��f�]f(V�^A�E5~e}
�XSx�XÙ�
A+�d��p�T�x�bDz�&1�ɨ�,�b���];A8�m��Ū�k���5�V���0A��X���OBü�e��3�4-k8sap�\������eܧt�Sf�$1)�E�
�t��A[�����5�+ R�ںN�Uw�^}��*Q�k��KC��d�B�""�0���s�a�Q�ǋ�/�Al�h���3�M2��欫���aT�-�$H��ᬓX�d6>�hATG�L@��d!�AZ�I��x��h�)�&�Xͬc#-�R>kmg,їHb1��'"$&�j�,�d���5�	��܏^#�u���ڍC'@��>���$zŪ�e.�ܒ�I�P�A~	0l�M�����<58���R�R{����TRP�;��\�����a��B4鳁u5"U-l㼟�@u���fkY��R�5Y��%��0]#�t� f�X���u�u朻�bڬ�voԽ H}ւE�l�LZ�(��``��H�(�1Ó ��%��>	j�_oE�jq�c��#�L>W����U�����~����H%/��6##[�	/�*A� \�9�xU2�%)�J�S��Q�^���w��=�{��C��oL� k^OԿ���p��䚏9��RQ���ulxdA���B
���h:a+��!��� �k��-P��"�t��տ�S߅�oZ��'�9rx��dkͱ��%n �|x<�>������B��'���;RPd���?<Vt�j_>}f��}�ȡ��SD1����<�����~��y��gV~�3{c�������/Z0o�tց�;���m��$ڹ�ٴ�D+ܹ��0�'��S	 ���#]U�ko��E�-#
q�TX�~��-����ų)'0��lw�\�K�+����,k��D�0�'13ee)��Z��"�F���7����oon'S���iB8z[A���I�ې��C�uBJu�㪖2!xLMWp�����!wx�˥gx�<4�SP��<�VZ�d�u=Vc�lUA���ַ���U�4A�;u�2�HA
#U׮^�V������0e�z	�E�efA ����0<>�Y�����abؽw���d6w@D!�Ui��(���[��xpx ��NHE�I������{2�!#�xA}9���-�l+77�}�C������sq�G����:�Y-15���O@ C0E���4�|��r˲@���O�X�ސ�H�GA��YȺV#:4��[�q�u��^J��� ��#(!1d3MMd ���Ē�Qx�r� Y��3�d���%g����E�q|8
�C�g"	�p��ea,�����L��Ƃ
�$��!�� +?��ޱc�;t�Iw����*v~�{/�</]<�D�o�

���qD�Z�kٻ"���t����CN�C7
���8f���b�j:!|M�ƶ.�uO�����h����QHEw��nǮ]��N	�aLLNQ�d��Q��)aT���͎Ǳ����kLl�0 !:���9=��6��X��xM��]���]��S�������h))'*��պr��U!����������j�ƶ�溞a��%�
��z��;H�������O��T���
���[0�BX�j�"�JdHb<�K&�����W��*���+ٽ���K^����� P����׾� P�Z���'Mx�m�N��.!!ؔ��V�� ��su5u�ӈg`P*D�.=��BfrM�|ouW�p�Q�%���������n�X�KgS�����g�=D�o��dE�6������gw�����h��C�G0~tʴ���;�3�]:{���_����Y�!�=������ޞ����w��j�b�JmL��	�5M�d����bƏ�UU�F�_�ꖭ���%��/s���iBm@R��Y���D��|,�Rz�u��a����{������c�Ϙ1	'�T)a�R6�g���7������V�!'Cv�.�	g�:\8f͂��62��uA<�aq@��i嗔H;g���6���(zʯ@"#@�AY �5uź���po�nt�='�-K�6����J��Ū�3�NSeT�é�ӽ�(e]pEʽL���yͫ�	^fR��B��bwgn�i��wHs�%E���"@+J��J�c��#��qhqj� �d��M<���x�=?>.�`���#AY��X��W��4,ʰV�9�Fǌ�1�4<�Q�u���{��J��'��h�SgL����J�`���]����6?]����=�1&��'�>z�^21}tDD��{�;I���Mt���Mp(�(˺�@&ƹr�!H�feS�K�Ӊ�k�t2Le�":��Ц��Q�qXT'�OЁS��y�@Ȅ�NR�F��6/�3կc���u6F5PY%�Je�v��E��m߁}<�y��L|�B4�&h$�w楗A�@i�$ ���4ap��%��	�6�或�ÃF��̻X'����|1�3ӳ�1�`5]�n��9cn|_�gS{��q��m���KL��Ս U��%a����{���~�{���v+��7��BK��V�Y�Μ:��bMR�]&ݬN�Ԉ�	d*�#�� �Zm[�m�����@S�2]������^���R�m�X�����{�� x�q X3i5)�8�T�T"���bдx���6X����0&9s�];C*1����8� D� @Z�P6�eN��T�/	�S'���(�ꢂ�L��>�f�����!�M����+�ͦ�����nM���,�@8�)n�R��о��Ć�\����wz`�����՗ί.,�����۲U�T�0m�L�������M��3i��ל��[o��؁�e�p#�b�[s����ϥe�t�Ջ�R��֮[gNB�'�{��HH�8���v��ry|NƤ���m8��{�����YT���9�C�Mr'�c>���6�Hˈ<ICq��ua���}S_�Z��~zP�JH��PeP+R�><8���J�ȅ^|<u��.��#d�Wk�\c݀)�i��KDP�-bpS��ĪǴ�r(�!"����`�&�M�Y�\8�AMp�H̎!�0��_ϞC<c6m
�o����m�ڑ|ő&��|�Yhھ�9W�X�6l�tYj�V_�݌ukV��x��n��ɞE�6�w9�ؽ������Z:cFBb��D���L�v�g��x����]Cig�Wo>��{�����ԱatI.��8Ȇ�m��؅�G��vs��G��P��=II�a:(�^A�2��������R���յ�{�ɔ��Q0gí�O�˩)s�j	��lh����]�$�i�:ut��j�O�CϹz��)v=t(H�M@X���q����W~��e��p&@l��8l�h�[��04�G���������
�2\��r ��abiO���5dh�����'؃���$��0T�
`nO6�X�4���זa�K�EN��_�J	80#�q>�i-��r�u��R?.�J�}�,C��}Y~�:k���9��rt�|VҺr<eS������ܯa��T�Y�c ��G-`YY9�dWTXh�5ͅ�3��l}�e�B��LV�C���!(7�X������ț�a��X&=���d�˗��v�*H��m}�W�}
Gz�R�݌��\m�@�rغ7Bv|�)��#Ep�g��@���X��3�_c�_s�>$�	��>G�U���!u�S��:e2\����?m��ʹv>����j�U*Sײ�`�>�����ňxq"FBdMI�d���ȉ�n��.���JQ��/�N�Y��܃*)`���K�u$I��SB6���7�MrA(�J2��إ �k�v�.�%=���?���_�u�,��~�џ�:��]�t׽���w��7۷��vkc�#b(}F4��HGP
nӳ?�|�jK�ҋ�޼��7ә7o~�H�Z�Ĝ���nm����^Z��SO4$'&�EE���������<w��,���LJ��wd/��&��r���	~։G���S��n[	Ae�۽s�[����	.��޽��a�s!�iZ�nA��q���cr� �J�]�;��+��?=ǵ�t������O��I���X��K5�J}�@�½��T��3�1�Hr�l.f��X�;qޕM�S?�z�yw���ӧfAt���N�����GN`c��[�����U�c��!�Q��5�����v�=�XVs��w�ʺU"cY
��^~eQr���F��?�k�@����n���lɣ�k�j�blf�d)Ā
��85�ph�bJܦ�O�Rw�%����A���0I�>	rW&=�����M�i_}�#��ҭe��<.q�;��m���'�$��S�T���3yޢ���� -w#��Y�UMr��'�'��X֪�����r�U��>���k6 Z"��������ug��rߊQ�[��α����F&����i�w'��7Q���e�Z��	� w���>A�����%���_m)g����TP��P��@^�O��? ���K��r/�{ݣ���������N�������9��-�+CK�={f	��0���H^��7܏q�"{���}8A`<są��c`��E�&���v���5[e��խ��e	MB�;������8�HML��(x�f�R,�tn�}=muK�Q�� ��<s`��a���q�l`���F�*V���&�="1J�2��"�Ρ�����yOs�@���}���{��H��Ha�x9C��bPs� ��q�T��#(�"�o�h����Z��ǁ @�kcm�m�O�	D�T;�t/�O ��	��EO}%Z�ړ�K'�2���5LER�a��"�F/�<Y�^�c9IA��p���1�&���K�Z�e�*��./Ū��~�Y�$�Ѳ#����yoD����:k�:to��d��OTv��%I����2b,�#�~�,}������������>��o߳�at*���\{]KBL\fg͕K�zM�#fŝK�Pq����x��������g~�2Q�:�����H1���7�~�轻���o�3S$_M!3�p����D�@_WI��j�1Ծ�M�&����q�~����T:��7?��[Եa����[�s��L/b�Ӟ�jܴ9i.�8�=��dwho�����?.c,c�1�'h��t����<w��e���̷�bU�Q7%"}���d)�~b��O7���[=f?{A��>=�΁4c?m����U^h�y?Ǌ$��lj��@BܺeE��6=w��3�;��wW��!-�m��y$d��F�@�ոH��"���aDn��0���1�fUe�ý�iY�����wW�^���v�����Iւ�~o5�=K����O���F7H�YUu%�͉h�����8
��X�Px�>�n������P�,��� N��u�g�$�R��UL�����jH�F����iU*+��o�EI	O��q��d�!�����P�-���2I��y��8���~� ��ׂ�听�O5f9�2�y�B�{��}+�7"�Ȑ*�����mSie�3?� +�]�~��6���m�D>C{A#n�rLdJ�F�J^FW
XC��-�υo���w��B!4BS� ��	���fcu�{.�Z5h�ZEi������[uk6uy����)�%4�	c�SǑ����wӪ�g0X>��"�A [\4� .����\�����Ǎ$c��]N�N���ٸ1p}�ixE7��o���N'h]�K�<���4:~.I�-h��:~�1����"��	8�x$\��K�\���z;�S0$��5��=����'a�	��`�4�pDbH�k�V��&Kp� Й [b�^�V�(�Y�[���� 4���9���l�߈�y0�%��~V'7�x�V];+����1%,+���c�����p2�3�D�T�n���eͺo�S���z���/@��7T��3��r����̡�ޓ:��������X	籈�O؎DH�2�ܸ8v���Z'������o��1��wХ���r��aj]|#�o��6�l�߉��֡�ۻ'�o��O?�s��DT�"4'����/��k���6S��`(ɢb�\yg���u�|�"pd+u��_�F|W7���7���ræ���}_w�,���T_NI������`��<jr�E�!�%<d�fd�C��(S�n����G�HfN�W���q���Ŀ��/<�Z[��=�� m:�� �\���T'S�&��U��3t%ս�R9�B����(�ѺB�����PwۊRfI��=��j� c8��i�6�9�!�H;��l7{:��T�m�B;��`��#�ǰy�-�c�)� �h;��o �D�n�t�z���bD�jܙ�dX�nni�[�Th�H�;}>�}��v!�A��k�"���I��j��= ?��}�:�Jظ��!S}c\)�Pl���L��l�"���GѲa"��SG�A��,� ��tZ9fp�� U�}��n�TM�K&V���-&#-ap��𒰕c�CL-�� :Vph��,�Q�k��Y;�xlc�~��ket	Lm�\q?E�� ��.�w1���lX	�,$*�IV�̜9%pk 3�ӊđ9r��rM��Np�<� �^�I��S�����Xp�X�f��א�ù ��S�p��.����J-҇� OJl+�� ��F�UduQL6�\�"7��7�'x�k<�c-rA��-��}8��h*#Hg^��P2m�8�$2��QP�e�F��l�qP���9J�Ԅ�E|	x:�`$'/��Iԓgs�� +^�_Y�^5]9;���j��Ct�����n�وK0L9�4�Z%Ѫѭ^�L���8%����#��rKb4۷�NO���p#��!"�r�-��Ç���w�F�j�Ԧ�XP��q��:}���tw�ek�h.����B��]d�Y�*7죖n�H߇�^�y#}3d��_���Q�e�rXG���3�d�}���CA��j�RBC�/�$V�p�@h�ԩ�`�z�oIӹT@=�Ɏv�����^e���	�X���h��	5�1Z�9�y����ύ�{`�z�YQBO٩�q��gL}qO�������KXjFo/����y;�����@� ��Ze�	
�8tF��z�7�w����㑣��^z�On���G��ۋ�4L�2Y����c���?�ٓ�q�S{�� ��R׭��
�e2���0u���g�%,������B�>��@��ȁ]8��l\�l�2z7���߇���N�8���ʷ֔Aɸb04$A��/\�}��_8o�ʊ���~���~i��i�Hnl^ի�}��.-��p�O@>!a���v{.cVqԧ�?���[���Ϳ%����"<��%�rN�]ʲ��`�_��%!���[�F���'Fq|:�r�(�@���pu]@�S1���RHY	g]���Jg�ۻ���X:�����H����.��'N���5��âl����G�"Ʉ#�Vv/5���*�Uj}�U%����Q1�՚"��N��D�@ =����}�a+���+B���Ѯ{.���^���ZL�����a�f"�����k���=�,M�BD��C��IHø��\�����j̥��^<�dD���t'�a+����,rY>s�ZoƖ�;�n�>���[w�Xa�Ji������.Y���=����'c�������I#iL<��n��b�^"ك�s�&���.�pz�]2���Fodڤ?�z9x$^N3����+�TУڻ&�P�o��`/�O8#2/�LM���ӿ����Y�t�YF���'�)fZ�8��6�7&
eBe�L�#(��E=�s�_	"���T�%Å��u�o\.J�H��ձ�_�#J��zh�J*u��=�$-�}d�*g�Hjn���-+nq��w��u�c�}K���+/<�N;f*cJ
���5jYˠ�G��H[ih�������,CTG��'�uhd�DB||��� �S�jm�rk��OR�]73n�V�1�	�5f6�˗.�J�, �Q9a_�>,������Ht�N���mԜ�'��Hz�v�^��;t�uJ	Q���[�L������pz��a�nCq�p�8j�+2����t��{���D�g/�}��A`�NP� \A�`y�-�m�Z��.Y2JR��=�9�@$�T��nހ���I���']�F>�(v��Db� �AR�	�I��pG��N���Vvj�6uV^fFZp��t��?��w觏Xq�������-���8�OVk���qT݆�e�>0#���in���.��ۣsUfBa'jb���2F��yk�6����v�����=��Vպ7���ێ�i�E����z�س�^�L=2�mdD]+��89����C�z�������1##�������8q���zмge�l���{� z��uCA´���MI�tœDй��0J��|���Vw��2j��h�O@z���:�]���;�U]�C袌lz�MZE6<�HX�Z2vjt=�!��\-��\S<�+F� ����"M1!I�8�ό��?v��!)�V�/����s��LFk��s��q3h�q$����F4��
�QK�쓂Ti"�[)G��r8��f{Е�C4*#=�_��G�|�5�:�ΥD\��� �x�'V'c[�֍'E�K[ut�^;i���Vv������M68oL*h��A).�;��a׆vg�"v��٢HU��|5c#e=?[\Y��Ĩ�i�LS�v"�( qJ�X^݈r
$����{��uGO�AC��~Ғw�q���z�	.�Φ�������eI����8x��{��hg���~&�05R�6*%	�cO$�l�H���\��K���J:����rh�|Ƀ*��N�VF�|�}l��]�|��w�edFK����aU� �����	Z��^�\3p����}�a Iʐ�����F�0:�kT/�T��f�zȸz�!��No,d{����"����4A�
lȍ'�uP���<�k�m�₩��*K�t/M=�AE1������ĶH+�y��ƽ���H�2ǀs0D�]Dᅆ�D�^1�7����3f��Kb��k��P.`���EM�H���ӾBƵ��{�ɟ��Q��T�W+����c/h:�@`���1Z��h7���Ԕ����y��3=p�A�nA��~<�a��J��������� ���WU���w,������Bl|W�G�}���g�P:<G9[>R�n�*B1�vD��[�l(����k������ҍ��dnm�J�V���-���,�n�T���X����L���%3�r�Yf����f�n�s�-k־��s����7���gN�YQ~�;�k������6C�J{s�f�1��q�	�D�8�h�bNJA,ßD:�s��d�u��ϽɏO��T��Zn��T�	�0ˡ��N���/V�D�%���EL��C�1���>�^^3B뗈@��+�����F��TkT� ����mz�������|	l��4�kְ�(�[4y�[�|%�4��*Rv%T�'��$㛗7�R2�a�j\��^��s�]v^4�k�g��۷�pI�n���n�@�S����\�@犰5).��p�	� ��V��6�#:z��pj���H�z��Hm�;�����>!���L�U�a���s<�q�V'
�N?.Ջ�@0	Ź�So��*�g�1I��e�cE��٭A�CY�`3�R��P7�z����If��(�HYlӖg��{#S
35��	���G�)�]L��˭�ԑj���%�Ѷ����n��g�7�nJ?x�`Jjd	�e�Oשz'T� 
8������c��v�.��H�l��Y�ʆ�Ho����)e���W���g2�����d�8�"d0%l""�"(�Ǖ�������+U&��T�7�1Ai��k�"ç�G�Sr��=��8�F�Ø���J�WO��N��R�$ۨ���j�\�I�O(hN� Ʈ��%60~4��&	��v?��\�
�� ���3[|&�#��g	謄�384Jb?VA�����D���{:�);C[e?V�Y�W�1Z�Zp$�P������w/��e�n��C6���{ �A�ݥ8���H�DF��9HG�����A5�Z��a9'��w���W�PA��t����tN��5k�"f��TJ���D5�G�b��@ȑho�7Mc��x�����o��N��E��k��!=��3ש��D������z�Յ��uخe�
(�=�E���܎�!w�y�3����w�\�vi-�g:g�/�'�����d�-�8w/�KJ�<\myt�-Ϳ���r�'�7A��VY���L�Z"�c_���k÷nT�P�\���-�kf�xUG;�(��ƍUS~<�Z�.���|;{jPC��ƣ�s�HVdM'��MB�_/^���W���+3��_}�O�^��i=S�޳4E�����(U̈́��u�DH�B���dl�BXy�ч������CO������%4���߾�w3���>w�s3FR�jw�`�O<[T��W���"¢�vly�[^z�oF�c1�{@��pFAʉL�d��{��Qd��&������������l�͖�f�b�[q1���9*R��pE�oJKKۑ
����/>H&[���:9<+!��l��0��hw��_p�V�%˲�-�sA""h�袾}�CB�l�K�CZ˔=Po������%,9Ev:H��D�[}�nA�K�3���H��)W�i��).9-�5����1�rl�ID�B%�7��)�37N\(H�(F3�ƭ�F��\���?E[�ow[�e,�&p �wE�*���� ��~�SV_Cv��Kuݚ�
DG6�|8?��2z�Ѱ�UG�#���a�MʟNp���e���ѝ4�n��2G&3���8w��^d$�}���v�+|4�YӰ�;+i���d��PT-\���#�Q�x�ٗ���`��)(�Tg� 3�ʊ�z�A+!���?o�w��Y��RU]��~Dy���*�T�iyy�	AУ$��WG9d'5�P�^&�FJr��Q�o��v�af��$#�IX3ׇǚ���Ը!G��� �pg`��T���r�)����֔7K��R�'׸]�G�Ij���O_�>1���:Ț�z���cv:��X��zvv����.-��֭��L��y%lP,<��E�+8�b�%1Gr��E!.����C�J�\�.Oe��k�%#9W9eA�	1�!��r�!�o%�oiiq�nݎ~C�M9T)NV+''�lk_h2��?&��{�#��?~����g��A�0B�ĳ��FpґO��?���dh�Z�֢ib2���C����X�w����w�����Z� m�JfzI�������Pof�jO�lP�^�� �Z�q� '��ښFs�:Ӻ�Ie%�O�T!"&�cх?���op��gA�.��r~|``II��驻�!�56z�k�ppWR�BF�֊O����p�\��fh�o*�d�R��3��{�?Z�_���W9�����=�w<��\���5�Q�
gD�m%1�h��:0q������0��`,H������|�V��W���������v���;�͛\XD��1�R;Riٔ�W���̍7��~�{����pj�"�(��X©����i����Q��"Ʃ�M��u�\'�+R���X6���i�.T-�ߟ?_�94����{��e�׮��[�Q���7�{������n�,��]T\�M{��j�����k��<3�E����&�]��4���:�(�!Tr�L����b���F�����ip5U��j��-cPA��kHa�%�nD:��/�HX1	´�}�뺩U�\r��eOr����Sa�jX��84�|ː[Z{�_���I��:��X���q�1dR��q��,p�J���״�u}��>#�Šw��O-�.B�CU.�e$2P�!B2��<b��H���'vp�zŬ}e��u��`	��f*7�"�A2�;�B^d�=o�=�����+��C�^ ��kV�;��g�D2jr �O�����}d�d�(���U�%(�����?�A�u�����9ym��0���̈���+(�,ɓw�(�HN���wW�1�f�۩g��-��E�P&?�CuhTR:5O�R�Rґ�mw�I}��&���ީ���0�A`#i�q�X�����A�L띟4ܯ[r�^����ގ�v���&*�q�	�B�P�Ȣ��G�׾���-��{�#�y���^��V�z/0��_�R�k���Q����k\ �;����o��&Id%^�M�L��O5z.Nڄ�p�R��dCBL|���^3�A`Bq�:� ���N�	0u�dw����0&�Qu���Ε����q�_׌2	�(Ќ����[+N�6����O�F=k��0���>x�����r��L��ܮe�:Bg��h*J�{�'e0=P����t_a���Y3쳭{���}��ڹ���nZvS~�����d8�bƋ�hSᔠ�n���C������:0���_���~x]�;��eG��hh/�2I0�b;������ho�\&v+����dc˅�ҫΙQ �_��S\4��Wq���k��p�W��'�VU}����OMR�+�("ũs�\s�9Zt�\�xxcNz��Ғ��%Ӧ�Z>���tk���1��B�,*A'�n��0��W����IS�B����>���Ol����uiY�Dd+l����g}���s�+���������ޜ֓FO���󗹅kuu,�(J,$����s��V��@�B0P����a&[w*�t��ԓ�����������/�r�ht��R���y�v��5��wf�CD�E��V+pu����Y��x���R~.� �[��}��0fs�ka�cc"$�؄q�d3���_}����}�M���h~��aHK2C6� ��]
��9j[s��*��Y�S���[FLNr�E�=2���T=$��J��D"/�������Е�@v��]�h�kD��Wt�cp����v���G0� D�"9Y�W�k`��g�aK[�CqX�d�2r���&��q54��Q��^�6>>ڕ�^6u*��X�N��@B>�~�	@��p��!�4��p�p���\�~�/�������!G��2j� iF�I��!��N뜐����͇���E2H�Gޠim�瀊�͏
��P�3A���YP�U���n��p���:#�4�5���>լ�>�i
�ۃ�zD	�B��7�@�~k:`b37iP��K���b���4�@f��!�Gl\���R�����*c�+��+��R&��<��v�׹��']z�t�ͬM/�V����qO?��H�K';|��I%��lV��}ݽ��~�|ꪬE�&�q(U�����=x�}�k���<)���	Д,��ڲrCU��S��Ȟ��������{&���`~��z�U��T��I�I���g>�&>Ҹ�O��UU���͛�%�QD�%HT�? �^פZ�<��x����)���|���;��OB�ޜ(0�����P�M��Sc,;�X�51�v�o�y�D��L�S`[:�̴�U��zWIL{Pkhg-H��`���vT!+.U��@	�����~�+\e �^�5H=X��\`����HT�Qv�	�>R{��"�&�@�v�^�k8[�ѝ���2b�$Ν��0k�<�@��i�*Z��=�K��������O0�|�#�A)Ŏ������=�N����X���p�����{�G�A�z����'��W�����҂�!c����?��?ϙ�~V6�QM�8���ڐ��z����O���䩳��ܤ���)��L����҆SBM;��a��N
�I�0�&2F�c��>j�����p�ѱ��K��`�+��wϞ=�Vn�˿��G3�ˮ9s}���e�6nl8u�*��_t�y��Ȼ���.�.�$���������;�>��T�[�����2����N��N��:/�ݺ����|�n#��wŻ��W�0��}��B��������"Z55L2���t���@�[8(����0�	��$�l!�q��hk�p;��ۯǘ�� F�iJ�9�L�ǔ��6�[�C0�Տ*;�L��f��}�=1l8��2|?��k�+�Q���^��+�#�3Z��'%TŞE���N�v�+``������r��cX=��މ�/���St�c �)� Q	AjnR��$�=�A��U��m��ܷ<I�b�W6hC�����ȇI{\C_�$e�,ixEjb"Ӆ��Ӱ�g� ^��Y�x��@��?w����M)&��_ޏz���Xkm���8`Q s�|][d%�9�h�#<�3�IS�~��q`y�=�S��;�yRt���Ѯ�l��$���F8�;���,�Sy��{l����K�}���h!`<1��dԑ���-rVR	50e ����(��l�� ��S}�Qd��3Bӎ�>@�F��͘|�]owk�S�l�f�)g(�LMOu��%Q���ad6Y4��QZ�o ǦX-��=o�|ӎ/G�����srhZ�2�<��O���]�齇@�`��r��'��;�YiŸ83��>��O�t����+��`z�����2��TU��a�;1D�ߋk�����h�χ����?ϗ lx��R~㚒h˧Ai�$A0	��R\`�`��>��F���*�:l��qg��X�� @���s`���� �B��5X�����~Û^��f1=:a#�D�T�F��&,�-�"�vN���\N��l3@��q�E|�-�x�`��O�p���~���_2C�������ϑa�;'S�l�&���d����c�]��������|&��,.#m���W޼��v�s�ԑݱ�X�1��c'��3�^޶oſ��_��/�Sk���i�ň�[u�Q� ���1=����Zbb�e2�������i���W	b��նc2��־����ln?q����_>����O��gAI٩�Ĩ������j�-6R�8H�	���o���V @�=���L���-5�{�c{��:�iE��;_�hyT��V�c �|L�&��_pM����{���qd��8`�S2�<��P�_�X2���:܅Ín�-en�B�T��֝dBs]J�H�{j�Cc=&�*������$�����vˎ�1�2�B&4�54J���p��;��&���g"ֶ�;lRY��2^�ˊ,(2))����}��azꂬE�QiD`�eds��EmP9���^���%jy����R@����&+�آpi,�1�;͙�����"锁����^�����q����nf=��QUM՚M_�����[m2�7�A5mS̒f���E�g��k�VL�S�.4�����p4��5�B�]������[��*�Av�XZ�7C�x���j�S�����gB2
�T�V�:� �uk�
��ҵ"�̩�2����Ɍ��/)��f0��r���/a(�K� �����fj�]�� ��>[�ד&�w 2���$����n�O�7����!̷�w�.��;��k�������"-�9��np<2В�նQfi�0r�ܿh:N���ӽ
t.f���T־��h�Zr~~�w�����?�=�k�`4h�A��vg�2gO��K V��ήf���/��b���K@HY�:tp��y�D�|�#���{N ����g�oYc~��]�f���k��U⒞��~i|�b�N����/((���w
qRN�ដ��d��'=�հo���5Z�k�&u]��s>���"@?���k0��!-��<�H��L�������8�X�fI9;>2�u������|_����p-"HJ��������4���������\��w׶Ƕ����(̶�B�8�����1c��[�.�N]m}V"_4�Ųe;q�?�h�W�9��o�c5��l���fiT坷o¡���<g挚���∴�F0��@��̾���ގ�X�V5���Q��l�M���|���~����W��_8��������޶�I�yG?����o/�ܙ���s`3S�2��l��>%nٲ�'~�3�'�R Ƙ�X���
F[
֣��\�u/���f�_��I���"���}��K���{��<Y5.�g��2�����m�t�d���?���1q��^��^w�x�$5�9��umd��ze<CEna�M�T�i��"���j��oҫ�Y�h���<�N�L�Ȃ=AI�'ܽw��n_�]�&`x��0�q8YҜ�������]����{���2/�<��Cr�����j���A�>K	%�9��Dcҫ�M�8Aځ,E�S�!YE���ײ�%�{��	��E��ۿ�;r���}��u��\/,*�XJ67O�����߼<�[𮌥j�m��	(��yw�ȹ1N�R!!����]C�!iJ��8�x�u��a��b�
����C�Ը�4*�+[�p�8��dP�8�֋��A�����Q���L@&L&����g�s�#�<�w9c�$���	��g����f�tF������Ӓ��ʤ����T���1tڥI_Qq� ����|���ƀ^�q����r��-	���1�J6⨈��D�搯Y��2J?��K�F���A�������ȴ��> T;�[^�sb����Ҭ?p8�{�&��3�G~���3�3�3�9��O~���Ν��Ռ�����e{�N�M"�^u��sM�Y4�X�>?:h)�4/�{T�K`���C�LW+���{������{���6�w�@&���2
IR��HB>���3ʸ���M��!�����R���Y7����_���Dě�)�s��
����y.��{��]��2y�_�O�N�3!_��%--5�w�X��@�aj��O7>	S^�^�#�>��3\�����Ͽ�����2����3N;�W�Ξ��zj-�@ߠ��ё��p�K񏪪���T��������{�#�!�בНR�H��ַ��9-#������^��C�i����MIK>��AL�}�jX�a�����g��i�$��O}�R[Ow裂3�Ǡt��������Gz�]ԉ���;v���<r�_��+[a-֮]-���O����cz�=w�U0�ET ���QF|������W]�l֘�|l"d���τ�rV���ب��i��A�4�7Xꮵs\Τ,��1�z���8��"�S>)�L����p���Կ��w<�=J��	�̨�L-v���Ĩ2qHvXr��(2�3���M{PB>u�8�;��A	46Q魌��]�����LȤ���5"�V�J""]�(w�o�F�ζX�2r���>+�4�֭^��lXA�����$Gi��2 �Ո%jc�Z!3��� +U�0��\c�ڠj�F��z�Eo��6��ۭ-��ޢp�e����f4�<�&i^5�jӦ�����YG��fC�wϞ=�L�6~�`}�6�FY�^�.��� �r�T|��`�y)����K���Q�<N<:8e�+���E���8=��%��3��ިL{��Xr�1hZ�%�ԙ�p)������_f��B��1� J0Ă8k��y���=���n2#|�A�w�(�Q��>0DW�iD՚��h:�b�~mkk�\C@�m�	qe�9�ᇧ0$����ūO���\c��MM %��.gv�:$l�4(�s�`��ѓV:�v�8#&��	�4�2@rj���U�>�q&��*��Ⱥ~�7>���Gɐ����+�.*�B+c*��,��i�;۽����z�Nr� b��w}��e�Ɉ[b�|�F����w	7^	~ƍv�,�z����9;��J�\����Β�}��xe�
T��4зn� 7`��L�F�t�>�"$���t>����n|��k�������]~�:+@�#��C�"1�`���'V/�ɇ�q����&ȉ�Hj��Hp��h�M7` t�����N��?�C��\�{�Ё/�޹탘�X��|@l7A��B&��$��lmON�ݴ�ɿ���_���̰H�ȩ~��;rh��S�������@����^����-��{2#=��5Fd;��ۓ��ֱ�:����ֵ"<��#�BnF�w��3�Oi�;��/�|��0=+-2s�i��a���iv�����,����ܱ]���eLHYn���7_wII�����Ԅ<�6 y55��О��y��[i�jIJμVG���Mݺ��D����˱��õ'�Y�:
$^�8E���A2�t�@����,,�N>a�9U{]����a¸��}�m�\M2��R�PVB1��ڈ<��$ �q�޼e���9�|o��L�2��=
���^e��(��Q�����lF�N.[��L��\�H��J
V0�wԞ�n���` EB��a2�11�epY���ϸ'�xʔ�b�A��^�rT���1N ������_��k�9L��T��D*:y�4����c3$
,��E9dWu�,�0l�	�8��h�"l�gm�P�����м� s�e���	����'�|��ˌA�[u��E9��Q��*�㏗�EL��5s�	��#��R�C�G5�!�Æi���7��QJx$g)�H
���������K��`���c�]�n�Z����y���@�	��9���͜S�֭����Y]p�g��������d��R4��^���P��IHH�c�ͺS��"��!�o7s�(#�E�3e�1��r|�9о�ǔ�0~���'�E X��A�H�J�Y�6qL���$������)���R�H��ܿ�_z�Ls���b�q�^�>�K�6-`^#�g$Ǝᵺ./F2���{ Zɐ�DbTY�j�:��<�d1���R4XS��s�:�`m)j`�.�̃Y��v}G5���w�>i������g X��=�x���zv��uh>h�����]�`+5%������$��I��s��A�Dn �齃cP���=�5sw��Kx�kݤ�ui�0$%ܤ�w��O���2��Z	�5V2 nJ��JB�|�@�����	��w�-@I��h����*J?3�㭮�W��j����g�`뫯�����.զ1(���CʿGG�fػ���vn��~�K����-$����t�b�ࣼ�d��}���!N2ƳHfRI2��Z;W�]�\�Ps��ߏ�qIhB��z�4�A�UE.V���?����s	����6�l�'��?��������a�[����M�8G��P��a�����r��K��L�F9�޾��o~��4oBg=��
֘˯(?����u�z��?���K5�mۖj}9��,������*w��񎸤���I�:£B������'.�
'K][�x�^��>�?R���.)3�ѫ"�D���n�p��[\Ԉڷ��#�1a���cӐ��4�M'VɟY9GK�<4�g���O��`Ť�D��1�c�]e$�km�\%�6�0A��n���3я��nt��_A�b����U�/�:Aj@�Bj�2��떩��Q/]p�,��P�C)�H���|�9z�֧}�Z`��q
�LD+���u��T�iӦ���1�]uj�J"u}������P)`'臓�ڭ�J��+s�������ЦK)S�3�eP���\�t�L"e	�����;h��>[A�i����8��V�´w��0`�k�S�h˼�?<����BY����V/��u���L�D"�\��گTJ�y]���ֹ��c�6,�1d2�@��lHl��� ����S?WQ�wX�bB�y�8� ť%RǏJ��KO[�ć.�,�w3��8�
�C�]q�L���/��xa�wJo]�ڜ�����T�Nब_N����}���5�8�>�`+%��r��fJq0�!�}�߷��B��[&g�Y�/!ߕW\2�U�5��&ҍ�~D\ ����(}0�S�0��,�������6�򒜈lE�!�>L�	d���(oU36ֹ�#z���x���ށZ��� ��g*E�{����c.��]�*E��6e���Ĥ@T�bn8#���~���m}�����Zނ�8�@���5�S��'��/�� ��i�$�R� �vF����N��D
�`�D:о��7����D�(�qx5F�3�v�����_��~����t����B�ٿ��a�^��d�J!�9 +�lZ�bO��Soj��d}}�'��nSkiF9��;������mZ������N}x�ޝ�9>Z���(m	��d�q�6��֚�jl!IRm�st���(Y�j��v�������q����~�>����߳��]Å��2�*�h���w�̓����s'/����'����H�`[�h�nA<�6�r�����-HH٪�j��R���҅�������g���a��٩']Aq�S_��w?�YP<T^��l���W�ۯ><
�H�I�`��ܕZ�h��$�0||P�����rᴀ��Z�ɚ,<��(�Vr�)�f�����\�6.���9,YyE.ֶ�-֚'�o����D�8[�z�J�q9m+����N��	�A}�w�}��@�v/�RR�^�D]�8-s����m1�k���z|T-5<�:�}.)V����m�ի�[颇����Gql�(Jc;V�`E�u�M`$">������� =�֏a�8F���9sf�^�AF���Lf���V$�a�6���Mb�
�N��ZS���$����w*a!pL�J {����RUl2�%<Z�4�� ��?��"��u�J�Y\��0�6���N��q~��)���by{��w2
���`Z[\|6��ͬ�������d��Q6Y*�jD��?kI��w$�w��'�� �\���QY�6}O�p�Y%�
� x�v�E�U9E$F�4����Z��!W�s���ر������<H�M�~�G��!��ع�mܸ�z�};3!(/|����Ν;o��W�uHCA#Ysɺ�P?�0Բ�� �yY_%�J$l�{���E��5���W�.4@vЄ�<�o��@Vj#JU�#�\�Q�����L{K����q�I�b���〳��GLe���$N	�H\(=#���[�����i��x��m](Μ��!x���X�y -�V��@������ު~�9:3A.�~��7�ɵ�2�P'��&�&VJ%��)[�Ec ;��)�����E�1��T���lk���u^����MLL�_Z?���?��ܙ��O?���}�w���LM���2�g_�����E���uK�zd!�ޢ�OU���0�#���K��J���n葃G����@�=����ډI4��Q�G��5���^_�%�*�>!��sX�`��s���~���<ulWԷ���j�|�}c��0�UGK+��.yC�H�@���0�/(4���g�T�mj���~h�i��|��vt"2�JՅ?��:{�D� 5����dr��Χ��:�t�U�����a�Q[#{�t��������?����?v�ԉ5�^}�w�x㵍W�4a8ꄛT�O�w\�g���%VƆ�\e�穝� �[��c���1�B��`�-G�+)���OP��#+�OB&��=t(�1M%7��H3���^\�1�Anמ�8�Aw�m�t��Uil�7�m�n���=�c�B��׶�y�~��SO�cWݽ� Ҥ���k@Έ?xi���u��5�Z�p2�8P-@�|tp��=��A�-�mh�4��m��������}���k����^��k׮r+	�0��lX`mJ�_��7-[���%��֬�Yp�&�i�pX	60��d
W#�51�κo^>�r@�L +ʡ�A�~�qX�:Q#�UFفCڳ�5d[�����a�t
���D4,Yt �!`��i���4�5���H"8f��P%�Luu�C�" qkXH]�W|���1�L�j*VD���=Qmݘ�j��{
Pf� ���#(9���#� ׺/b����eΜ��\#ߩO[����?�ܳL?���!lpI���j������$��>��f���)ϰ�fr�Z=9V�o�@+z�v&ǭP;��@{@NM�Q%0١pJ3Hӎ�{(�U����M�tZ�����3�'Pʱ��0]�j�7֐�5,R���x��+��}8�"K�B;G�g���g����=p|�%���x�����e,s%��nk��4@T�RO��|��}eCo|�Ll ����͏���>,� E�#�����%���(�^��Y����A~@�����r"�<6�M"Gq�������N�i!�����fp��� ������1m�����;�����©�C�Z���������5�{橯u�G=����ir��x����@W��<�������@2����\A(#����T7�讻�r+V�t�-�cmn����~���u�Z��9���/_�Tv���ܸȡ�	�M��E+JeSϾ�N�.�r�'[٠W���+B�B
G|�a���$�8��"�������N�wU���J��qFj�g�e�������O�݋U-OY����U�n�q��[�Ӫ�����,abT� �"�7�f�`��Q;��֬���l�2�<X�P$&�"?]��^y���Ѳ�Ҹ���v%e��e�8�.:�5װ�9 2$b�W�T1��ו��Yf <"�X�X��J<��
my�%H`��;��{� ��P��̍Z�$�(���#8P����̹��~�Й-�>;~��emL���F=] ���0וΰ��Ԣ���Lx`��fM+���n>,��<��aF��20b�4C�8P�3O?��k�u7����j����t��1N������݆���\c����	d~��O �����L]$����b@��v�b�5���in��)�t���4Q��6^��ȝ�)pi�A~km;�*���9�bP�S��԰̿�}E��A!�ju�et��sf�^�%�d����C5�L�P"I:���0�[P��l���ڪV�;�ѱ���V�:{y�H��a�r�9���?�ᶾ�
(Ǹ[�r�K̤V��J9O�hDuU#s�k��K��Ì�zUu�m�O�����B<)�	Sl䂔��^ɩ�R6�0̧?�9���]�'J�	M�*t��A&�j�"�
�Rq�Vٟ>�������Č��O�s�K
������@�XC�&�d��e߄V����Ӹ^j��R{�u
pU�8�k�}��il���Wף����ĞH`��4+�	uQ�����gm�>@�
l���wÿor�:���e��5ʪ�������^�}��� ���� j�� ��ΔX�xU�ә�&5:�&�tOeJ� ]��x8o}cm�~��$�G�"�������/�����C���L<v���jk��d�Ƕ�E���H���?r�7���gD���X)S�ٍ�$�Z�y���>�43�����r����V�i
�֭"���گ��B��%� ������J�ZA�R��8H-�D{�m��]W6P<w	�2��ɄF�T��m����b�����PH��f�d���jL��h�{� ��⸛}����98�	� �w�,|(��34c朥.=������e�q��|��+�ZM�R
��&Wa�Mv���=�㖮Zc�$B��&S��
��ƐKKH��������=�k�ݾ�RAT�z�)�01Kv~ٝP����%�a�h������?誮^��B}�q�EV���� ;�����h@�bf�-�2�̌1$q��I�w��e���o��I�4�8133�dɲ�G3�����>��ј��������3��~�^�g=+3yØ�1>먿��O���%x
�Ѡ���L�f�]��ٖ���b=�9@�^ڝ��q�k/�V_�rE!���o�o��ِ�M���s/l6��ɟ�yh�{� 2�ht��D�T����H)����.C�)��r���ܹ��i�Z��hY�x�s�E��BZ�Fs?��O\����|�S�Z���FS��*��tK�D�%�0>�p��VHk���!�ȾF7�.��qoj�;+~�nF����sP��[O��*��،聛aP+���D��JU:ɠ�$��Ç�)�1Uow�)�k�_��0��V7�J�F
�~���t?:	˓�#}�ѻ�w.c�r��ጢ���a���G2tdB��mb|��i��Q�����V�C=� �p���Y�j����2žnҤ	 @W�>��|_B��Sڢλ��e�G!6	M({*�G�{�D��O��"�u���]#��Ed�A_h�����&�(��~��i�x �ز#�덄1�^/-6[���Y�C��Kg��WD��݄��F�U��4&��6K@c�|$A�DJ� s{�葘�����X��y+o�˂L�N��G��78�f.�u�ի���3����%���BF>񨍁��Ç�"�ӱ^Qr�E��V��٬=s�S~���o���П��3���<�=���P�*6ev���UȠ|��������Gd,!JRO�l�O@������?����_����/�{�>t��?�������^7 ��4{����׬Y��	�����!^p�Ei���x��2b����<6���Xt���:�=��Cns�*`���Q�52���j\Y]��֦����:��w��T�yQ��㏦э��	��N#`,�}pl��;�Ww^��	�m��thǕ� {8!U�i?p�u��ݛV �Y�J��S�:ɋ/�����lj�\v���d�f��������Xt�]뒵��_��6i0��>�������߇��ڂ l�h7}�d��ӏ���t�r�~L�Na(P������d98)�4n���y��1IIKP��$��q�Z�y5��M3C~2��!ʵY��m_�'_]�$=��a܇���4�U��E۟=��?�R�J��G?r]�uŗ��4�Q�uF;�)x?�8��л�2��9�V8Y�:k�A���f5�����-~F���u"eJ b���08B�¢77mX����[a�����d��t�yW (4�|n)2����\-V�0�@g��De\�Cѧ[�O&�ݺew�6Ϋ��#{^��_߱���< 26IC�h3;��ѵ��b�!�C0M�I����݈��^X� ���Z�	��}k^�~�dB��9��(��*�/�2�u��<wo�hwY.�6z�z����8o!�\
��:�Vx���Kg�}�4�b$�Nۺ�S��L�-YrzLBB���gk���&_���:j�<��;���Ǧ� ?{���q3(�����g�J��<�H�6�	�2[@z�QF�~0J5y�W�C����\�rg���%�X�,.SR0���C�z�"Kp����r�PJ4iR�ݳ#�&R#��g��M���[���k(2~?���{�=P�>�����[A~áNy-�>O�S>S��VJM(:� �B�yɿ�{�u+��EPQ���ρ���?���1���d�O?������W��k����v�A1�>�2���_Bqf#�K�v��J/�b
�	��Zj@��.��҅�'��S��w�}��_����1k0�C���1$]�+s�.�����_�9U�qw�Y\M�Ѕ�
l{� DǜvPCR�݀%�F9�N�y��/�<y�eÆ�ڎ�4�Q��\hƌ��n߳���~ځB��l�;��ƞ��s�K����'3q=�ԯb(
f�v�:*U�����މ�f�|@�^��Lۘ.��tڙ研W�H��t���;����0^BTM8)u�uh;)A4�+h���5�,��qH�f3��������6�)4����F�L��s���N]�CG�s.�.&w�@c����F[.Y�2>��gH����e�/:�T��EK��p���B�,Ò�q�x�����X�-��+֮f��]H�2���6��]���� �d8���/��:��W�3��n�C����_[������M�5T���{���0���a��C�6͚1���qr]: ]{�Y�`�p%��pd~��ڋ_y.�^�T�>u�!d��e;}�����nJF�C;}�<dui]1q���+�&�5���>B9���\q������[�&kfE�n@���!��qF�qdNh,�@YRRT�����GY������Y�*e�ǘi=6K�g��CT��U�l�
��4k�|2�q!<C��s9����n�����_�z7 �6 ���j��W�A���I'�C��~�=�!��e�����nAp
����3�3z�o��fV�+��\��*����7oܑ&����ۇ�m�-a��ؾ��oq��#`r����c��_C��:�ĲN�㏟O`���q���m?[i�\��%;)x��4J]C�R�^d�޳5d�zchI�C_�f]<˩����s��l&��RH_ʿ�px��|���tk�M�r�/�Wq��_g��������j֭� M�]���=r��}Ӧm���Zȷp������e�U\Û!%Zm?�`��.8�/���_���u������yﮭW̞����B+������ʇ�����^qDn�U�DD�f�ٙ�\��c����ٽ��sN�:c���˺p�qwv��zQ-D��&�˗\q9K`�*��L��>� U��>�`HD�5�J4��ɋΓ��}j���ҵLz�ٷӤ!U����~�c�����K_ya��=�PMm��j�G�R�Fxx3����,N5�֢��Fs���e�M5C��d��~�g��N*x�ϕ�̨�_:��h.wp���h��X�^�vd�%/>���'�rd֢1o��V��1�+r1��M�7��*k�\���k���v��@x�QCfI�e��&~���}z��S��W1`��lJN�T�b�[� 3~��B��˄6��#�!�MLS�� 9mK���e�T'db��F�{��%�x���讏
���G�g����7B�۷oO�w�ʂǩ�im��Ò�.��Mfn���KgR�v�}�eY�=��gp0�y��\��d�G}T:��3A ���+N��HJ3t��Q9Fֽ���t86�P��z�1r����d�f��6?~�%h+��B��O�1�uϞv2�ᐛN��H<w��d4H�rj���ǐ�P��%1O��vb�~K�Kt�N��]������US�A�Ĵ�hC��ؿ�A=����xF˹V�mx���lO����f��}m-���H^yie?zƸ'��1׷�R��W�c}v�a������%���&�����0M ��}� �:1�*��O����)���ש��Y����Y����c�2B:uL髢T�i���> 4H"���N����q��yW@�C���znf�c?�z�瞴���(�P3�<��$�V(DXԍ h���>hMtv��6~��Dr+���V���^:�=l�Z�,����IS�%tɒ�A�{N�����U�Ou��	_nֲ|�@����g?����<����&�����<o`LcT�a(�W^y5f$�b<��7ϕj�f�J��Xt慨Ma�ʹ
~�[9toܸq�Ϝ>��yT���k���}��r�����_��#i�9��b<d��HU� Cd���K��G�('|�)�t������҆�.��4�&{��3Oi㺕�?i:��}_�G�ݽ~}�d��/`����{$	 Ӻ"[Ua�=Y��P���@��L�6�<R�Ķ0݃���J���X�3����G��͜�W2w������K�=9��d�d��/z��i_W��bn�6�W#��@�:1=�C�̧a(��q��Lm��R�.D�xJ����8�p�����!�SЉ���߿!�ߵ	~��x#:1�Q�ܝ���������1uh$�[Y6)��Q��@�9�|�!n�Q�h��AiŒ�ө'�������1y�|�[(YH-?���X�)dm3��҉](�2#�O�Ӂ��=���n��洖�}V�*��wؐjD>��?��4r�ܷn�X��cn��0�p��~qu�͋���}U-��Ϯ#�C�!���6C����MkI��i�������B��Jx"@V�y���"��� ޵ѻmX}�3��6�뗨���P�#��+��[p�Ƃ´�����!<g��zg�7�w�����Ӝ��ʅ��0����c���օ+*p�:bZ�"�����qP�)s|�F���uצ�m' �	2 �ξ�<��0c@&|��a冀c� ������D|-��/՛�o (\gҖ:��uuRژ��Ю~�{>|jZt�8JI����1�uo�J��al��� ��@�S���s��}�$�ֳ�׏��繃`n$��&��:xd�f��V��޽��@mAZ4gb14e�;���f������?�^0�����8���u:�1(f��-�`�(aR�ƬY�Q�;&Њ�
M�#��ޑ/(��s��YG�����N� s�H�#��f���F0Ȫ-tJ9c[*)w�j�-g�CO���;η|ˀ��i�Q��j8ŗ{e��?���O�vE���i��I�w3zly���;~������������U�Z�~�w�&L�ٹmkZʜ�%/>���HZ�a�dF<���"S�!�Gr������Jd��n嗽�p�>�c/j�°��o�|��Ys�4wމHC�������N>�4�g��z������p��[W��ukW^�j����]�|��5�~MM��.{�U?:���_������l7 ��!��a�S�^�x�Su�r	��wyらs���V���K�|�����T�I�{ȳBe)�@�n߾C���p_��<�X�ބ1i���fu�
]�C��٬Bx5��ԥ���K�q��	c&�Bt ��<�G��_�Z���}�?�޷��1CҮ��Ӂ�;�իS�r�Q�J��\_3P�>�i� �ft���}��t�M?J-;6�A����4�#:||�&T馥�8�1��a �!�l��+P#
��(��hC��E����|/|�%�?�%��T�*٬�����8�)�M�pv&Ŀٳ�b�@V�+���@��?M��֖}-�{�!���S�o A�T}��k��۩cfiq�:,��p }I,��ȵ��t�|�!-=���,�U81?�rA�tc;���Ա�±ĺ��}�]�<�{�����A`n��w��v��aM�g3�}+Y�(�o	H�Ƨ!����8n���j]	S�IĦ0n*�]���饆m�/�� `3��P2�hWs���뷢���p�����6^K�6�y֮��SL{���4G�BX�
�S�z7�קN:�2-z���Di"&��,]�c�3����a�A�<�k�TF�����{���WA�,3���g6���Qsf����2 r��k��H���������d�ty�C��ᇼrn���NO�V� 2�Y��3vO�p�PI�\�E\_ �ve���,g��םK0��}��r���Ih�<��,)�9����Y9Тn<b1�&®�BP���1�A�����e��5ZҢ�#��8�f�StѴ�/�_�2t�By�������,Sd�؜e��7���g��W~&%E��6n�i$��իWB��Dޜ��5�B���Qr��g�#�o���{둾�B��~>���z��ͷ��0�P��ƍң�<�ƣu�y�F}�Y@�!����k�{�����QS(��a��JJ��h]�YV�鍲�j2��������]������� �`L͚r�B2��l�Q������C��=m����9^|����W~�Y�������~��?&�.+p��0(=u�mi�����C��W��g�+���ӏ=f~5z�V<�2����<$�����v2��PC��Ӌx�A�gΦ�y(�ju����5�`J/��*#s�#�v�˅��m�,��g�d�m�n��ߧ�f�M�{�����t�P���"��v5b'_O����O�������%�Z������o�<� f��u=z�T���t�,J��@D���5uDeD̼G��`�J'g1����:��x�B�-���_�_��`���G(�	��&�2�ޥ�����>��8E$\���<����g_\�p���� ��%��qƩ���-�y�䎊��~���%A�+�H�⾏��py�N�9���ܐ����"���e+�=�Bò���j�~ڢ{!��#Zm���8�ٷ��q0��u�$E�� ���[w��~��((;{����^�	mf�I��N'�����M�=��F���=�H(�ͧ���8���W���ӏ�q�ׄ�-B.꽋� �Q~��� #��к9dȲ�� �.8�;xfk����i�kò��A�'`����ҜgsP)���h��'���4�F9�O��4%�j0�
��s�����q�"����+�*؋C�֧���s��{;j��t>�Iw�q:�5<�Fj�u��u[��yH��MoD�x���؇vi��^�b���.�a��B���)�v��0���c9������\0��Y"t����5�Ʈ�dLHz�6��SІu�6b�M�T���:� C�$b�g��s�����7wI����3H�}�'�v�g>��˲��{7C�vR��l�g�E g$��0\Q�k2=�v�+Db� ���
ދ�x��@����D!��㧞z��og�Q?{� wj/M�2�����2�q��~�iS����`S_�WH8/Z>qѸ����2�^�(�eYʢ$,�}o�(�5��͑��!��0a}<�D�:��m�~���������GG|�cW>|���i��yS�ʏ�����7�t��v���_ph��N�y\Z�ܺ4o��S����뤓N:P�0���h�4�S��{6�ԉ��
b)��ԾƑ'��1v�=p�7R���i֤aԊR��Xǃ��>�9I�ٴ�t��5���"m�%
&Q0� DO9?�RN~*F냒E��V�z!��̣��6�6�m;���$�tD�JS��	L�!�6P�ax� ��R�sP������ӗ~v3�M`�s@ D#y<��>��h3���
Ij���vB��E8�v:Ře�;�HBn��5춊)�t�=Y�&�g�uQZxܩ\�>���Q�L�8n85x��-h�����ʈ�d�v��dJ��:�bL^E;@���YSS-�9[d�y��^
L��/^�*k�L���n+�*��sF�\�SO>EP|V8��f����R�U�o6��V�!hm�T3��9�f�SN:>�2�B.!Xu��:"����� @쿚	?��77��GF����\W���޵(�3�a��x��
�d�6�o�>��cXJ�mL�B�E���A���L!ݦN6*�BY`����EI�O3��R�mS2�yy���WL�����1�R������+H��נt���?�\�|0�� (|�@,|����\�����\*�1>=}��I�>�TZʨ��;pxc0�~&��������SÞ؅`��g��yD�_�5P���c���Q���s�B�����t�ξ��RkTQ/ց�- v�y#\��S���u�{^�	�#��!��̣���` e��s�y�����A�!��9|���H�Nn���T?[ipWŞ�L����K���ǳv��i�����hK�����Ŏ����K��b���/;vP���@~ߍ�w͡CH�c�ɛ�a,�P�]8
���N�|1��9�=!z����R�\8��LnT�4�(�X��w���_��ES��t����H*lMm��>���>��ǟ�\���/�����Ӻz�[�͘yă�>��������WEL�w�䙌��:��2
M��������;���[�%$T�pJ����;�Ԃ�Vˁ}�h4���6�)�ƅ��=��{~�&�Vn�D_즴�C�����s{j���ylν5=��Ҵ�g�ӑ�-<�8��ynZ��#���@���l	�u$F
�&͜3�	b��j��>EJB�U�|ģ�́)��Jz�%���W����5:;���]�]꿛a$Sӣ��R�>�00���C�<S�~�7~r��.*�h�(a��0�Cٯ?ư[3�C4�K{g:��&��[0DudX��1u8���GB���u��Cerv%��l����>��ie�G���/d@����t�	��X�R ���2�D�[C�����
��0gWyg�~5kb/{!"	/�b�	�<Ɏ
������52����P��r)S�|ݠ.���ر5���cRX3Ĵ�F$s	�v��=��������\�5T�
�uS��aėh��` ����E�ٍ(Pw'�l�Dg��kq�xD	*�D&�g@�u�Y�Ԟw'��:@e$8*�)B$��,\4��6�^~%=��3 8�́Z��J��0��E�`�L��|{ث��wȼ����4���-�acg�gX�8y('�̅�sؐ���Q-�s���S�8;m޶�ŽLu�����ĸ���u�CQ8�l������Eu�������)��S�#!�����t�3c��MRgg@'70�!ɚ�P�6$�__���D����_�:��H�,�b����wK��-�?xd�Xe/�W"�eH�b��t�ޮ\�3f���?���ڒ� z5
^�-��c��_EL�]_QW/�^�_~����z������w͡sS���9+�Q���Ԣ	=qU�^~��t?���3O��!B��,�����~��#�ղ����/#?2��m[��G(�޽2_Xy��[:hlzj�9G�@~��>������_�diume��g��k��g����DF�W��8q�΁��z���.i����G��`f��>��+/]�|������0Ҋ� ;�N�U�6����	;f��g��&���;&�s׫X{hQt��A�y�y;�g]\Z=�42D'cU0��ݨ�,�r�Ȁ�)����1?��3/f���i��L����h��2n��|!^MJ�����9�)`�������`�Y��D�Y��&>�l'���{�%�8�Cn��l��ܡX���#f����Կ�實�{���]ʝ�@��������o|3-_�"����*�9��2�w΅�̎�������Q"���+�zo`p�d�!�.�O��U�ץ��a��+�pf�_����c~����ޘ���2?�a�1`L�ʯ������~F�����Pϵ*&�������k�)�z����h5X�D����A���ӱP�.z�ɠ���N��C6��=���v��H�?�7٥+u�8�����Ӓ�n`/>�N?�� +r\��o�䰡�y%�뇱���W�����N��3��<�_w��6u�|:�޼���(��1�fH�	J��W�N�VGR�U�3t]=}��7
�*{�,��!�����c��z'���JO?�T��9QGwZ�)����3N�kq[<T��~F�Һ|��	pSp껶o�39�C"������S֡m��LcǍK����U�a�\�����p~Q!�S��wޗ���al_���@.w���©��N���f��[��֕��J���6v��9�hg��8��":�y��"&F���>�������]-�ߛ���k����_~ӟ�,8E�~�	H� Ƴ쵥 �3� u�<vѸ�@YK���&L?� ;C���.�P���ɛ|~�����W�MO��o���CG��a�b�QX��q��j���+��Oa�7�'�|&͙=���!i�:����E�mDP9���6���pk�l8�m���{����@�܃ ���~�(lM.~������_������[�hЊ��h���}�M��51�}��U#{����!�"6�WOG��%��p;,�|����� lww�
'�1�E깧�L���4��"IFL��6m��`��ݸ-���~8}裟H�g�O�6��+����K��B�M���U�섳e�l��j>/"-�e7�p�3Iif,=�tՍ#�އ��(�u�-i��8@���l���)�b��ZWW�v��N���gd�[�E���M�b���G������V)�I�n��~�`��ͩ��5Uc5���y|�8!���J�{'�T5��8�"'f�	�������߃3�xi�{X)M�?&�Q�vR���W�\Ko�Y��d�fФ0Λ)Y��5�׭G����0��
Z��2F7(C��?�r%����Nh����[�m�%��O�}l&o��h����F��� ��0F��x���,��.���͑�E�����^ ]��@��B����\�3��s����oa��q����7��>��s����d�}���^PF��_x�:5.�g)��h��@����4�с�A�?H9���8rg�Ĵu�~�n�马�L����X�c/�5x�^3�GR���p���	P
��DD	������>n&�l�Y��W�\���>ܗ��g�'�|�}��^ȇ�����:+�3��>Dy ��
�7h����y���R��_���^h����`�pb�� �S�b�;BO�D��~$������C7�q��4��aĩ�3_�rGn)(ٶK*�>7P�����9E�	�}E��ސ�6	a$ťV�Zmj��}�y�*�Z�v`oW^P��H�ʯ��_�\��'Oo��C-Ё��q<q	��3��n���7�����1�� ��)��Р��d>�[�s,Ô���[�8�!�%]W��>1{c��g��L�j�u�e��]s�D)k\�`k�}���"k�jD��A�g��{P��M-�!:jU�����ۘ���s"$��ۿf�!���|�1��s�����n�_����uۆi�h�մ�dm�������~m�ģV=����s`�$"g�m���-9*��0;��zvV;�ϡ��������<�����e/<��:�D���o� �,� �
E�����[�OǞF{�Թ8V�(�q u`}E1�ش�K�����A����xP3}���:�4�j��4�p���=�f����D��}�NS)|}�:Ws��H�R�}����K�#0C6�u�!���x�_���W�<����uiܤR=�gl���u5�Ai�ѹ��EfQ2pAJ81[���GQ��'M�@tBێ������Q��#\��3��	Gn �k�P�{�%��?��G�1��87��ɵ�eR�p�פ�@������9 Tt�l\����i���$�S��۵�$�atI�>���j�����G�JG�;��>��;���N�{>bxR���e�TL�ׯ_��ʳ!�Z͸�O`��3+���i]Zz��z�o���D0�����A��K�o�E9����~i�b%��{�� {��X��N``_��'����@�T������_v\�9�`Rn��2�#8�S����a3��;w���ԩ� .N���.��8?�|�A~:$7l����P���n��D������$������̹?��::0�����H.H�a��x����44�B��E'/b�fs��L2#��~�lں��|�c��Z��1���
k� ����H(�a1K���2J_��� C�)�I,������L;<�SvP%q)I�r �P��od#��K���qc#S���5�2��K�ɛ��-��r����}������;� �@�7u'�Oaϔ�,�:��{��သ6�K�S�LD�RMwd�9X.���8�|q��W���ĵ��a��o�O�H]]S������<��O|͑����&?ϯ�ܵ���'�\�CV+ʿftYY�4ZmG�cLxڿҬ��C�8Zڔ	B��y�-�=����d�@2�����C/��4��k�5��[�C�y�z����ڙ�ۀ@ɘ4��'�N��3������)۷l�a٪��8���,ZB�v,�U�SaEe>�I�K��Q�)����C���OmN�g�H�@�m0˓���>�^���YF�ℳ/Kdo
_C !s���w�_�v�y!:�����5(5'� SS3��?4���v����`��ѾTQ����=�ԾY3�V�f�$9����M�Wu쟺玴e�����vj?��rx\�P�%"#�"�'>��T�D�����AT|��U��l���8�CM@<ck�U�)�&�B[C��m�X�"��yO���H�҉d�TH�W����J�#H�����<=��fU�cNeҜ�� �8u�-���a?�+y����Z[4�|�Y�w�fg�c-��
�}���c'!j5���Z��!{��`�"˓1_���#����(!�rK�t~��(�_g�_p�9��N�:��'f4f�������?�� �9�lg���X���/�����=���gߖhU۷��v�y�F�\�񶜃��97]��\�8�3̘ew{�C	'��=Fg���?���3&�!p��}��v�h%�3e��`cplԤ�׻�l�k��m'�
�7����x :%��P1�����?�Q�9��0���8����8:7z�c�2�ݡ*x�V9�9&�NR�A��-7�4:j��=Ȥf�<�F&�]��1D�gH��l��M���Wv
}�*�C���z�B8�h��d7�[�������<�gԹ	\l/s?uG˦ckW�M�6�WI���YhZ�������Ό����*��w�����ͽ���ʤ����>����c��b72�={���1����޹+��37p��e��Qܛ�|��܏2�T~�=���Yd��{z� ��ɓ'�������k���{^�&4�ܡ
n���ΠYIĒ
�c�?�Q3�O�&�7���1�E.~�����Ն�}}��� yY?��j��y�dn;c�MВR/ꩌs�jӓ�>y��G�_;�~ؖ� ��[XYw�v���Zf`��jSݬD��V�j� ���4�uW�4�������ğjr129zma�(VG����N�̊V=4��pÓ=�w�ߍQ�.�!����z��S�f��Hq���8Օ+צd�*��E�u$��c�]��̝��pP�&���#x�hY��k_J����Y�lluT��b��5 	�)]��)!]�a.Z(�<��0_Z	kW��Ip��L�:5�r������h4T�8U9Kl������8�2GPf��a�l������n��'P��gDXh C�s��Ƴka�	冞��ޏ�LK��@1p*�V�A �ɴj���Ƕ�e�K�@4#{�ǥ�.�����R���"�:�M��5�0�:p���#���}^�O��4�+օc�`��g�@k�Q�qCr<��t٥g/o���x��W��~�c����ē��൜p���G��:Fc2��v���;�����l�>��y�X�(���`ؠ]��T�L��-C�t��ڳ9��-�h��]��M����DIE:�M7�}�.�O�E�^�#��c����y�&�}�_�%m,�TU��
{�4���矛Τ�P����Y���`��n���`3����4�-��y�������_I#h��B�>��@l�kQp8^˾N�e��%\�k���}]5�=���0�YgF{!cKg)�+����~� �=K�$�Y�(�� ?��2s��AbH���a�Ja)D�?f���� �W@���o�����i*M�\ܧ5��	r�AJ(��A�Q�n \M"谫��ѫn''�g�ƃ�VXp��@��(2��� ��x����C//�p���W�`��ovϿ��k��7 �dk��lP��h���q^��=�#f#:��pEC�����肋�M���HU�� 3pK�ڐ4�PFϖޖ	&��[�h��ŗ/�F��܍��Ѫn������V�2��9H:�2���3�U�Ҹ��{?h�?o��n���?�=w�>����������׃�۪zP)�D<�����O����:�1������a�p-=q�����}�$b恫��ʕۙGK����N߯� ��J���F��Zp��s�xbX:��U)�Jtadq|W!O{�it3�|������n�R`������^N�^��.�Hm�tz1`;Vyh0��L��� ���q���d��r�$��������(;��F��#�zn:�����*,������N�ݹ��g��V��?���׹V'|�����!������ਹ�JC��_�f-��H��>�,�ϕ��X��$:a�1�B �ğA���OYQ�P�$ۙ4vZڀl��+^O�wm�������ڼK'�����o��ػ� ��J���m�8���SBW��乬A�ɵEoo+����z�W ����P�+�nuh�N>�D:���(����0A�Qi��I>�xZC0w!3��}�g��=��w���}:�� �A#���%�`ٹR���K%U@�u��0����<�{�C ��݈��f���2���Yh�w�.h��0�|�(�s۠�����)R=$b�^M��}�1����_|5�(�g/H����W�L{޹g�E�er����a�=Z9sCi���vp�� q5��?�|����9W����ٝ���r9WZ��w�:ǡ�@G���� �r�?��hϽ:��v�v��h��kYˈQ�T�{Xr��7&:p�V�3!8Ef�-Sa�"��cɢ��1L�^�M�}��'�@?�Z�*�*f����RB���B�%�ę�,��+�|EE�]����rNS��*�6��N�u���9Q�Ǿ�0l�DC��T�����n��޽+�De�8U�j��ؚ��9��ŕk�����HRTa�HH|�e(l~��Aq_֞�_Ƞ�L+���!Ϳ�n;s��]u�DTK`~@fn�U^{��NZ�>����_CgzlZ0��c����s���
�]�l}06�ٹ�S촼�n�#j:�0�PD+�*��*6�ז��#A�dA�-h1V������������O���{���}��?�觻[���d��T�=�:��R!5��p���_����t�L�q�m��J���D�<����4z[鱬	K]A�܇<����b9a�N�_K�b�Aq����Tr�_x恴a�c�������twl��#I͸j���#::W���nZx�1��P(�hІ4��S�s�ܜ��ގ$6��a��J!�?�]$/�V�A���7�
�o#^������:H��õ�8�eĤ.��˯,N7��'!��e�]H6�ی��-��/�-P��KC"V��:�﬙s�����]ЊN�0j[��S'�
%��C�}Ę	|�!8
��c�c �hzDe�����b�T:vWiZP�Z(�ž�D����t��RCF����V�0C�E�M����f|��Y�[�:յ��\�=�5Dg�[^���,Ma�`L��#��й��w"�y���\}Vڽѕ�9o!�QKھ��pp���7b;����Ӑ:��=��z��X�F8�Zi��?e�t�� %|a�@��͆�α5����[� �5u5�J`�c؛:^��&�ю��n���ȝD_�ɠ-@��Q;Sb���""41�����]��0���ӟ���u��YO�F�&w�qǦcO8!�[��h��+�ԅ��$�z��H�enHH�Q�hc��f�C���b2ƴa�JN�^�͸���Gt+Ⱥ��X��;';t?�`�vI.�_>5�˗0AP9��SP���b^��d�+Ҕ�������o�r�3�t����A8���K���nV^�A�y�#�
'�{��քd�:>$o�=ƿ���Xkc)�<��i��m���;������Wy@��D�b���Ef��c�9λ��n;��{� BÒZѼ��쳛�~8Jb.�h���D������M�R�����*�`�ć��O�W  G:��e���{�
ޯN���7����x��?�����?�k��y����U+w��<���������?��7�����<�F�RaC��>�+_H{��#c�n�w[�"k�"G��#t�C�	�Cx���4����i���Ȁ6��V|FF���@�ܧ?�T���V2��뗥q�:�8�:�C8�hkHC��X)D���hx���8J#� �/�2���O�u�����;�\�\��Q�H�s晩���G�&8V3jY�!��z�ԣ�mm,ڿ<�z� Ed�5�ϼ>]������x6.��eM%��9
��}�}�P�Ӣ3O�33�鳟3{Nھ�3�q�sx�kݿ�9���碳uT���s��'b$�Z5��9!`��~G��I�5���] 9�/��[�u���t�ͷ�=1���K��!2�p�8����������}�Id��\uŁ�Y��K/�(݄̭μ�V�*���^��s}մ^�U(���E���4��}0$���t5T�����@/�<0�x��x��ṯ�ȫ���r4�o4h]ܼyW����!���Ə�A��7C��Nf�qvm�:ŻDA@�[�Y>���}�1Y`�sp7T���T���r]�	�t\�9��xؑ�"�e�`��M��_�)Y��t�1�>����|G[�u�ӣO>�^�%h��E:9�l��	d�3!�n�
�z�$pl���p����c���(v3pV���Cy2����-H�&U�%"9��-}\�>o��)�/�~���/�p��a�ԇk��s5��#.O��g��������\\9��p��sm:s����g:�]�6�>&a�=$Y�Q������<6&�Q��ז/A<g1�G���y��Q|z����b��G�,�K�i��~��1Y�`�c�t�������ֵ���̓/�הj1�,��<}r�tƏK��3i��=i Ƴ�h���L;6oL[!� Pf�Vv�|����I�K趗����%�nF\��G�)B�*��KY~����w�[=���7�لc�X��<��Eܺnc˟+�� ��R�M ��vLԑc�8Z��8%�ht�J�7�:Ώܛ\�vnٜ��/����0�Ih�;�"2UɎ>��O`�G��ٌ��j&�i� "�0�m:yo��*�A�zjJu:s��8/k�fÇ�=���"%:�ѓf�^�e����n?́!@�N�ߺ0����Z��W��l�f�d�q��U!]jFq>=�q��ñ殁G��޷H��H�]?��bO| h>��9�眻(;/�/F��{9������u@f>�u��*j�(��7�:�4DC
"��*�ā��G�t0�4�qN��`=��r	�߅Q�@J��6�������Ȍͭp""�?�pn��R�u�d{�������/���4x�H�98iG�:^vӦ��P�ć�*���\�h��de�W��9�&�āƨY�]�>9H`�
��*U�,O$�W�Ti';�I����`h-p�mk�_>(��0�z��i���Vz���	��Y������d:�� �=�����X��������8ܳ���A��}O�լ�[T%vɃs�I�{�ڢ$(��)Ȃ��^�XG�����X�JQ��Er���r���?S5���1�9ƹ�޻+�r��y��<��ϸ =���i�v��a�H��S�������d�-�C'��`�����K���(G˳�"	
_8~7y#Q�}e�c{�(ןA3*"nؼ)�pz�U�}n��Ò|m��v7��-�K�~G�Ƽ������N�@V�>Dkl	�Й�+�ϧN���rn��p}L�~���Ah�d!3Hl��䒴҆����mG��m�[F�eĪ���A9j%��� �}�9sߕ!,o���C����ؠ�L���N�Er+	C���q!aـ�i:�������@z#G6��58���6m����HnJN�M^��5��fR"����{]�U,V��z�R]�@��-���mظ�3��/�~��9op�M=���uw�O<��vA��r�lf��1
֕%T�cd��b�Td�
<h6l�s1^8��y"-y��4o�0������S3u�5�3��������/�K/�&5��$��rkQuH��������@r�v*�=�����rg��3a�X�zؤT�̘A��S�LD��`��LtL�L��I�0��.�����f���T��tY�6Z�V���E�v?P���Ӫז��z$}��I��M	�b�@0"e�B�#"rk�����5FM���C*Wv{L��p*��1iH:z�8lm���ω���$�^��|��\��B�����h�4*�a���v�(=�]xQ)׳�;�Q����6w��v!3�ۜ9�2���Y���3v�j�\�4���ǡ��t�	�B�̀�u���=�H'�$B{�5fY���b	=�F�R�>��N�r"�шY�W5�=Z�� ���*J]�Mm�$��ԕ�}�_�����tfmt*�n�a4[lKUcf���9	f�J�q.�x��Vz�@|�FԀ�L``Ƅ�C�L4&&��ԲG�3�x���1�fӖ�i�LJQ�h�b�u�ޚ�x(@�n�7������jС�*:R��<�v���;�:�!F��-Avu�{W�A�)'����M ��l�)i�_2�� ����Q����Z��,�[j�+�#Dm8<E���M��>e�Y��=Hđ��~�Q���& �:"���G���*��-Ď,ո��s�<wZ	���Q�zo�.��-���/�wy�T��`Eb[�Y<��&1ޙ��4'�98�xӦ��i��.	��G�]�O
����^;�,M��] bN}hp)�����Q��d3���Y:��̙3�?c�t�����-��_�Ea *|��!я^j�(�43�¡gĜ�#�xs�`Z�{��X��T�iL�W(h�z�vF@	�b'�9�>V����{�.�0S�*w���n��f�����L�9��͘:큦!�`��?���Ǎ�V?q��鳀��1�d��������!�
�oٶ-����j�drBc�늆��E�.�c+�+�ݙ������w;w������h�b�4Z���9����դZ�)��顃;�*ƙؾ>:�?����V �@�kW"�zΉ�hL��L��پfm��S2����rK����� j�Ȅbt���>�|�v�hw��G�� � �m?@�&�/��+m�=>򉏦�����a���?�3����a���A��AJ씬����,�W�.�U"����,�!lnJ*�{�Y�����V���k�,7��Pz����\�5A����j�3>A�5�'����>�B�9aX$:�!�����G{:�ba�.���GB���^h}�rH]�w�7��}Q�*�����k�f�xa�r׈���3H�!��_���n��r��N��dҢ���؇Ӽ9hB`0%*�6t�Qz�@z=��NК�JlB�uH��xh�lo�H�F�F��Ӥvn����p>+�`: ��'U�Mkع<��g��ob0�7�,=�̋�l���ܸ��B0���A�
.ZtJ:���Ys�g�
8�^��������G�S�8kX
����M'�q>*+��Y�.�� ���@�r+"�YNt(�z��a��m�pq��� ���K�|؄rd�H$�~?َxm�Sq/D�xg0�Y릦`��XB_��QÃ�^8G�G��3�Ñ
�l<�������;��/��_{S��t�GmA��P$�ͱQ�L���B��� )/Xx�a�?`���$���~����頣˖-�l��ŞmFslt�1:�n��+Q��R I�x'��~����2y�^���������|��
IԜ9����YZe�ad_�S���.e�30\���B!;Xf�N�ě����@�|fD9��xW�	-y���Iv�GDʥ(���
���f,6kޘ����%-U��o���n�����-�7m�ݎ��=�;� �@9��dT/��2tĺ��AZz����4�Re:����'OO�lETƖ3�0-�Ϧ-��L���)��ңn�� B�q��E!k�&���7}�>�l2I�ɽ���8߻v�!2�[�zE��=����m2��R|�5�S�l�^�����	���9h4&����J\��Ryx�'���ջ�ipOF������.�AtB��k��؉��G?��`Q��:����Jw�}Oz��Ǒ�%0�Q�#W�=�s�^�N<�؀F��EK�D&dH5"f�^����:6N%��u��P*cU8��>��U����shѐi����Y�"1�lpڼ~�ٌ�d���B�1�E|��)<��p��K��a>w̨ ⿴��f?9���^!���P�(�"Nr�mp�k���{"1	G���bFB�>�\�������%~�"<L�h��￟?�Nl�e�w�qX�0��*6�~y2��%�<Y1��H���5~��kd�81�3��_�2Pr(	�0��G�F]��g���F���H�^��힡�H	����M�<|?�A0kU�jb=BHb#>K��]!L� ݀��a`�(4֣�̓1�����D6-A��pvpo4��μ<��F(�;��� %���TA���a*�(�.[�zϋ3h	!�\+��}���,S��5�~��7s����>���.C/޺<)�vZ�Zz�N\o�y�^�=�:���vgqz!�$�%�6H��#e������XӶ4{0�s�	_��d'�>H���G&�|��&T�����ՙg��{o�@���U��{㡼�ԣ�Ѷ���;�ϩ���c��6�cjc`��]-i���h4o����<$2�j�Fr۷o#c��[������e����2$Sdo��_oԙJ�U���`���Lݳg��}{ j���Ѵ��ASq'6��~���i����?�'�f[���#�a^M]��/H�S�����?��������m(fz9�7zbjټ����t�샭�f��^t�l�T��<aҌT3��H��2 '�M��F�8�~d;gh�����f�JDKB0���	H�7���>�^|�~¶"s�EƧ:^'���ĩ�����i7��Ѯ恵�"ř�DvVe�#��4+%$�!�Yݍ�V5�*��^�.VD����}_����1d��}�#��{3�&��ZC�9ƘrB<*���+ץז��Zf˷p�M���LL�"ͺg��Q���:|���� 65sG��]�I�6���Tp�
Y7�k����%��,����/e����rpL�,}U0w�i o,�fP���ǐ���>6 qm�����=��c��� R:邝��.�ʲn���;���$ø�HIÑE���;s<�������fLci�Y��zd:f��H�2f��NT�E)�um�΍�j���G�%N�yH~�$�1��Tt7��U0��bq�o������3 #�����3��A@�
eYB�T�!lv(�;��`�@ ��t�ED��L�Z�1�16ldz
����6F)�V��gJ�^S=��Lw%2��H�ȓ�Bڵ�TϬp�h>o<���R��z���&�a���Ù�A����#���sQE.�xf)>�u��r��HG�[\`.�I������5k�V?���?�#�:��}��_�d��^L�%oc�f�93�C���T��;ĨG�k��@r:���69?�@�ZJ�>��Z������VՂBe[^0�UI�m�~Yj+D��4���O;��I]�������]w�D�K2�ؚ�2o舀x���q����x08H�݋������j�%�<�m���C�kcD�Pz�c�4�@�0�w��o�|��=�:����$	�僕�s�b�ԦV~�� 1�){B���"^m��|��7F
Z��������I�LF�8����}���/{�m7��!��c��*��lV�E�`�4����{קUK�Ng������FEs��i��ũ��iCԃ�\t�1��� d ����G�m�桧��C�(��ņn3�@�$ �2��4��Wu�����T՞��V=��7�J�p\�d�V.��H�6�J��'��u �ҜlA�s����w���Up ��Vr��(�|e�j%�hN<����}k�,C8��7/|��F���U���h�G{��s�3���w�M�0�.��:|3G�-�W�^x0}�#����v+�ݣH�Ψ	b&�=�3��J�SE�t%5YQ#C&�r�xr<���t�i����8��t�y�ҥ��>�yH�,�g���[-�`�jX��P ��׿�6m��	�1��5�:e|�����,=���XM��d��w�B�6H��{�T+ z��d�νi�,Y��4D�g�p��A�y�T@���X�h��^Z�kI����?
Y�Ǟx�䧢?�����-3�=��t��j��B����1�  h�e�$�1ħ��V� YpOuwӹ�b7�Ɩ\����i{������)��6�](�8 J*XOI�V�`9-�^��R�."�lz3�e�V�g�#�F�~�L޷�y�#����H[!r�����So��k�����D`��q�^�e���i�l�Q#�ƅ�f�(r����[.-�W��Uh)_���;}}��k˱�@G���Q�����?�N~h�����~T[½PG��
`����K�472y0�>}X��@��/�a�n�L���?����t ��$ͨmz��^c�O��V�7��j����+'�x���imދ�����3��h��Ȩ<2u�a۬#�"����8�cfOJ?"c8i�1���NK�0s	�v�s50~rİQ�qLmh�nی����.v+D��a�%N���E�����zy��=C_����If���U����*!�#Zhz����t�O�^~�q����-�5���T��I�w���t3]�!g��$�TM�#Ӛ�K��o K�T����TC���L�cH}oE]��Z{6�6#[�([t 52�������5���C-�=�������>�F��a�>�/��,>�f��<��^�U��GIO��ө_1}`���S��>��*:pt�B7<��P	%��2mf:��as�����xua�-=d1�������ڍ�p��&=d�+�~��T�� H$4������#��q�M?������!��p L����o[�/֤M�u���?5ެ�6��1��J�T�Њ�LhЊ��~��-5�y&�8̬��ۡt��Y�+�n��8�s�3XEBJb�sϽ�>����c�q�Dt��]~�%Ԡ�[u�	��F�^�s�^kX���˛�4o�*a�Q�z;�4 ��B��[�d�]�����ux0�?���Ѳ.̓Ӱ"�ˋ_�=��{�?�~����+/Og.Z����3
ȕgw�'�����*p�OA����S�F�K�L��˶ �����|�xk宴6�w�ەP�Ǝ�R��V�A @��C-���I���ٷ����l�`q�Y�nl�2'��d_�B�$ׇեw���D�k�ҥi4�0G���9h�m_���]kor�З��2�O9�Z��Ĩ���D����f�-�HL�r���Pݪӆ9���V�\�@M���C�{�>�i(K�FٚGp�<��KJ�i�����{◱^���|���)e��l�	�A��W�<
,՞�?2.��;�(�o���/����]uQ�Mtz�Mw�ݛ6����"U6UA�ڒF!RbO�H6u��p'�����'���nc(
Q�����\c�_}u����CU�0�E�<}�g����_sdI��O`�GFPd�:^P";���|�tۦ�6䜉(eM�)�-�i�ģr���r#� I��j��뷹� �M4!�(IL�e��N�#ݟ6���2��Y��93g3��r`T�[�]���ȗx��w�]�'�؄�k���q��i������*�GFZc@�0�)ag��>��3HH
�0s��������}�ڍ�FU�?�{�QG�����:j�zh��(W�}��5q�b�6mZ�CXr�h��{]¡�%�逕�8�Jq�@"��iᱳ�нG�����:-��9�H֌� ��g�{��(�ȼ�%�ֳ�(���ϥ�y��D�� y�|w�o]55�������:�X<��C�3dl3d0rhՃ�<u~	|:��������Щ���O�xJ<��d��X+ѣ�����@�*�E��燈���.cq��u����@.Z�剉h��s���J֘7�đD��ׅ"��
�3���}%�Vȕ#]��q���!!y �$�r�i�i���)I�ٱ��qP�>�B���;#�:�y GVO+Ә��=��9��r���? ��xv��Dߌ�֌�BE/���eX�yTk>CE�N���G��#꭮?���]߸g����_�'�3���_w��6�BP�	�wS*����1PfΜ9�NX��ٯ�2���%;�#���ϋ��	G���[�����)���L<�����kh��9�6�i�^Y����i��Vs��X��=W�:�(�q%%Έh�_o@��c6ʾ�����4l�h�+��z���r(���Q��̙3k�[��?���:�0;X��RC�:l��K��"�"�M�a��%S�է��U�}�H�_y)]�����4O;���s/�P��@Ic���[��h8D�����>��5��_5����}d��&���*E�E�����<����*��X�t���Re�=O�2%-y�y�Ng�%b cg��L�jAģ���c�!�3��_����P�o����gE0k�������c�~r���N\��E�m�_����%�%pP�s��O���=����G�P��$�Y��g#��:��][�t.f����>z�s�Y��y���-�F�C8��Bj(�M���L�#G�M���K���9�XW'��H���υ:X1`CIK�}((�u�`��NZ*�l.b="{k��h%y"��f��'��6e�e�lw��C����~�����=��/�v�ݻwq��d�@�|n��h8*A����}#���K��i\   IDAT/@��伏~�a��,զYtAL�2+��j]y���!/[�,��^���D��&� �C��n]_�8��sa��u�t�5����/J��r"��@,�@��D(�j����9��Eݿ�Q�Q�(�k�K$"�-���jE�e�Ip����f�����d��ظiP� �0*�����< �0��� �������a#+�`��wȌ}�O=�4e���j߳gk���o��2v���M�u��qv�����:�~�^-B4-(	Zv������y���K���+� ���7���l���ĔA�A�ʏ:���Һ8&z���@.X�0�>��q�*��Gf��b�,�~I�2����[����k<�#K��~�-x/��V������7��9`h��۔ wRb?X����#���w#�Z8��ga�J>���?@r��iӦ��mi��`�u�N�����n�Q�!6���;����,2jK�-# k�A#����6���4�������[�׾t}���KR�H�o�u�m��c�C���uۖS{ E�M�q�ɦ���7kt'���m�i[Dx��.�_z�96t�^��e�C�����o�l��f3���3\�a�<HVb��{� �T��H��Ǟz*�ɨ�~	hV��T8թ���mOf{�J��Tf��h6���� �[~�q�L�w���8(�ź*<,8�j�� Z�n����g?����`j07x&�[��}ڽ�IE��<�؎p�o��m�u9��acǣ:Z�f�p���Ph�\����Y�ݨ][��&�Ё���~9��Fjl=� ��:p�"�v��헿��;��t�嗄��_*��1�w�yL�������lh�9p�TA�ARÝ�bL�1j���	��h�6J�s�,D����1�öI�A��埡�瞵� Anæ��6��J M-y�DQ���hAF��t�}����p�VuĶA�w�M��^�Y.�"�6d`Cy;�3J�����������/b�ld��.a�|���E�F�'��#��Z��1�Z���
��o���.�Q]#s<q�v�m��K�]x%��-\�Yq!?ۓ�AZ$k���+��tR��7a�Y�sW�޵��	��9ˎI �P���sω=�κY�5��Is*���mc`�@�2���[��<��3�vSp�|F�^	�ӯ�F�1��!Ǟ�����(�V����߅�(���<Wd���{��������X$ϐYw5��xz��6X�n} P�P��gn�K$�@9��%nPV�б��lӊ?��ʋ䥸�^#W���δ�'e}����?O~LV�+����S��p�y��Q�a6g���'ȔC�(�ak���)>���s�$���~�8�-�:Jɝ�&��z�;k֌��y��?�wݡ���[�Þ�B1Y�A�l��0�A��u��h���C�bT���	������DZ�lI��'7 
2)�y����} �s'�ձI8v,�u��������0_͎�,T7� ��j��ҿG�Y~ ,�����������x�2:`=��Sg�
E�];�E�Wee��Q��UKơP�~wO��{bN�a2�eK_� �	���H�Μ9%�3�f�/C�nO,n�V�ل�cּ�52��`�!��`<�a��Q��gL�>7Sܼw[�8"]��_O/>�xZF�zK˶K�4 "�k��v�PN>�d�2:ls<��N~(%3�A�V������s��6נ�������ƛ~J]�Z�a=Xq��C�uN�{x��X�3"��>~��i��-KO=��2����$��9�A}��!�F#`RUIM�5�j���4��	w�A�5�G�:�� ��l�3X�quz��;JfDy��'�Rid+8ɲ�Τ��)c��}ɥ��Ka�1u���X	R�(�aV���o*�����/���p
¼�uM��������,q��i�}ƾ-If��n��6��d� 8t@:�ܣ$rT)���D�SCZ�bk��7�,]q�y�H�R����R��2ʧ�y�E�)ih���YDDр��N�(�-�G$b�Dm�F��qg���|+���Yk��wx�?��?�aB����I��]�b��UX�f1嘗��t���DŤ�R���P/����+&���{3��+�l�o�'�����nM�0��h$�K��IGі��Y�d4�g��i! Cmk�j������!�Y��_o����Z9L^$Ibc'2o!��u�Ӧ&{�r��j�!��y���2��������'y�|�_�}�����w�}����Jg��K�d���zȢ̒��7ם*4D8���L[Q=�R��b-�̋��fOM�����M���w�%W]��k
''��́�v��mpb�|+�-{`��9J�V+��I���?�|���z&:�����w��oE�[B��dY�fs���ҟ4IX0|'mjٹ"[Zmg����������Kp�j����Z�~`Yz��!��#�O5����a8a�����L��g�z���,y}�B,����"��vZ�g��/``:~�I��3O�𴅾r���"J��B�m��qv2r�,~)=���������f+Y���3���8-ujܡBg������.}�X�3}�z;�Ț1yg��Z�������YP�8;|�u�Yl&�bk׮Ef]�Lv2�k=}��t�1'�V��d���l�)^���g�@< ��m��N�� u�����7޷�Eo�s/=EW�L�dl���kʙ�������ףFק�({�v�Eq��q�����?�����'��	`��C�!nm4 ��z�I��5J�W�_��ٯ�p3R�ĸ����w���y+ɧ���j�x�"�q�}�@�kW+��3��8+�mb2P�;qQ������]��Ȗ}?���_q�8�a���
~�k`DCΐ$-U��N=)��^��WQB�B���l0�UMMC����q�u��D��>"����f���=>�=����A�I��5�arZ�nZ�@����o�~�#i,�&�3����⠿��(���@�ʝI^MA
�=}F���N���Q�HF�0��}�9䇧�l�H�f�ͱfN��zz�&B���7��#�+�W7�%{�b�z�,��JH-GX�6e��8��&r��YP���7��;�O����K(��Pv��-:��?�%/�/���+��������ܥ�����wp�%M�Ȕ>��=�#&ɪ�A�6 "F�8�������i��k����4����;f8����m�9fdA�����U^t?���]��0h��g֣�D���g�F�1u�җ�\�GyZ��ca$���ɢ��d��ګz�(!i����ӡf,�����4��5͘��i�V,��D-d6KPU�:�_��M���_��4$3��6A �q�+�`�h$�	˂6zg�d�b�َ9�t!�(J����=:�:ƴ��.�ܶ.�����$D�F��*pu����qnM�߻�	���Cz`��~�����_�5�8��
]�6P�Vd;�1�֘3#�l2"��_җ�����v�Ѐw��%2�}�� �9j^L�@
�� �>v~�
�����M?N��Z�XC��VF.������Z���84ӷ�V6�:p�}|�Xq0��}�aX�VA�0���ѹ`�;A�mp�!��[{.���&�a�t�Ѐ��B���$é�~�c��6F@����Uz�Ҁ��_zy1�K1��](S�5���.<��%<� N�2���ck׬]�M	ڞ
[��zΒA+3F𬬑���t���s�z�����7���5x_�<��t���e�����Y���Z��3��}Ĩ���՞A`�u�6����t.CuZp{���n'���|��7'�	���r��vR�F\��ܢd��l�Z+ �m��/";5Do���m�z˳��罼TW��ǑQ�>B\��|�Yh{@2��IS@��"S�/�&�<���"H��?�~0 sow��͋�G&����u��/�6�HS\�����'^���3�����a���|e؋ ���%6�@�(�� ��2��$��������7��2]�c��>�1�;��c�r_����w���4t�,[��7#��M�L/�b���,k(��CT��賩gφt����v�-@����	����8J��`�Jw�v[Z�tIz��ѣP2��Ħ��WmFQ�V}�F��nٺ���-�^�@kR��Ó�SL��d��J�s,l�[��^Θ�;T:�>)�|����Y5�q��F)�Pr�����;T���F�|e$n���N���˞�`���M::-:�R�)�P��
S�d���-_�23m�˅c���~�k��N���1k���{�c؉=�B�ag}�0�� AE8{�~_qPb�AN_�����B<[��A��%�;�M�ǋmr<�Ї_��_����	�O�2]���nvG��5�nF�Cn:f�<#����+��S�=�/N�9k��ϞwC��s�?FӰ�5��5>J�Z����#kXE	���\F��;f��&��3M�1=�q�	��16$ C~�՗�SO>�J�V��ס|X:���dQ����{��ؑS�N���j0�,�x)��0�Z����`���k��AN����7Pn�� �1(�O4q0IB}x��?�=8�b{Y.;'r;���[���&�2�J[AQ�;n���8�u���X�0��Ґ^~q����<Ѷ7`�9~^�D�<k"
��i�	��;¬_�lPR�����AĶ4f�΀�I�;(���n\�����~����u˃'o�REf~�7����V�����`����  �^{wu0nv:�,l�8�$�8Ϟ�L�+�L������X�BG|_����ap���Q3�@k�^5г�McC3z	�kp+�)�$�I�@�:�rⱏD��	cof�ߐ��{QgYܗ/�3����W��/޷�ﻟ��� ��h��|�;�L�SҲ�j.��Fn>���=�U���	�b�R2�?Y;����Q�W͝;�:���_�Cߺu��>�E�ٿ�����
d������'�8�WVmN/<x[��O}��ɶ��.��ed+^]��?�X��ɂ*����A��52��9Nֹ1e����&�7��X�0�`Nv`�Z��J��F�Ț�l�
l]$|�ak�q�J�V!�����$�P~�尚��u��C»���}�"�﹅��:���l��X�$3�E2��?ݐ��1O�>/�v�-�]�Yg8��<�{�i۽CqfB�*�p��V8Đ��YHZ�a�+ɠji�YG�?���޽+˘��!*��� �c*gh[�St�Uf1����huop0IWd�C�$��drU8HY��a?v�8���-w��k��=-y啸�̿ރֿ"�fHC��l
u|~/�pe�/�sŕ�Հ����M���<}-�ߋ҈OE�y��?$��6fO��	�+iKXWռ��4`�;X���Ʀih�W�(Cd�����M/�)M�A(�ɦW�X�3o��`p�p���ʚN"f�4��#{ShF�Dp9�dى=���A�=�i)�}x�f�_�җQ�#�&�ͳ4������<������Ι=3�Z����2=����~t��6~����:�{��XcQ����.z�E�C��T��U50X�A�0 �5����{�v6�mf�������:��_�O	�EՐ0&��?&r��N/��6��1c����W���`����}��F�遇�+b�p|���e�BlȽ������ʘ�f �3�p�왌����Ϭ�.ڇ���e���#���G�J�E %ҡ��̼tf�����n�_�gv�V����<v����A�����E:���~���|���I���bO�.�lQmYr�	���dU���>©�T����`��S���D�{���q��]=}�u�w��|��CG�w�#�<��ߜG0fZ�Gs:s����:�w3��O���ۿ���E"{8!8����T�a��ʋSe�ؼ��R^����{�L�r���+���ּ=�i���鮽k�����7���'vv0b�,�=h7����|�5lf�������������;�<P��Y���pD��iYh�)��;6�Ζ������+zh)bǷblj��~�<}�Uג9�'#7%��/b]d�Z�UE56��l:2Sҵn�x�ö�QY�a��{nNO<�@j��(�*�\�$E: ��ui�����ԀS���Y�lYz��;S;pZW�}N��s7�~>�6":j���'��k���܎5�IqXc�dq;��� �_p�����m}���Ű*Ho��h?����Ct�>p5��#mz:���M�& �?��}��� ���bt���D`u_5�__��� �kv?���!1�}����尚�X,!�6��V�Z[y-��#2dn0���cƅR�*k�N��f�Ou�m�*l��)W;r�F���Q���{a���!���Ll�C�d赗�J�,�AG=�����\����f����w�N��}Wz��!�*�o�Pj�H��2��y�g�s&R�#!�eE�(T�U��I�118޽kAP=���k��ČIy\_��|�>��C�h�� I��U�9���ﲥy�#�A؜�9~Jڴz_�؇>���k5?��e�י��~�#�w�c�� �K1~�$��F�����8��!G=E�����o2c��2�+O��˘{������h�ž�8U�����܎3��PA�ht����'�Rc����������N�r{�%V���N�����i�I��ۦV8��?L�e��r{Y�jϼ��+J�^(��)���3��I�[��������I�ȳ��n��Ck�ڹ3<g��$LΈ6�7��7�����ɬ��,6g�c�o��s3�Ul��!$x8y0��+h�=��t�M?J�'�J_x~htW�v3��L��Fz����"�Y�(Ǎ5vFVV]	�Y�6a��_���>z��<�GG��������^�!\!Q*>Hˆ�����ҝwmO[�?A��0�Jb�q��qpCц?炋R3��%i����m�.��b��x\�,�i	��	�D��MM~�ȁ鴹��Bo'�h'QܿG�������_�r���`&���˫'��1��&ON�׭������K�ָ��@adt�]O;u���Q�����d%�e�����@8-��
�X� _�4F����$���ZS:�3��&k&�}������ۀ��;�\��5(?�G�γиΘ1'����xY���eh0���:�(Iv���r+ffP�Qی 5�빿�4�c��Ǟ�І�q-����o���:�T��U�1�����q�	)�Y����a�ҥ�]�k�u#a�s�4�FC�8]�4�5�7a@�+]��+9�̙u�p��|4�#2�χoD��C��(1�Q��z�
p�k��Z���Rd/z��\�z ?z+%����h7�ՖV3>�I�wH�s��̐�q������N$p8�U��!�4ԀCS��w��h�����ٯ��)�.��z:�9��I�g·+�J�}_8U%e�x%6��l���>���LrX��)e�oVo�!%q�����3�G�=-�8"\1�|,봇@oM:�Sr0 ���J��%D����K��@dJ�s���ǻ�7@�o�|��~n'Z���}���{�ޛcQ]��~���#1�/������l��|
k�3N��TE�?�ē��?~e�y��{�����{��xh�Ǵ��O����xv>�U*0&5@�,2��!��?�����_��V��e��|�|��i��5�3N�{M@�@Xf6j��Ua��]�R��i�ů�L-��4�Q����r����6ȶ����;��I]�:�D�ud���2oO>>ņ��Ć/E�E$d��HX._�x@&�I��綥lX�Z�B=p@�~��}:�{���	fx���ܡc#�?H TE�:j��0E-�q�d��� �����m�` E�(S��wݐ���"�J��@F���v�����ʗ�nV̅{�D7��>���h6;��'��|����7�����JCn;[F��h�^vi���	�ˎ�}��ꐵ��J��<q�Ϣ�TM��n�.�P�ǔ���K_q�%���*�c{��"�ֶ����?��� �%�����!��bŪ�-�X�j]@�ĩG(eڌ�\��N��ƥ���P�x2tX�jQG����RFX�:8\��4���D�$9��P������G&>�Q��M���(Z�&�oy}#�^��@N-��Yf1��������t�</���g`���4�n�㏛�>���\��Zg&L�XK!�L>��N ��<���,��n��Ï<�f�!z�e��Ub�4N��*�>��O�q�m����z�N�|�����v Q�a��Ls���\v�N�<�:-��)��Iu���N�v���t%��1��s5�\^9�Bc�\��d���D #�}N�����^�##!� �<fB�ꓻ�G0\�u~<ߓ�M	(:��x!�hv0}��y������ݹ;坦��w��n,D�������̅�F����op���������#5��/�������*C/�:EP@�j�����2��_���7��=��]0�?/�M|d��PAD)��"��5=�w�Y���#k�	���X�F�ΐ�6��g6��+Of�8"���Y]�(���w��A�99���h�z��Y�����R�0�i:pP�#��'݈`�a3��-d�;h9@C��Y�ԦV��e��,jjE��+���မU��$z����Y���d�fM��m�phJ8~%^3�ށ�=�Ƈi;E�yq�᷾���d�B�Ρ��~��t�u┙�!�B�zhB��Jo|����s���/��%׈,�;dA�}���fR��lU@�u���2�����`��2er��TI�N�x��p7BaV��V�5k��q�zBO�pum<��uӡ��˾���/D���930"��"Z��3~��-���6�L��I��B��FUrY#0�\��[q�2��
�gB�+����69�v�	d�C�#�h�M��8��jbp�GA��CMT�k��� ����eO� J �8�9X�n%�Z�����p�J<7�_<cIE�c�� ���t�9�$cn,A��+R���?�0�{ҋ���c*n�q)�S�t�Yg@&�4�~����Je��J� ĘSQ��>��W����o0����F�`{( �45��ڄ�G�nJ�{zz��GS�sg��.�<%�����k�yN�|'����Ta��Uk� �j+����.���{�Dr�$��@��#Ҿ\O���R ]����_��1��*�\q����W���Wr��I3Pk��'�uυ�"'Q/�Au�^	�d��n���l�����(m��L�S���C��P!�%}�ۧ"�	�]��Y-�7ɨ�/-�8�rE��wF [
�J-j���k���8}_���&N�����~� pOEs��p�?����={��̡c��]G�P'��
��~�����c�#؜�@���b*�%����O#d$�Q~�$&Fof���L��݃�2S��&7~���ۿ���λoM�ů��?	��i#$��6j�����5���cǍ)��[��ng�֐�	��D,`��P�[(�ƽ��ѻ�+�����g/���x_�YH��}���P�D�;���IQ��^���u��}��u�w� �:��� ��0�+^y6�����w~��0�8���J`N}r��G�ab�J�~����ϳhFa� ��)t �� Rq�5�����2\-�3��-z��fN��m�������q�ƍ�W��w���D͵j��v d������"�r��%ƾk���v�T�5�-&�	��PD&�˗�F_�H e��C��mO�y��W5�Ȇ�O%�F�8vB:��(=�Ꭶq��P���Жf�"3�>�%z�,~M�V$-�ĵ���E�q��$�jt�A��`�|�1�(��0���TP��a?����h�²K:Ak�ٷ-�ꑥ�l��)4kص�^�J��i	�<^cf�bf�2�ǏǼ��	�hQ�j����B�ܮ^�J��K"\nMw0���8�=#-�8f6#Cw�$Y���B���˃8�u]Ap:<�;z
��umӼ�R:z�	�~�#� �>kNz�G�K���[�n �0n�А��1u&��S���ӓQj�Z򓲷�ӮDA��y�����;:DS-)��ܓE�����q&��X՜�vK���iqm#G���-����ܣ�EPs�?�=R���l��C��������㿋V���x��w��������NT���~^�>��ާ��p�}�������AU�V�w"��k��jk���P�'�x��im�o��{�Щ��ʵZ��|x"��U,�8ϐ$��#s7~�F:lDڼl�&;~7Cey>���`.SC��-3��^�P �̱���S���]���	�g?�)-~���.��d_��&�-�!�Ԥ	���0�R˞-�l��$K6 ��q*m"����\���
E����H�G������-b�#j�?	b[������`�*�]�o�q�Ȍ�𑁊� |B�b}3�}V0�����+�>C�:��I�Wn"�Iv��>xp#�Io3��l��n��8Tڣ0�g�y��c0�f�<8"W�Й�vC���Mh\�נgE�'�X���,d޷�ygz2���ρ ���C�J����0�|_�����ӯ|���߶.�ʔ���9�Ig�Ӗ���;�� "��c�����K0���y�c!ɕb���_^k-ڞ�Z�4=�#3���'���w�������n�)Y,~�(�Ӳ�6��ٯ��<�R�L�\�Az��R�p��:�� "�������.8Le@�m��S�Xc&���I��9&L�#�������8��D:M�t���=���c���FrL�������8O��#��{�JϿ�J��ruʼv �nܖk��&-<�X�f�q@�輟~��hj�V�\�C�C$sN:��8lH-3���t1q�/��Ngt(���	r���~zg�{v���(�ت�hX�b�%"e1��
�`�6��o�@��3����m�ړ��k3��y�k�tj{
��@0J�z\����A��c��N�#�2Y��Q,� 3��_~�qt;��b����<6��c�OCd'l#�,�t(FB�+j�w��>k���oU��=���<�Y�T��^�9��_.���v���RnGq���wоW!�]Ŵ4�7�E~��ۯf��w߽��PSL��ϧ�|����TM$��Ӧ�-�۾�~�s��@
Ñ@ĂÜ����O�_v*�u'!�r{���W�[q��t��fe�J?�`z��G�A����Exe�n�ۆ�iu93�xנ��^�hq۲m#��1ٙd�*HaY+Y�e��Or^i���Ӭ֩h�����{_�~���s�#�	  ��;Ƕ.;�y�II<����_�*��2L�RɒtY3�7<G�~��Y���4N�Z3G!�G�Yap�u�[�,���gf*S<�P��w2�-�>$��/��=ޡ�mK�ſw!�c��
]b��
�҆�j����o'�K[�����K�#3E�n����v7k\وX́����@j�c�Ng�N��A���w���;�Z�*����*�"֡�h��WMvR���S����LTs.��S�X��s��Z�{	L���M+�� 퀃	e�H�M�]w�q5q2�[����RJ����)ą�v�݉����7H��󣚿����17�������:���������x��Х3g�!t�΃��{3k���e��.$f����A|����7�� ��W�s�ly�87�1�U־�S�oV�@["G�3�z�f���v9U��n��y�2�a�禣�bA���: f>�־.��_��?��B_�WX�*����[r������}N��J�:�l����女r���|�6&J;�1��|.Kԝ@��ki�E�ɘ1cA����_?�E�u��DSJ*6�]�ƨ�M�ຯ�)S��Htpma?|��d����G��N���JkԿ�ߊ�w�Ũ��u�ޟ���P?�]�>o �<���Y�� β�L�8�G5��_�Y���w��7߼��T�Dr$��p�E�(�d�g!<�|��;/I��V+fHz�X5Atj!�m�"������gշl��w�ٚ�`�:��T�:9;��뿗�{���K��E~��v(6`{�.j�����;9:T�v�ⴝ���ٰ�J81>�?F��f� {�lP��ҡ�Y�����(6x��̻(eQ�����B͎�P���:q3�!��m�5�V<�x�g�m��y��w
)�IM�� ���U�����`|+�� �%~~�vb\�JP�1j���+o*4���C�G��nW���L�Z=��9հ� =�q�
�ه�f���l��7����{ax7p�zu3�ܓ���7����`]CZ�go�Vf�"k����a�(�4�U�rՊڜ(�"C2�Ն�T)N�`�#�5�j%�J�w��N`p�eIw�QZ�.V6�Y�H��f��Qw��
l���L���8(ÚY#'c�OC��zz�g�`2K�w�y0�eR�O�Q�}A�4�A�md}�'��/:rJz�̣�{��G��A֧p �/��
%��~����1����;�U�{Kr�9��N-��\��g7�;��s�d�Y�e6э�ۿ����~� �4c�p8/8/U츌�J��z�锾���ߚR�`�g���g*j&S�3�""��8_�L�#����{��m���f_�'�H�^T�7/j�Ey���-�xN�u5�P{~U&�e�]�օ����?6�)r/E)i�ĉ�N��r�$KM�ڕ(�hZ�Sv����>���W� �������E$�2շ\�_�~^����¦��W��ޗ��]�����{dD���Ϛ=��S�L��ſ��̡����/�1甯oyM9��p�ƾ��8�N�PϝL�V�v��Ե�j��T�	Qn��i���ƻ�ΑZnɱ����ܖe�e]�Z��I��N��_����/�/����矚.�o�4AbVo�X���	���� M�n��@1�J�56��^r���6�����̰��ov�]�^�^��{7xdq��00}�A�sƜ�i2��첐b$��qt�Ԍ=4:��q?���ŵ�����5fu*�E�n����X�z@�\�A�j����-Զn���ܳO��A`B����m���Ap{����S=�>��#�O
g�}c���gϙ	!qs��U�#+��Z.��%/BB�$7k�G5��ԧ3:���3{��Е&��/�	e��2��=Z��8���/����^�"^{��P��Ե͛� ��ư��(~f�q��]�ek����w 6�vdYcQX�A|v5��n#$����qf���@��H�K���{	s��G��X��N��ڷMP��oSCI�?�������kՊ��O<D�C8ى��7��,��3�&c��pn,[��'߳�M�����/��<��p�!�eD���+W�g��WDd�4�,i�M�����ڒv���ڵ��ݰ�;��a�L�J�8��KP+�������k߾i7
�ݔ��0aq��"���h��b8�g*�9S+��rp�!�7���`q�|}�{	E,�W�K�RBQr�0�~��ܻj< �t��ӓ?y�4�uuz����f؉2&z�����f ���Ȑ�I@�Ya����~�	�sDv2O�́��2���_�{'�O�����*iU;#~m����b������������=��g�y�wP�+7E1�$W��W&2a���=��x�FÃ��XՔ���/���\��M����j�=d���?�ij�;����`p�����.N�^ô9c�4���/e�A��0*�Q������O�[?|x���Q���FI��ň�8����fm@����n�)�w��d)N�4׃���G�-���כZ��G��3K�(��/:���7�!� �^XH^�vEz�GRce��vW�}�g���^ �=��0.�M^-o����e$�%�أ���0�-7]�����:��e�8��p�>��Ҷ�k1����:b]k���cZ�R���k�������{Ȳ2���Yy�aS��h�zR�@�k�H�vvC�jN��ԇҤ��.�-�$Yz���R�ߣ��d������6ͱ�5u��8]l���8�)t�H�?�dZE=�_�Ul�~�Z�?���c��߫�m������n��g0�CNi������!���m�RL��`d<İ�b"��=��\H|�L �L�$� ��������!�Qd
N�<�dz�v�!#j����8Gg#X��_��:�g��_K�mJ�3���R��{�K�<��U���C����9��r����rگ��g���a%��^�kA�-����!w�pc����J��ҥV>��P?�P��� L����r�`��%���������G����x�9�o�v~s�^�e��,�}��n�e0Ɂ�������fі�2L��82��\ߺub�6x*��ئ�Ii>���NX���?[y`;"8��ۛ��I(��3�˄�� @���_�x�6��%�� �<�᭿2*���څC���N�Ϝv���{�7����ԡ��h͚5����-���������2���Jd�,�Qߔ捭OOX�cibh�/��\��Q2��X�q�9��������at�8��B��!��]��	��0�N�2k��aؘ^xz	Y��0�祓O9��;�&,{�,T�&9����]�8(� :ؾ�rᒳ�uM=��͚�H�P�Q5�8 嵮��5~I~A);%���4j��C�u�q��ui'��A�ڜ2�l--yh�F��
bf��3X{�G�B�ݳ���ִz����d玝0�zFtw@�At,ݏ��f������n�C��<H�?�'�2��J%�h?�R�G�}�E8g �cdTa�dqw����o p��B��i#��}�P5~:�
����)���R� �nk����c<���䳺���cmJ�dɗfP9�IL�#�V��އ3VGp�7ۄ"KR_f�w�!����Ǜs;��>�ؓO>�����O��R�9�9�3>�vێ2�g �FONU�b=%��C�5d����S���L}�(I8%34�J���}:-~�Y�h�5�d�l*����N�p]0w'�W7mܓ�y�G`��g���N�NP��~�18c �Ef��L+ZɚzM*�����O~,�z��A0(�Cs|�m�V\�7���DIr�b��t����.�"�p>fϝD�ZL��v��k��Ae���>˵4�\�qLX�ȲKxa����������X�c,g�+SN�(ō%2�$�)J��͜=�d4m��@Z�����L��,�a�\�9�ڲC?H� ��D�����-��)cM�>�7!
T��I@�����zo��Y���BH���rN9�Xا��}]v5�k鿋����r3���
�ޝ%�RP#�}gcCçN:����}��~�=u��ׯ��d��
G�Gk��H��_7\���Y��~����Ծc}:���1d�����7?l����_O/��R��^s��m�����$��~W<c[�d`�����9g��ƍ�\)ӁB���'؝�E�F�Ya>[�d�6�4��(�fv��$;vn��nfq�T�.�5�E9 G���(�Py�P�#ziC���F=C�9�عe���)�"[�c��4�� �p���B�`[�m@�w�?�����FpGDCBNYs'�8ߏ1�~O����?�*�m��������qS�fM�3FHš.8<���/΀?y&!5�%=����0a�;�;V�C.j0�}3b9FN
�H�R�� ˰�s_���4mꌜ��v�m{���{M�ԛeU��/��lܲ3}��G�j��q�:��֮��<jv��d�
Jq�q��u�&�P��w#��u��_x�9JB�lB`9�o	a������Qgj`���Ҷ��k����*�s��.�ڐ!W�5"8���A�Hy�:���t2"�
�y
p**��=�#'q2�T��<��3̎
4g�Χ�	b=U��3sF���K)Q`���"��n���z���cp+=�	�[ �fq��,��6P��ؙ�ff��n�=��桃�t�[��JХ���
��������c�}��V�0NR�3q�w�Ź*iy����C/�@A����OTL�ˀ8`r�Z-�l
ʈu��]��Ă�W)�ϊ�z��Z>��#;s���؍������ދ%��n�	������;>�8P�s_��aK���}�Ϡ�	2?b-�ާ��͢(�r�]N�+���:�;����(�ꏠ0���r!{�g�|����̟?a�������NxF�VC��r�!e�3L7�P�z����K&ր�Ĭt۫�9��<�i3z"f���ҫ:=${��Ј����h&o�`�C���\��p�s�y���_�?���A����T������1R����,]q�%(���Z��ٶ�H�h��'L��B?�"$� |���@�/l��ES~ �|���v������C,��=�7�f��=)`�i%�P{&oٻ.��v�`ζ�Ԓ�}�����C)p��m�6�:��:�U��?��!��o��t�p`�y�1cQ��c7Fh f�08'Dk�}gm��P3�k�
A�` �p�W�m&|�k�%�>�Wg+K����T�:ز'\<d�����|�~��R�����G�8�����\q��i�i'G}R2�~X%�f�q?������y�q�a�"?
���`˟��$��E��Ԍ?�x����6�[��
͐u�T���u���	�^Aհ�=YޢA�K���?j���ګ�#��L�qԲ�5�w��j!Zۖ]_�㭶��q���A&�R%��2uu:�UH���n����<_t2r�'D��L�"���7�F~D����D7KrG|.U�<�<�@(����$����-���K���)Q�W�{4�3����-ѵ���EnJ��H�p���J{�q�;��K��4�iT8��y���9��q�:�2~��^����"hN��P)�p��o�"�7�^>bD�8yR8��:y�T�t��Y��:@d�!���� ��4A	��������3l��������[o)�<�D�j�s�E!.��ُ����z���:�*G�ۯ�������8~�k,�zy)�s���I'~`��[�������4CwAo��5���}�E�^l ��=�N��tx ��Ãӓ��.���jGb��Da�1-8� �U�C|�V����MS��>$���H�Z��#� �ƫ����������o��}�R���1ԕT�I��N&I�膯���c8�ƴ�Z{+3��8�2Ł7����2��6�N2�v�<U��J�v�N=���{S�Iw�����q0((�[Pﴧ�\���5zY˃_��y�Q�̐pNf\?a�Ì��=uؐj	@��䭢��9m%�P:�Vh| ��&��/�,j:�$:(�fv�]�ނ�:�dh�_�����܃��k�!�Dv��ēCEn ٩H�mOA`���r�R8V���|a� tD�/)�T�e���@;�lQ�\N~U�Vǝ[#kj��/�(���r�Gcm��@&��s������疘ϼwof��˅C7(9�c�4ql���̀"�e�lu�0�A̲3!_��L�����>��֤��U���2�����|�@����~�T�u*10�v<z�������Ŭ;Ϫ����f���o�w�!o��5�h�I���2�XֆZ-N$h83����� \{���W��P����u�b��nK�F40[�)$�-z����nZ?��nM��g8c� 8R@J_1�u~iɋ��:��h
~�h�!�Y%ښ�d�bj�ݕ���c����Ҷ��D�+�y/_���y&Bԋ�=��:��}\j	4=��.#}A��UD1�,{�a?"�u�i[<c1U��F��Ҽ*�'�5��TAxt?�\��������p��b ��?��y睗ϔ�-��#����|���y��%� �1)
04������h�Ǟ�K�Cͥ�#zy]���I�;���wp�Y�����{���8m��ON�<��m�_���ݵ����v��at�du%��8FP�-��H��q _������ө瞑����6�3{.FE�i�J�M���55��?��KV��s�A�f���F�K�or%�p�&���8�r�)��������SN�>g��b&�.� =p�c��K�H�1X�Vm��r��*miIɐ��L�����0:;���P��+���l+1Αu�Yf��9��%��)�c���Nq�s?[8�0�.��9 �[�tJ��?�P�H�������kݛF�1�z��c+�ي�W����R��R�<�A��-�����s(��,p`܆������]�v`�w�x�)WdV#�:g���N��ύ�N܌Ӫ$C�&�4��dv�@���P
��D�@�i�=K`�z��iS�P^�K�����h:��b)^#��$~�OneX�z�jK�=w�K]t-�w۝�K��	&�sTq���7<��ә�w�Q�k�X1'�[k��8j�*WiAD'�$�'�"�8��������}��v�D�#�T4����!c"M�Б)3Ǧo]��t�bOı��N���?�L���i���+��m�t��Ʉ��o>cƼ4u6�	��}�Vmi܍�`j����v9�d¼�̬3�4&F�\�-��}���~6��r@�A6���03��汔�^O��,}�cg���@�c`��|�M���-k��-5�W���g�D5c" ��ҩ'�Β�ǈ *�*QF�t�$��p�N0��'�,{��|�Y��/y������e�nz�=�� �����vw�	��G焁o\C�� I�`���B�����M�[~�����kp0�M׼�#�'&r��3	(�y�������3���#���a� G-S��8,�-eo�ɵ����8�*�l aj������3�S��d�VC����@q�����t�{�����#.s����oE�+��ޯ"Ȋ2�3�*��y��o�������s��}�q��Pj���e����hR%[�駟O�7H���W~4����Ӫe����>7n�f�aC��YG�)9�'���oJ�y&�Xѐ���f7���H��Uw�8unjM��/O��|���c���3��Fr�����}�b�/<%=�hǭ��>��RUC#��[1�c�6X����,�!�iĹ�Ș҃���J{�J��}�"
.��>RHbK��J�y����*e���37�����cv��3_�x�}a�z�t��A��gPN��D��
� �QM �!v�1eZV�D��!/��"o9qҤ $���6.[PJ$����� }���ӏ��T�Q���\z%`UN�����	:�T��F(�k��h�fٲ;�Pj�a�KY���� 2^��׫�=tXS��u�w��3PT;���Y�^_��sW�S� V�4ir�;k%��� 9��6����d<G`�}2�J���0�-W{��k�c$f��9�]�jmr��(ښ��S^Avz޴
�7�ŀHMD�X�%�2sRzq�iἓ"P1��L����+���^}� �5�thl�0ܒǌ�Dy�	8�L�r�w����R
�7`��F�a��9�NɁ�T	��4/��蓔7�uV8���
2�	pvD�6~2�j{ �zƟC�t�0u0��ß+�x_Z�����$�H��kg�7�y����(�\7�l�;=o�4ʳ��{�~I���<_�g�V��g`j��4~W��)tB�x�5�g�^�m�>u����m脽�,'H����#������O<�TZ��O~�SX��Cp*B�z,��X�R�]B%"{ř�� �P�q��H��`\��
�e�sE�
"E��iPW*�͗u+Tؤr��X˼�}�Ĉ8ʼsx�,��{ qVK���"�QL����]���^�诏xh���=w�8�W��e�b[Ii�ѡ�����e�l@�*X�<�Hڷuc���F��g>������߿5�v���l[��@�&�);x ���@���xF��z̈}��`�(��A��
U8���&��~����O��!GqMj��ux��À�]���ēO�&6�����	��E���8s�6�w����6|4�Zf]ڵe/�a;�T����d�8�խ�y�#͓�失�/_�Q_�pǴ0�9����Z���^�*r��)��ڛ�e�o��c���JՇv��7��=���1:�Q]i�Au�X�93'�Ys�q�<%�2u�?�X���A���I
���h[�W�P0�[@QF�y���H����)�w�4.�p#�aZo_�����8]|��ҴYSB�Eh�z�*�s���V<�ɲ=�8�̖7����*��[O��0a¸��r֑�g�rPO��5e|��:���v�B��~v �X��NO"Ө��ӝwܛ����[2�N�CX)����w~緂pgPcajس�D'ރ����^�М;��.�$��$S�L';ta {(�u��n0fAP6�I^��Y��	���g�d��)h�":eos}��?lش!}�o���)���@��u�lf�op�E��2��;o���l��<����$����Uв_���	4L	TC� #�U�(2�3E�rDʜG��3���0��)�/�^)hU�B��2�vɔA��v�	���GN}�GUֶ�j��Y'ٍa2�\���IbTc�z&��R�D|�q������!@�=��w��wG�'>��QĎ4�'=��	��|Kg�8���mɅp=jD+��rhW�ݽ� ]{70���Y�Q9����J�M͛;q��o��g�a�K�F_�=۲����XɩG��~�
5�q>>y�	'�����~í�����vq�	�k�M�!��1z3HOj]���������?H�"Sz�y�� �|���&�IW\zn�3���o]�;����v�jT����G����A
'PD��C�|f3�'_�KԬBَ0�QU���$�^�}�0���u�����vG���~���K9�Җ�����^Hm����#1���M��0�7#>���5c])4�����/-��t1�p�Ev�V��~8"I>�Ni[h���� �鳧�-�I}���i�i��&Ѕ-�d�����*�>�ܓa��J��ٺe8n��\Im]��:���EO ƙ
��$��;�?'C�����Ư�a8[��'��Y���� 4���~05�I8Ro 2�q3��������MU	����3� G1Y�w��������j�r��@�l�w��@�K7�4[����;� �
�D5����_��Ɇ���G-W���F������?�?���	ջܾ��j�п�럦{`WtK�Y�����#����(�B�^v����=	a�
*�����$�5�b�l�Е���<������"Pd^��&���M�2�g��q�Ζ�����>����*�I�i����l��y�q�/J�?x'��N�ZZ���U�	 '�#�K^ie�}+i�5mV�:��s�n+k;k����i[��O���:Υ{I�M��//A�N��'�
Kܓ�;�2t3߂���K�D�qĤ���j����n��ṯs��3����<��g�Ű2�08l��QK�	�k�_+�z?I3����f�]'к�
�brM��h��G3̞�o�cՒĺ?9��쿃�^��ܘvt�I���;�_T�v�?��bJE�cC�Zbc)i(G��,>�ܙ�g�9�Ιy��}�'	�p�9Y)�+���27[o;ضx��Q�.�7��u�G��{��i�W���^�V���7oև�����c<�_���e$���ͯ=M���t��K_��ϥ۩w~��M�}b�3�S�Pj��i����m�i�`ƣ2�q#=�3f̉�z[|�9�2��f��c�Y�}1��\b����o���e5M;v�
�3۩l���}Wa�֤[o���hY̹Ț�
�; ���}7Y�Z��FT1f��7����:��m	 �V0ʋ:U_�iQ�
skU�n�b�~U��ȸ8|�1F��]z8�"���Udw��kH��>?m^�+mY�2�H�>�)�T�c��Pf7۞���u�,�}��h�ٷ�@�4-���_�&��� ���{��8�t�Y����L|{}5���pLl�3έ۞��q�f8H������2�cK:�F��<za�w�ӕ�.HG��I�>�PZ��YB����Od��ٴ'�r�I����*��)v�P�j�|"S���F���Ľ��4��Tɭ�^y�p4����w?�^[�&�u����Uaj����e�y�=�:�}��K.�c9G�"�y���ٮ1����~�N��!�R�٘v�H�����y��g`QG��-�-	�t}���;�SE9u����yqKҖ}n����|.M��lEF�Q�����Ug�.>8�~�1i��e8��4g�1�)3��}瀒�㌞|�1��dV�iu������F��k�]m�Q��vb D1	&�S���l�층=cA��?��5#�Lf��ʜ�E�܄7��=����=��V��ʵ!gJ�|i�jX�	���D�w+];�)������!Z ����<����+�y
wf�5�S^�ڵ��t{�����L!{A�H4\Kt�K���]B�{vx��������üI�!ėZW�݇6����P�LUM0��s??�LD{��E[`���ڕ�a����p3�Gy@��jY�F���~��|�d�=K�Y=<ak�̚� Ŀ~�[��ܡi��v�m�9�*y�E�-j�X��y��HF���� ɬws a�Z��,����D���«3�}wܖ^Y�6�w�Y�R��s}�ijCGF�{͚MD�C�Dne��I�G_����`����~$}��?Js'6CB��W*˩ѓ%~����[9�U+V����i�dv���/�Fz�{����t͕���7���0X��w����3��A Sac��~���)>#څJ�>3W��)����W�"c/~��ʵ�C�a)k{3���F'����3kF}:j���H����q0�T�"2/9�6ږ��/���v�)G�'èN�a`?�ċ��L�fMM�}�k�ƀJ���Fv���\J��ګ��H�Ð��H��Aj�w��)8��t�a�@�= w� ��%���5��t�����@�v�h;��Nn���;ւ)�I������ч'�XAmyD��	�aι�y�ܹ�Q�QY��-U�r-/�D H��!G�zo�������5��/���^-rT�0܃�J��Zr>�up.��O�$P��h-;�^�&M�8��Ą\O�h�"h�eH��c�L� ��0�+^�9�f��1b=�ƙ� )�we�d��\�:�b�9 p���m)�D'q�`G�gS�}����N5�3�b:�l8O<�LZ��� ��ݝ��kƤ�O<B�q�_u ����uP��bPJi�ȏ�+�np/J�[��z焠��KYfQ�(�`�۔��V@�A6���|F.Da��Ǐ� �r,�W��{�pv �Y�҆�|�fFm�jh�U���]W���U��fG<�<�u�0�<c�LP.l�P��L�E�`��������d �ʣ�M���tpM�ֳ&��A'Ic�5"Ii��0IR~Rs	0�}������_	���-�O��`�,�~;o��Tr�֞�?�>c�'�L�D!�_��l�s��EG�cCN,T�7���y��u��Ƚ�O�?��m��cf�H���6��rg���rZ�.L��g���N����-?=�?z!��ڴc5f��`I��<��;::,[�4����e��L�w�>69����0�ҢVIM*�8^w��_x�1��(�@_K�OZh!:�y�ndK��L~z㏀憤�q�;v��0��FƴM�&d7P�3�fV^t�N'�a��	#�hm�N��zԑ��ܱ��Nʡ3�b�a�H�##sL��<X!4������)%��d��u%Z������4e��4������m���b<f���<fv�ao��������s��&�̜���9N�6	��O!���z#0�z�
1e�A洣�_WEMe�����Q31��00- �[�R2R3�
���= �M��̔6��A�m�2:��W�-ol������}ۑ F�Sjy�@N��|;d�}�
2���x��;3�1�{
׽�7Xr��x�>G!�)����-}*��r桱~��:�+�SQ�xD�zFX�NX�; I�Hv�_�nM&���À��/�;z� lAN��:�=鳚�@��>�� ��D]���{>��>x}	=B)�t�fե�0�Pu��[����'��>�䒋#�l=��ez�̦�>\J#�-{�x���}�rd<��=zld�q�Js�^��>x����=�Ί�N�p</�r�/�&��E���a֦N���E�f̘���x�{;7u��3 8A\��(^�knyo�E]��;��lJ���g��	�T�c����oEn{���Gq}2ۙkPLZ+2�R�S�A�4�1b7��io�f���Ӭ/��A�#k �,�����?GNy$�p�2�x�9Z�[�7�[y�(!���5��zFF�W�3�6�Y��ߝw��_x����v��r�)_�7 �lR�W�d�9 �`2w��uک�v_��ΆSā:�Qi� ��li�6��ի���^�N?��t����~|3ʠ4o�4�_S8��8�Y3�1��)nM�شiKڴ�zpo�w�lj܇�^d]s�U��� �t���v �-�j9�+¶>fD��o�n�15����&0��4����M�pq�d:o޶�ˮpV`x;�A��h�A����B8$�/��@��O�x�\����MοX��?lV�fg��f���af���?�e�SA�Wk���=�g���H��L��?��ݑ����xa�ԧJ���pd�o�)oI'�<7-{UҚN8a[����,�q�F���9.}���K'�|L����S���q0M?6]J��bh����5�~�8�P�v���L����:d��ϛ��,-���B���7����h�G���o"+o��v�ܞ=���W��1�' A�]r��u	�5��Ӯ���`�M�������˴�#�gFZ���_fՇ�Eas�p�����3�s/߇�p��Ӽ�Ho�ճ/=��������mSj*�NK�`���=i��O���7����68+ w�
��̇��IO�Pi�%5�}����d���u[!��D��E��dt+��L4p8��h4�����ڂ�/ZQC�BQ��*V��J�x���0ý��p�rbZ�����]��b�����H�9��������~��sP��R�ϿbT����U�''���ET#\F�	'j��DR5�KL��G����=���t?h3h]��v�K[��o��ۙ>�������&;W���g�HW��}�g�#9p"GB�}�}�Ͼre���]7�}���	��j���m0����R������*��B����|��$�X�7C���.�S��0���:�m��H4%�	�*BJ��_�y�����Yd�8��ekFϓ�3��#5���!�y�	E7��a�
�C���o��M�Ƴ�90��Ӓn��f�{k���\�>�a��[�7���t�yg�9GS�v��H�D�F�4��azSz����E��f���|�UF{�����V��-�C���	dd9����v�nO#j���]@��Kz5�%�'u�Ѣ�����~tCz�ť��^A�� �i-m���JC	`���U�\�Ԡ�-I�%s9X���J�5.�3��,�Yg);�a6R��Tc(�c�uF���rX�R6�R��]�y�<�l��������i7��! N1�	���5\�!`����ӤTW5��]�M�����4吺it0���ԉǝ����q<� ��J?�k�8����	䯄�Yy.j�ة�L��
8�� b>
��ӫ�:��y�z�d)d窪݃�@�٧L����(;(dN�x�}�|<}�CWk��&��7������'� ���KA~
}|�;���#�A8��$L�d΀�W��G��$5�zX[���8�6ꥇ鍖�`�L��N�x+B>5��dq�CE5"GNc3�Į	 �>��)��oM�,��`H�p��s �M'���g��fG��o�/�"^�.��7�䴀v9��ZT�7��ur\D�f%��]����OdBQ(��U�3kvW�����9}s��5��B����S�c{��GQ����F�^:v+�V͜����b����30(��ו������2��UFǄ���7��l,
]?���-��d���L��}~���z=<�z���Q�{�On�9͙{��ώ{R��g����5#��<2��l�B]2h©e���깷�1�j�gaxbs�k��Ж��cu�7 ��7,)3դ1�#��5$;9>�q��H����,cC��B�7p}��n�w����v�v��5�
9�4eE�=�#��d�ڌKEDh���ښ��:��S���}�?�^W�Jd7D��)��\� ܬ�����'X����S�#a��u9�S�\��W�]
�kc���s�uW���[2=�x��i���/J�&LN�G���5�f�<�Rˮ���'>�q`��d�-i�1�(_eN�10B�CWM��\�#W�R�ͭY�a�vp�9 Dc?7�1��	C����fz���_����" y��v�55uuiCF1s���k�PVC�0�e�u�۷W
�*4������B�f�f-a�V.j��^�P]zrM����{�L_4���j�S�;�3�?#��.�ZI�j[K;VJp��@��{���.[�:�3}�� ��AuGd2u����y���J8ܑ�Bqx��uJ#���xk���Z_�n43�_|eq��w��oA���64A[��\x�y���k7��>�l�̮�AJt�4F����Ƽ0�׵��|_�CZ�m��Gb�Z5gG0���� 5����������2��P�`$�Gq��[�E���k@�ǖg;tHsh�/�س�ϵ��(ap������申B	�˖.�aª��S]�a�4�
翣zşN��h�y�oXGKm��T"��}�'�x:���F�V�f�h�Z�lΙ:���<�8Q�@@4��Q$f`�{&�7f줴��Q��k��[�l�{��H�`z�����]��gVʶ���Ks һ�K���O�2{���貅�Ps"����W������u=��Ѱ؝��]5�/?�R�~����!�:T�#.���=�g��H�xMhQ��[&Y�z]̙��K��g�y���X�l	=���?߀x��G�H�!�i�S��ݔ9&L;*m���}l�� �sI��mO(c�~t����p=�*��!��<�A�h(�[=�^�"A%g�V����QBB�������FiRi�!�ݨ�rX"6�gx~KAia�g��m`��u�Ŀ���Y8t&��YvB"�2��JYf����N ]y�m��Ě���:�v`�N�!�$��#(vVC#��M��=�~����ǽ�N�@����=�<������K�9u���dT����v������Z�Xrx$�=��sA�R�DE4k�]L�r����8�G�\�J�p�k^_��T�fN�jwy ��>��t��y�?�>=��S���]e�}d���{�����I�t�OJ5;�Z��u �7�_"P�m>�s�A�!��Q*��9��㗖�_�#��j�6P���1�b}_}��5:��#ǎJ��"����l���v��Q�|���U�-����Z�d������ut\k9G���Y���N����ܶ��9\j;L�:C�տ�[�f�yԳP�[�ku��w����������t�gƜj�ۡ�Ϧ��t�A�@ꋹ����}#�:#�Hs��AU����ն��~�aT3:���&*1�����ߛ=K�X=�B��OԞ�
B�1^������o�C@�3�ϥ^;*F���+��<�۶��~�3,٪g�J���D&�9��i6���F$S�fT����e�o�����څc���I5�\_��M�ē�H'�|f��^�9O�ÝD�G2(`��֛��/�.�z��0N%-n�ҕ��BEq+"3���[&W�/�mi���.}�����r�;Ձ�\�r]��N��T�
`�y!Ͼ�n�3i���`Jr�q�֪�;����a����y����\a�|3�R��q����a�%�=�`�":�}�$t@m /|����^KG͛�n�iA\�%�w�Ӿ��)��l/�mr�#�z��E�og�洿���؉C� ��|L}��������D.99:�y�rE��.ywn0�k�-*�/��P�j'�sW<���d??���X}KȋϠ�㹉�_;w��u?�+��W��,��1��ӷ���4���:�r�k7��e.��i|�h
J� >2+��� ��*�>GߨZ��+Q\R�����~=mY��t�eW����ʒe�7���V� ����6ni�l���C�$�6j68��3���pyh��|��A�yN���E�h�3��#|�L�,��z��A�;*�@#1�_���M�>�d�ۯ7}��kb`�6�v��X	Zp��j�`OWA�jtHF}݁��u�Q�P���Е_]��';���r�\q4�z\�w�A�W�i�q��b��M�����?ºз>L���4�Cg�Ao$�L֨�E�k�t��f38-m����!:�F'����f͜�p:��~�K1���m%��i���v�^=�NE:D;n���Ȗfͥe1�ߑ�(߱���u���aܮ�gc��箨ʺu뢯^e�.�
��|������r(r�7L#�Q$E�N��q��F7���;~ͺ����}$��ص3��)H4�Iq:��˖�Pw����Ⱦ�P�ڣ���<���/�����r��F}#��ں�s�m����ثȢ������!��K�T�̊��Di������~�I��u�LԺ�����?~
�X��k�/�	�A������E�Tnj�� �Yy��Lǚ�K��.��v���kr�)$���<g=�Kv :P#�0BBUxqH����>������?iz��+K^%c�_r�%h�)i�:�=k��y�gZU�M��9����N�����P�����Y?w:����?��S�4@-i�,~*�|���7R���m�����b�l�c=�����gc�3�D#��4�q׊Ơz��T�F#_��ég^�#I�5�d���w���>�m����*�5��:�s?�*& �2Ia�Ò����<u�9s��N�<���~�cW��{Z��w�'������[��u�nλ�y�\fdk��MlmKֳ��Ne*�Loݬ��ts�*pfBa���fP3�秳Ϲ(m�J��u�kҥ瞝FN����Eͬ�jt�{0t�e�c�*b������F���,�E�sɒW�U��&�9��1��*>��\K3��zz�7 ��~U�!C��:!i'��-?�Q�0�\��m��%��:�Ω�!Ѫȴ���/y���@{8w��	)�h]\�m�@�f)���%͂����~�x���]盳("~	J�0��f�f{Z�ae�͈д��S'��Æ[[x^XY]�8�ڙ�6a��(��Z���ڀ�[�oA�G�ty+��}�I/�,w��7����ѶV� ����|;ڭiB�bb�FP�m+$>�k��?��v��z����3�%��mA讴|��X��a�r����D>�y�����]�S!Z��m4���h�_��7u� D�;���;�^�+���{o8��v� {YSQDdXG���w��㏦�|�c���u.]�hv˭7�)�����4j��-Bx݊A@m�8�>��8(23ܒ��Oݵ"P�0fm���ec�H�����Sɡ���"��6\��$d�8������v�L]۱f_�쒫h���R�Y��f��K<~Ŕ�B�԰��$D�z�"��|��`�gE�l�Q��f�����hAN��$:֮߄�][t$D�_"й�㼔x�7����E���Ď4�tE�l3���iu�.��*~7�c�ЃJ�]��R��4v��t,j�W��0��1���Id�#�yw`�Y�7����c���<���J�_��ix0mmݔ��,��*	"���0�2���N�����rwZ��D��1�ӌ�9���@����n�@I:W� x���cy�ե�1�	�9G1��T�yϣAw�q���TakT'̪~�̿1k��_�0nܛ�1����ޯ����]vݓl�ϯB����7S��iD�&�8�KB��Z�S�E�O0��x��� �y�~u6z���������z��t�՗��vEz���ҏo�/?g}:�<�U=��lŁ8Y,�M�L��,��|+j�#������y�����nI��*2��b�Iӧ!';)=��#�c���>� ����3
��Y^�n����k���؜Z;�Қ+�Pꑝ�뜫N=��1�:�F�+�Jm�n�x�s�[C`"G����@��:�?fi#1�eٲEf�Đ8N�mR�Ma�����r�۱cf�ؖd� ��̬�fF�<��s�{g>�i7M�4m5�D�������=��<'LW�<��y��e�b�|ڟ�Z�����B����T"�\�������m��q<��-J�d @�r��R�R�!�@T��S���+2��ˉ�q����魥�����>�4��k��Ъ�ƕ��2Ie��Dݖ��g1nB5h$u�P���|����zk���)ރ�ПX��@�������A��K	A-B��,2�"�i�U�^�|�I����e�=�~�FqQ+J�r��^yy��1/+/#�hvg�^zW���%$��R J�)���:�w4��¨��x��#�$v7��1;[��G�rw�6���'`�7�xRG7mR�9c�@�
J( ?����z�ة��>��:�t�p5m�d[E�kZ�Ĵ�>ƄJ����R��j�p��Q��y��JF���S��C�u:<�T�3F3���6f�=��ӽ`Y����=����f~�&����f�9�2|�ԕm���cʣ��	*+�����Vi�<+u���|2�8��1�:q���H�\�9 �qK��K���^��JcO{�1fA�b�^^RP��뿭c�3h#9r4�`5/��������K�''@�
@����w�D�o���u}m����@R����r�+}�̺g=Db4  �&��p�%	��Kڠ,+L��� }Z%�Ãρ�/&(F���I:�I�lC��4e
��\g�{He��%Tp�5Bz��T�$�L�?����w�+��q(��� �﹁�P��Ո@������8T;�(rL� cXN#MpjD����=	v氣�*�f;kڬ�?��f�����=�+��[+���ŗ�k#+F�2��p:����4%5ʁ".C��u+`����E2X&u7�VɡV����K��o�f��e腇�I8�q�������N�k:�r�}�d�H�6�ަ�A����#U��\#���E�U�q"QP���ęK"��gȐ+6�N�u���M�f�Dlz]3�e�;��Z��ό��Z�0���&���W���-<�a�Ad�r�N��I�z��i�Z���,Z|�;]A�]�]�f+G����&U�PFx����Fd��PʺD��lO�&ͮ��Q-f�)�
>�{Y{�&�Q�a\{�釶��}n��u�o����o����I$<)PڌB^�yY�\��2g�L'浢ݭ�5��{g���n��䡰�G��}�ꂐC��M�ʅ����eY�����8S����[9�b�Aa�X{����J�\\A�u�ܼ{��m��eN�K������m.�І�CF��~ƚQ�ӘZ���p*�e���Lq�JI*k�� U_51d�Z;�H�xKaF�������CiH�Ze�!���bW�C\ܡ���y~L�;v�a<m0
A	����zNkXNxݺu��K�I���Ñ,~.�z7e��QYC�ZY#=�d� N�}�_u��t�3rd�֝��;��d�+�^aS�V�TFMٻ��[lÖ�H��p�n�A�p�+9`�E(W�Bae���j����ffD2yy^Y�J^��^�s���&`y����3&� �ΓnM��A�ҁ���ұ#��mI<wڼm�Qp�������}�������Qg[2�2~c�y�=�1�t�����p��>�h���U��!�Z���%��D���p�]Q����>6g�i���� �}N���Ėf�f3-K//�\t���3v͵�����SϬ��U{m�E���!��'X��\�L��rFSҮ"J}D�_���y�bZ~g&�s�\�{ﭤ}m�͞?�ֿ���EaVr2��d`�;�t�N۳�C{�W�<z��_0ߍy!�]�A���,���
��R2}�yF�ɓհˑu�<��mg�EN�j�+Եb#.�k��&��ev�,��<��>�[�\á�����j�q�S��CwC�qۆf��E�{�\С���L��R;^�\.A��X0��x��\�h�p��d8���Kl���VG0ԥ9���競���e���S��	DC_T#���/�b\�u9Z�I�A\��k�d-8g���-��T)�o��a;�q�O��DX���ϡa��&˖/�����
7�> #�Y��"��{���VyY�d���r�?��g+9����[�.���Տj����a��6�Pӕ���DmK��j���1�����+/Ad[�@�7<S������/`�}!�Qu�����ڕ�,�P����_(����eo��ȍC�B���4�W�	t��L0gi츱d�
|=��g+����_�q.Id�G�����m�N؋a��v�|�r����-���F�8��(�5����Ǥ6A���!,z�0OR��R������a�����3���5kl�ڏ�3���
�������C۞8ވ&�C?�U*Q��~���V3�h�g�TЦ�!)ȧF<>��Ĵ4�@��8�B�f�䟲ֺf�*J&pBZ8��P���l�B�V�=�2�PW�w��>��D�H��gf軰u�7m���'ß���Q�[gE�w��A��@P�����}��7�3g.p�ُ��
��;��|�۟����3���u����$�Q�3"Г37�Le�Q�6A�� ���&T�B8�N��5S9<ID�2�{NjS�,B�C>v����������Ys���Z������ �?>l������=��傊����Ӣʙ�u��-����
;BOp6}��D�)�Hf���|s��2|�l[�i�͙:	� �:򐥭>xԃ��zXL6����w�w��HTO��<f���Z`�v���l��YC�;iq;Fo)u�V�_J�<S���o]FP�S�V/��e<{w�o��]�ˣE������$�V_�X�rB��sDKrn��b7��
U̦���0�G��rtA�ɺ�ֵe/utg�>�h�m��$ySA�-]��Y5�d�3����3ϷwV�"C.tƱ�L���s�l�̠~{]���p��l��0��e޲�Z�Heb�+0j�a�qk�m��Q�֚��d���	kRǅ3��X^)	�;�.p����տl���Ϸ�Bz�5)/XL��G��/|ў}�E��G<�QP�C����W;[
A����!'g-�U�(���Y����{ݠ%���vP�IQ�-x�*ֳ�����w@��|�Ns]<bޗ3��C\u2�u톏b��|Ζ�s�����p�� �˟�7�GX���JaMqKk�΁$�!p2lH�M�0ŷ����9��	9q8��Iw����C��mp�,�B�$f�G�7��J���6D�祯��I��C�Rm�mt�@�3AP4@(U	���uV�L(!(1C���HNX{\퍴O��z��W ���]_�-'-��9��\DJK�J�����	�!E�L%�n�vH'>�Z�;ﭱs�=�@*�ϦP�g�eɃ��d�"��K�iP�5������jD�N�_r�?���5ww���d�S
`�d�!6"e��Ю�ڹ��U(��;� ��?;8�w��&1�p��C���Q�v�k
���PP����ݱK��<��S��y8���V��͡:|4�O��O����|��*�*�0ȸ@d2�S��Sv^�)5�.��a��Ci��S0o�t䔜����Y��jSJ�piڕ2�wW����^�R���+�"��_x�fNE����M��e�u)$Pܑl��C��lD F�"��o/[fG��yܖΛn�q8�`Rk��޼H-+�=Jm��9���]鈯Z�̊��A�S�򓟼�>��������}=�]8ە�R2T��n���n�H����2F��.�~F�a�p�薫�Lu�x�`��u�Uk�V�F:��?�M&�bt$�l� �%v���C�1������"ƀu� �����3|g7��m[v��I�^F���@S�t�IX
Mv��}�t?�g�Ĵ�?q'���UF�E���bzl��-^7�믿Ik�0�Š+2P�+{F�\>m�d��Tꂄ��d�fO՞�vC�Y��	Q
�o�ͳ�ʄe�;����-w�����"�u03~�}�+����qz��H3i��(�\g*Ն �g��.� :��u��u6z?�E��P�гV�Dm5tn�A5�QЌy}(����<"Ue�N�$��^�@A�pd���ۋ�L=e�\�A9d��9V5n�K�@���V�A��U�;��T�8�����<�'Ù���� q9Hu����_�m���n/�^8�P�vXs��r��H8G����y�f��e،��}|��S�y{�ƽ���z]9w9>���[3�y�u�(K�@�c�=�_fw��i�9<Hx�Q?����mE7`#��o��vЖ�p�����[6#h��g8j�6e%��^/�Hu@_,B6D�1������B�)���c�5r*1�V����u&YI�Ʀ�m�� �Iݘj�B!N�?c[ ��H�e��K�C%RO��G	N�әlYA�me_,qh���1�G�9nLU��y���V��š���K�n���656M�����H^_�Q��\qD�O��D�4E�=���K�M�I�����3���%#r5-6��L��{�(J�)88��!v�ؖ��a����}�3l�9��F�����Ʈ�b�E�XX�t�ӛ��iC3>6�HOyC!�3�2��sw~�V�)�)p%��O�c���Y��SQ�[��u++J�5l����6�>D[>8���T�B��<��o~뻌f��Ø	۽ֆ`�i�k�j�,�{B��ѥ�	N -�@�ގ�B�.�ue����w_}}-��p�OH�#c�G00rD�gF�~.�g���u�D��ukR�|2��z�'�){��AM�}k4d&-z#F����K?���v�W���}�Zl��;�5m�fg��ȁ�{\�%��B��w��C�裏��Z'�f��z,�M`���r�UU#�7�׀�O����YG�S�Q{~�!~*8}I��q�Z>G2����zm1Lx�=�pb���d'Y%��K����E̚9��94;e59�H�Y����_�maRA�k
9���",���|��7Q�8����iPP3m�]{v�4�tȵ�"��eNӺ|�!Co���gV��it�M�-�B�t5o���GU�x�@/���,r�jÆ���!�쐬g�f-�c>k��20�A�40�k���8���X�i{f.ď�?�Tu)�ׯ�7��?�� ��Ǵ��%��y�`,{Q��σ�ni�Z[>�Z��O<��>5n�xI*9c��r��"�ڈ��u?~�0%�mvA�F%�۹s�]LB!�d ���j`S�Z��|8����^�u�$%��s�I2�s���0����$�4�B�%�YYF�������)�tX$>�QWKd�@>�6��g;�4����s�k�>���������V@��:��	=����/����ٿ�<W������_�������}d'E�g��C�6�ZIb��e�	<
��}ZQ��u��2�RÔ)S��~�;�y���Ǽ2f��Q���9'ۮC� F`FmN�8�#B�k���c8��*T��C�����2u�-���ȴ~�\�}ϼb�N��ys�/B���c.5cT�Z5��[��N��[l��B����ΰ���(�!#�����a���=�=��hE+���Kuѐ�����|�s�#]gO?�M5����v��1 Y	�dZs}%Cc �d����5��򈜏�HSe� �^w���]D":���t��%T������������M��=���kr©8��/�ܞ%�9
�}��i�;w��x�'�G�MڹfϘfׁ�H�MN��Oy1��)w�Ū�!"
:ϲvg"c�Be���߭�٬Z��M�6�^f8���B9G��R�Frk�m��ڷ���={��$�$@�V7��N!Q�� ��9�b��z�k�^W�QF�(^�t���@�)U�`}�	��Y�2� c�\�`"����C'c*�lC��}y1M��c�a�v�q�f����M��r���7o޹h˯vF��vV��A�B{�3x=��=CV�*
�t���P������}Ѿ��#��Il�o���p��D_��>=p��uw����b���{�{b�'�y5�����8
���h:X�$�r�)qF=�=j�Ţ�g�
O�C�F9��.�^{A��E��K���^?)M��R��o9��
�qBx*H�S����>��!���.^��� x@EQ�%�#ʌ,p�Ͱ�{R:�����>K"So�=�Ʌ�}�C�(	�D
6& NȃQ�I+)W��2d`4���E��E�O�'��O2��h,��f�U��W�P�/J���^���]|�E��y:���u�
|���B�������>6E���F<6��ӆ�C_�;ijy6�rؼ�H%�>�xj���1X�R9�H��<j��@�yY��э���m�$�`�r�<
s�TE�1~OmT��I�Y=���kjT�kמ���C��uoڒs��5���c��ϒ�塞4 TZ���GҴ��n"�K��!�4B�i}�8i
�+=r�Y=�� �J=�>X��axe��y)Q�V��������5q�����od��d�?`���2��,S
l���RgoC�,��]��1U���� �����R�ʰE�y��h�	�3>�N�b�������D�3@wʚ��Ȫ3��Ofc }
���>������#����B�k�������7b�3�%�~�$ϴ��旅���UL�jBc�ֹ�}�3ꭢ�{;G�ɢ�"����\�tj����>��2�~�]$>�t�:�_�e`�w0�w��7�|���J����4�OkR|�#_r���?�Nb�%;3
�#/�@�jqSi&�}"��F9�4qF"�������{�u��%g�,��1��-��?�MPPy���{��Q�Q�)T�,�	ǌ�����Sz�ԓ���Nn�8�&�e�Qæ:"&��P������0*��6.��29QN����
g�g�;rLQ➊�u�������nR$;��gt?*�)�k	:_c,C�>Ȭ��ԧ绞��p�!@���]�quRh�|� ��$""?J]/HѦ��w߳7�\fw�q�g���׆y�� RD�C@$t=*��`��,s��JJ}
�͛���*��;=c�R?�{̀M��ք= ��fj�=��F��$\5�.�7����~a���d�`�9�6�	A���O�e��i=��*����6��I��S`���2>�����|ۅ��u�@�����f���9c2�z)���ə���v�@:+6�!�:X #��C@�L6�f	c0?Z����l�k���U-T2�j�4b��>�FfΞ��g'BLS����H���HF_]���r}8��)� u�l�I��o��{�+/�[o���Z���m�k3f����	?�:�j�Ȇ�4��ľ��o|���ŋm$ґ�����e���eb�H�2k"m)>ͪ�h���
�Z ��B�8���9+i�l_s���O�g�F+�k�YJ}�����:,X���/��8�\���9	`��Y���(BW6C����� �!V+R$���D�#��{��3�k��8G;Ȼ�/����`��/�D�>]p#�_R�F�j�fFImm��7�5���#3h	-Qjru�@�Zt�9���}� �a��sS<�KV�j�x�՛ɼB���n~P�$����e���xH�����-��.[��� ?�bb��^�y�w��ջ�8{�g�6@��@�Z��O��$6]G]
����@5���z�l���X��|���u
� ç{��I�0W=L`��E���I��
����p/��ĭ>&x�oC�N�=k��[�u��BP1����G�A ���>B@��&tKG�L�9�C\Aj(�d��!���ӝ��j�w���!��O��g�Yt4�rM}�Ygg���Y3X�h�� �P������^r�]�ꩯ��AA������E��*QB��w����pD�����wm��U�9����~'u7~w.���td�wކ�9��!>�'5B��}��^����zw�q  M��
��h����hgdjo;�-��,�@��(�r
&�J��Gew"\�X��G~��kIl)��1GIyd�,Dhd�:�Z�F�g#A�x�d1f]r��Ó�u����������4��ު�J����\���q��!�L�9h�G�:�Q��k��E5,eBW�zg`��(�S�"l�l�gk��s{�̙ԎO��]�l�~�R�z;ο��K>ݼ����(��GP��o�Qį�X�evW۞�Ȗ`�/�`��R�~���lǏ�\�Ճ`���fx|�fWC��~S�����6�j�1�i
��g��:���&7���o�^Y y>]M���ʕ����u�b�6ԧ9�Ca����������o�c�^9�W��D+V�[a'd�&���S?��W0#4@}��{���zܸ��ݸN�g>ʔ�a'��eX����d�Z#;���N�~0tU7L��e�{�}�ѱ%��)�	�����G�D\������?�6���㭹�!K�QƧ�'�쭷�ۦ��������*g��{
f^�v�oA������>���o�8L��2�ЊaN�K�Y�\]:�o%bw�wJHFp���.N�X0x0
��B��A��?������é���d���zdA�m�|��ȩH�FA��*1�3�m�����.-��b�� � O���NSP�9�lEl#9��J�c�Bk�H�ߣ�P���
�? j��92���:7A��g��q:��/�VB�(&��z�ؑ�����؎�S׋ ���&�iOla)<��1�Z8W>�0���Х� �7Ϯ]pF����[{yT�R���% *��v{�G�.<�6���&���g�nݘ���2��C5��L�\r�E�o���R��m�J�)��կ�����&(�w�%{@�@	�?W�H+6Aj��J&XI���)*�t0D��Ć珱�t�=7=g���gV]Cn:���<����lܲ	&�M�6ˆ��!�Fe/��6hmQQ��gL���~�2V������+D�!��ͨ%E�A����u�(��n�B$ ��YJ�{���z�*B����Ts��u��i�.�d���b���(��Ǵ��)�F���ka:���c�2��Q�n�w��ɣ�^OT��S/٫?|H����y'N��Ʈ�P��t6��A�Z��鵥q�����73�̲�|���#����1��ڏ8*����|Z�$2�l@�P��NՅ�VJ�Nr�I��P���ӟ��^}��[V�WT'����4�F-3z�\�#*GXe��.�����G����GL�}�ZzX�8s�)���! �ܼ��$B��|���>P�6H=�d�p�>��!i��V(� �+���ǞA�c�?�6f�����1�E	�x�3�/%	�[�����`J���ϼs灨 �JYDӴ�V�|QP�ܰ� ���D�k~��_ve��{�2�R=T�+h]�KM���G�����z�"	*cu�J��������է��H��Os�8!��}��,������qTb���K=+v����
�k���O��P��Q��cuv~F�m|1�]���E������S��7��˱�9
6>�yƬ��/ܡ���yU<M��!�M@�J���Je	6������w}_v$.A��K�n8�ʱU<ߵc7��i��q��er#�c���f���u��5�7=[Qh"@�tn���|v��W^q�e$���0����o#����,��s�k}���ʱ��m�˯�"�ѳPۣ�_z�E�8L��C���ju��;���_��J:�"4�+B����J����Y�te��쑖�G[c�_�<W�Ձ�Q�+D$�(��3�Km��[@:�X�	�O��D�y�!��I��=b�Yg~�%����������%��v#ʒ��]�-?ʐ�P���C�Z)cg�rX�^a�&�v��L�&-Lη)ÆڤI����n���D �����#��)jY�?��k�A�D$M^����6��Y�:b~j�F���!C�`��]S�Dѫ!���ZD���]t酶���d{b��M�!��ɡ<@�q�uS��$�T��������nb$�ۨ���3}L��(��� ә�[LPpb]��<q�ƍQ�L�Z�0'S0�0b�U�ܜD`2zD����5�1�Q����MW.�c�~TZV��љ<�c�DY��p' M���]�zjR��G5�$�B{�'~2�:�<;��}���JW �(3�׈�n�;��`�Ӹvw�����au�ZO YG�קN���+W��S�=����lK�$%�b��$�iؾ~C����8�r���uq6n�l[��tG�]~m"/q_\���f��l� W?����U��	�m�^���k�����m���H��y�4	��¾���=�
@r�����(�սy��r5���cO<��\�7" =Q���^|�b������n�����Z9
�O���.?����TqM��"8�����H����Oxo���^�=���z�[2�!;Wp���� ��A:���Y�R�-'�^���^����P~���%X �"��"!|�5�	+`V�}�;�ψ.��!p1J	�<�ܘ1�a����.(O�E�gE�y{|(��!0��0�%�,�}���4����Ā�n���a�є�*p;���`s9���V�ܖ�b��#G�=v�m����C|.F1Pm~��u���՗^m�Q�;ʰ�����Ѕ
鼵\dSn��r�x\���=�U��d��`�+�Ѐ)&���Sl��G��^f����f��D�`�1�U�V���}��y�y�h�2`����aQi I�$�͋�,�m_ĳ����9����6H*]'���4��W���=y�i��B|Ou$ĝ	)0���LR�aǌnc&L�g���#�-B�K��e�*Qm���~`;w��Ģ��G$<�y��(�x<�Q6~��,m�}��h0LrZ�sү����f{�mW1X�TD�"{���]�]O��nM(�5r?s�,���zh���;���k*�đ�f)�o�y��E9����j ��6*Z]8M����+�X}�3P}�Ir�e��l�y�Y[�a��p�%�bC���{}c��,��$�\T���'�3 �Te�2K�꜑����\S?���Ԏ���2&+ń���2]�Z6�icQ���3��/�E��gq��%٩HҢ���[����x��^��{��k���@#���sr��1�S�N�s2#U�x=�IG��B�1J��U��B�]7�A��r@U
��߂R��-c�JC �A(h���ȉ�V&w�|(N��;p(jE��|m���>{9��mЉ0��/F���-@�t/�d+��2�]�-�`��?g�mb����I$��Ulz���R��.���TYR�1r�ɩ��3���AƄ��n.�^A%3�E�T+���>�L��+Fnb�W��P��<�@�?� �:@������������sf�2Ru~�-L�2/*�jC(��lv���0�L�:cD�s1!��ٜ WM�cO�^�F���Kf�-yl�Ѥشi�}���%8�w�/X��Fz��]��t&�c��T�m����W0�}�����i3�����z��M���?�()��:���,��l���GV �s(ڛ&R�.$�XTbb�,`�V�YfȻ:����;����Hx<�r%z��>x��7*�$�Vx��t��,^���^��_�+�Ks�&�m>��%�y�1��,�#4�P�o�����V2��1E-���4�Q��';m�z4���^��uܨ�&w8s'c0�k�Q\�7���B:uń� /�wedh��@�|dh:����,ۼa�nw��W.���T��Vڮ����G��������h<�m���l��G?|�a3qȩ�o����/�o~�NOYrq�{77ظ��q�`0��sBi�v'�n�v�0�%�W�Z�E�.��~�����m����v���6�Q��o�[��hV�d�E�V���˼;���Lzké��/���^e���ٹ̡�4��Y��y���8 ��D������x���ҽ��J�KSȈ�2w]��<�Sx���@�?�o�T:A>�?����#/^�<�P6K� -�B�n�������ui��CP�Hb�����޻1����Ȍ�r�V��؏����]��<{O�
��#c9�%d� .jj����w�3�/r�������Ơ�2w��^��Go���N`����WK���H1N05]����v0�Yb�淾���6�t}���͠���`����g��`�]�ϝW��?'��M|!(	."�������l�J�z&ԎO':����kג�TF�|0�l��õ.�$2��}�� G"����8��s%x��ل���l�	�/��+H0�n~�g?��R�j+�,!_B ���[H$�SF'Φ��	2�x�e���69M����[Y���G���W51��g��ת|õ)�lB�|(��
P�絸<�JNY(��v#�CiC�k'�	yi�6�h��%[v�ꇗ-�(=����|O�?�f����^�4*Ja�)��p�#���8��_�
���n!=5�]���Y���J�'�.B�PG�,��� ��h�qIt��6�t������ϻ3W��F��߶����I�8#�Nu'����}�g=!{��
U���g�r�e�]����.O�1��H��[�p��ζ3�o�K/Zd�.O�o��v�̹֋$i;�/�π(7�V��B���1���m� ���߿�]���V��^��V��Z�HL�� 6A�:�{`�V�boB�Fh���N�g�;�Y����d�HDA�+�Ę��[��0��|f���z��:������P��y���P�I!)qt?�X��vл�:rQb/kl�cG�Y��G��0n�§�	e�w�q;R��dQ�$���Ixz7e뺶��<x׻ށ^�2�j�r"{ʧǩ�[��ڟ�٫�HA��KD�q�5QJ��dk�{jIR{���w#���L�:����������;ڋ��~D�o�L7���j�ss��K�>��\�5N��m�5(P�B�4B�#�;B�Vn�;D�V���j��S���;���}w�Zp�7����F�j￿�.��b��S�g�v���m<��Wݳm=�`Z�稼�KY�τ�0n�_����%:���y(ǩU�65e�΢�QS�B.-��k֬��2у�:/����:B,t���5��;�	ׯa>"4z��V02�Ǟx������nB):`\þ}�w4^U�"h\��'N�ڏ>��A"Ġ$<�|�;�ݽ��U@�b�`eS�$aE>�w�- �Jy�3ăh�"5}��>�\�1�  <8���u���}M��|����,���.)a΄��P�g2�bB�>B�+�l�_].�eWkT��~�R��ӧO����ǿ�
�Rz~NfJNJЮ�ɣ8���Pϒ���GW�r�H$�f��Z��H�p:�l��p�)�4�y#Q�g�~0����!Pþ�3O���A�ʒ:y�p-�<!S���=�1��ol�S�ԭ�j�I�{͇[��}�,����'�nVa�^_�"Գv���%���f����Z��� h#���54~���	^@:ơ���X'����]����$�q�P&���#x��G��ŋm,��i���A~i�����7^{��������gs���?z�2!����ֈ�d�߭^j�M7�h� D��"t��@5�6�[`4kpɀ�d���sƴʱ�;�D;rqp�RGdh<P!8�T���wV1���;����Ř����L��rY�x�RE�Z�{��?*�J2�v��lȂ-MuVG�A2��.�w���ߍ��=��s^rN_@���RX��}�H����j���}�~���ĳU�Z�O���3���߷�x�@~�v4�UP��`J2��Xo��&3 s�+��9!0�PM����?��*��%.����<��t?<���ӽp5�?0���!�l�}���T����_�������� ����gF���R�:�C]6q?����s��c�1c'�Q����2"��җJ��i>��Ԗ��.���L�<��3�&�>��&���(��놠(F�Z[����։g�Z��O?k.\L��w�ZHq"�	y��g��7�2��um�m;���W_���F�H�({]�=2��^_��J#b�K��g-DA�Y��E�ܺm��V�m�~KHq.�̿}��{�8��2AۺD̔�q�2�к�`��;7�+E��Jt��c�[	�2�RA7���&N����L��q��){��������/͡��{r�ν�2�ƥ�&B�ZGvm�Ꙃ�������h1ٽ{?Qi�tW搑�(G1c�WK�:$�9(�:R�%'����l��3�W�����\7����=�Z�͚��~N���\�ؚפB�N�Ñ��`Xz?�㓙J�̪^�W^|�F��h�/�ɮ�	�jZ�O�fgW��������� o���HcZ�L��t���X���-�:�:ܷ��}�_m.���
Ⓝȥ�9	C�����<�q��|����J����E�a׏��|(p;�����9Z�}(ӹ�%KF�����2۽'��"$#�,^���*(WN>d�����Y����؃D&[��k>��xR��1Wf�����ϧ��B�l��b�:䔕%K���3��U��ʑ�;{��W�� P�=P�ҠF��G���k��6
�8&�'X�A]]�;9�y��Q!��u���Ҡ�n{��z�q���<@�9�n��4�'��&��{��=�Ю2�!(
�']b(r *�h/K|H���ڸ>v�@�r�$X�R��	�ՠ��e�P����H���Z�mf�b�w� ���|��^�j44fr��JH��.&7��Dvb��[���,�˥�i��K����1_%�[���(@�m��L����x�SȡSc��t���~G��z���r����Ӈ������OZy�B~D~SЩ�^��^���H�p� ��B�)����	K(����)���/���l���-Z���,�q\n��7[F����3�9i��;i߉$lVv��d��$2���`�T��*�\�%��;nQ�NR͟{�3���<��]�SSՒe��l�?����3G���98��)��/T|{ո�M�|�u��
�R�w����X�i�YlV�,�s���`-	mx+�4�ө��[0i)��Xd�1�!�������<��

����h���-L*
}�1l	�ϑ�r�����V�rFs�ԩv����{�<'����Hnl��FGУ 8M�J�:��+jQ�����vl�7m�vт�6�����l���욥�Z9,x݂�5]�KQ�����!���R�2l6�Y&TM����;hW\�k �����dܤɶ�	Mj�SQOۋ��j��;�(�>��;�Ǿɾ�O�3�e6,�C.<{6�G}���V@A֐	�*a�a5�:�[$X��KS���X�2�B�������Y���e�Z�7�ف�}	(�gtNLS����6�q�91� TB-W^k��k�h�6Ė/�y�I7����i|�|�ZۚUk�7��y��J`��P�֤+^H��ճ��a�p&�	����uǞO�9)��[�&M�uK��i�=x�����aes���eR�>e��(���xq6xo�q]�tNge�e�ז�h:���!�]��!p�PnWZ�@9d�A4E�Q}ZeU_��	4Y.8 ��8S.D��e��E��@"�B�vL��'�%�%t�?�?�o!$:�r�^^Qi��i8ɐ�"��mb^��2�8+Q,Y\���"�N�L�Tm<Bo�	
tm�_��Jt�٧P�Ӹ]���M!R��%Km��I4��7!��x�>5FGx�o��K������C��D���l�Z�n����|�F�>�ش��6
�%�C	���8
L���m�b2�g<L��`���l�s@b'����|D������7� ,*�(��]b[=w/\x�κ�_��x
�s��7��ض:a�X��=�����/E�__NY�A�� �Ӣ��ލ��if*�V��jAB'�r������� �/Mv>C&�j�A^:�ÇU�:��=�Ǐ�C�mʄq�E�B��8`�ގ+�y, ㌅MK�bjTٹ�����. �>���V{�����������7[���<�������J,ƕ�D` @����j�L'bb�,Ku�.�Beڝ���͚;�z�Q�{���K25Q��0���OY���1d���:KVk�F$��܎���p�}�w~��j��w�	�C��cP/��Wuؓ'kh�#{Q]�Q�
E�JֈP����m	�;�9=���fbU.6���6���O���&�=��o�뷪#+�S�w���4)�Zy2<{��ȧ�I���_Dk��{t� �/	�Ȱ���Z��$�r�'ɾ��o������A���,J�\{��\*�OB¼m�x�$��N�+q�W��q4�7O`v;�P
:\���	ym�8m��b��=�ɂZ��.5,�+_�C{��+�;ɐ�t�4Ɠ�&�����*��,������z;����,Z��z0��5a���x�p�A�Ok0��W��;V;�Y���%�!��+q}<�wb�ݳr���xz0���B��8����o|�� S�C$��s��iB޼K#�4�>�}�3�N�����sϹ���>w��눙3�Y�`����kQMkYA��`�k�K���7ޠ�3�ɛ���>���S�W�tV�,]�k1�uݼyjv[��OR�G�l\���M�]�5�F*�rҮ��پ�t��4U��:�O=X�8H�� 'j-L�����-�Ե9y99��:󟳣�9��/ԡ��W��y�� ������hr�za������@U��@�+E�?[ۛ��N�(���0��L����8�T�Ӽ~l��^�&HΦ����.C)F����)(bivt
p�[/�l���s=��Ǵ��}�V[�vFc�]� �ϊ��2Qr����n��?A�E������&��۰��fY�{�]|�T���Km͖��УO۱��-��v)���F� s�#�)&�d�'ʑH���B�"���/��8�l0��N �6+�0���$�sc7���w���H��ȝߧ��R�����fw~�N;o�Ev�C�؛�l����v�D�� >L�EW��Ú��u��s��6�q���w9��3�n'K�)��jҪ�'��wAj7Ԡ=��8bǎ��,�R�)O&"�7�G\Y�r�9gx���h(�p���D7��{��N��r�5���ē/����AV�S�$R�:�#ʒʜ`��<�$�c��n�����.�d��z���L�-�T�f
B,m��=/]|�]u��V:�����u�"�v�p՚�~|]�2�к��P+�����¤������}�1bSu�^�[�d���k]ci��VAj��K�:�!�V�-��� ����-���)�KI�M�<u��g2_ӽO����m��@*�����]L��5�D�o�vGy"1��HD0�JX��MMu�����1i�>���<SW �-�0�q���ל�C���z֝�і��N0�s�A]�D���2{�[G�um���%8�z�>i�r:�7"��A%)��R	��>`o��v�6C�lt-�t3���������y~M��6j�X���x�Q`����B�I$Šb��o��;��I��,�!������8ݡ�T�Cꑙ� �(}�uk�������CgPs(��T'T��5�]5<o'�x���z|�Yپ7]&�}�y��ϟ��9�2?���A�l�y���T�U�_�du���!�����jّ��B��Ym���m��ct�_K5��.ث�lP����Q��d@D#pkGoc�&�Gڌ�ȵ��Gd&��%v���8Ԯ�����NR�j���mD�E{�1���*�Wm=��X���e�;"����
L��<�Vy6��'zh���������Ӗ^t�}���6���I=x��;{2�N�1������ �-�`b�&��D0W�yk3N#�Ϯ��:����7޲ŗ]��q��ﱫ�X�ٕ�|�7~�z\v�7�aH�DaJ1M}��=�,5���
��j��KYKmOoƻ����-ː�2���惼���9�Zw�vx>.��<�P�!��Dh61덳��ݝ~¿����"5��q�|���c�X������>Gq@Sd���LwAf�%[N�-/g%^����ȑ��嶶6�.@,h)�-�����,T����[�wLe�g�<w�$ ���T�opX���j�b2kϩ�}*3�0C��ݭ�0�u���0gi�Ut?ii��_�?�-e���L���
E�V�S%F����=vǧn�����ܹ��!�J��<�.`r�doS)ʗ<�Q$�^�e�.�0��ѿ�4#ؙ�SI
�Kr����Ã �3�GCk�췛����̙���)���k���'�LYy��W`!"�$���G� ���b���j4��ɧ��/�ys�:�'�6�$�]�y���}/I6y0��Η�Ld�!y!�]��k�1�A�J�g�m�0� �G�赴.*�il8�y쟒i΃�(�Q+�,�$���[�Wj !�s=�x��<<���G�mB��_Wu~�,5�G�Y3�?u�	<��_���;��G��[����w��V)�yLn�V?�m�L1:D8����sxs�\�;1t��2>)w�K۠&�f��������+�4�"��Y{$r�Bվ���Q�1�C�֏"�r��t�O�,��:HV���~��ἄ�-�m��ѩd�H�������*)'�px۝_jv��7����.X���H[��k��^��^���6���]�����'O��U�a�"v�
N_���/�̉uC�x٢�A/���;���r$Jt����<��yd�zӓ�����\8�G��i���,���՜ f�����h�����L9�R��uu��RwWO�c�"�Aޢ�7�2ŭ��u�D`��;��Nl���^����g~��ҳ�c�p�Ht�e�Ә�&�� �Z2���e?�*��ژ4�Le��<{��|� R�L�Z�qɘ3=���6o>5r�����;�X�+DDt�G/ѓ�}ܝ�i�
)K}�ypRثS(S�./���HNP��Z���d��r����IqCTx� �4O�%�*��~2$Aۊs*D,�V~�נ�A",�3]W+���N�#�O=@q��3j���I�3��t'�}�WC� Q�p �E�E�82�N�}٭�d�e�^6�\�d"��$�ה`��m���k���!�f��ZOca����P��g���m��Zf71'^�/:����}����v��f��}�ښ����΁�Jq��f\i������ L�&4��P�:h����Ï���D���h�ؓE�+���u{;%�UAc�p�'�|�����5*+&��Ǚ��3�J�?�lݯ�����(/�f�qԟ�~�*���ա�����3��~r_��T2�ZdwlM%˫�=�݂��Hq��r�����k�z��0R����>r��2w���4�*ĦPàf�k:�.fϞn�岔�:���؍\5&eNK.��닛֮U� H���p��Kx!��^B_T>5�265���ۼ_TLV9{���T�H�,-����:��¸Hw�"�8iLE4���y���O?mӧﴋ/�ʾ���؊w>����4�l��� ����<V���?9ݏFV:�����u�JWfdո*�O��$�b�k]4��͋��/*Ȉ���KD�Idb�
��/ٷ� ��K��2�5���1�����Y�V�S�Y��{�j��t,�Y/�E�� �p'�9�*�x�b�#n-t6tTGv%�ƙY�O
�L? 'z��VU���\x�W��ep��ws9~�Z[A�����"���O��0��@G׫ �e����K�WC�68t�'�B=ڙ�|M(G6(՟����͜�5�<U���d�`�徺�(���!Z�.8w6%��.��=��AƋ/\������5{H.��L�-.b�0��T��X�>�M��Hh�.�jC-׹+�>�[��4��9�O��.�X��mr����D';�Db[ܶx&�⃏p��1��k�%>5ƶ���A�g
�����ۂ#=G*�+��F��U��H�_�
E�q�+����3S��D�y��,[�;�����"��F��]�M����:�O���>�x$�+.��rM;3����.�  n��@�?�p� ��`��qm{)�)Y���RO��0Jd9�W�[��5ا���+p�8�fj������d@��'qb��/̞���@ڋl��{��Zq�ت�����k+�sq�7����5�o����
d�U�Q�S�d<�ޙ�3§_�����JG(�9$��UO���|xӥd�8�5��i�>K"�n����vF��괲L�e-�q}8��e�伔�PV�]z��ԷE��Mc��Z��Q	vȘ��?�3���w��}Gl����L-|�&5 CN @���FN\��q;z����2�;�ԽdԺ%�n�;�(�%�Z_6�F�9���Vsp��;od�d� �P��x��Sٵ�/.�#$�'ځ���G�V[IYLಐ%o���8��`�S����"r>��������[n��p�}�)Q1Į��J6ϓ�����9�����t���Z�jЅWG@/�N<���4���wԪe�~��ر��vA@`�Z���zq	ѳ�g���#'�s%*"]��~���
�m�8ۤ9���0A��&�z}6c�t����X6���k~&8�~%��3 !�����a����O8���yP}�������5@C��G���y�Yd��f����c'ϲ��q��0ixHp��>��ҋ|��T���P��Ju�A!���B�&O�B��4'/� &8,&���-H_�/�O����l��@!��O|vg����i}aۅ3�ǘ$�ʾ���ڬ�A5��.��s*,L[%��z'�* �R�ȱ����V�/_��f�w���P*%<�-}�]�wq&�ˋ[P�s}�gl6㍫�џ�d�+�����q,b1b�/[�����l����.R奡�f��=7�p��=�-[6{I��.Y�JP'~
���x5e5T
=(Q��@���ɡ�6Ct Rdk���KV!Ȉ��a�M�P� A�?s7H�o�>4QMk����ۯ�
��z��}������W.�u`?:y<uǡ^�Fj[#���s�����N�~�Rk�%I+vj ���5R���Q+�7v��v��I�ֆc����Y���i���C�LgϾXбq	�a��2� ��|꾰�'�ש��e8��ӧ�XJ&^�X�{��UV	3��k<Z}�5�>�|>�\�/e��q��Yy�Aq��jJ��h�S�.�*��ܵŸ�.�V{�D*��K�����uu�˥^=N�����m"��G!I�"�7���(�<�������W��Z`9.�uh=S0��'.9��?x&���������0���w��>���n���s��:u�4��6%#;
���2�q��z�=��A�sv��t�x���72����ę�ߪ�e�zg��ᬹa�ZxT�����+f���Ļw���LU'Q���#m������`�)0�CVMtx�H7�u�EJܽo/S�V0w<F}��݃��Qj}]߇�4�~���2W����!;���``ɓv��6.�%�(�&c�.o9��x��m���56{���L����Y�~�Z�dy��'NgS�L���~�oN|���֟�<�Չ\ѳ����X	��5[�c��������Q$?�@u���qq^�z�aҙ��x�WY�x���!a^�Pov�r�B7����x	��h�"`�=��e��޷�7mԈ���,",��xM� A��&�3���'q�H�\��D�jhi��	i𚒪� @�ּ��q6S��HgM�	H�܇�_%5�<�%�2
lt���(�����Ҁ�z 3�\�D�����8��_��IG����w�����;��9�בQi�`l�[��Ԏ���
�՛���`6y�&7��5��mH'���T���.���5)�C�	�tHN��p��v㝷���Kl��dڵ~���6�.k9%��$a��>b��!�ab��U�������o'�mٹ��H�2{�Ojl}��dD6��EF�b,_e{�P���AN^A_����qf�"���*St�C%"����y1�Vө���V\�nW�|�=�(��� ſG=:��_s���gޫ�1bL;D��U��������W���z[��7e�n9��;_�>N��cʰ=���iqf�I����,�{�'B^6ˮ���fj�)]��GC�	ʡ��IU�!j��!2bdA#ч+�� �^�� �Y�YE�m\[�@���uE���}f0��vDD��B1t?b�+�	�Inf^��a�x����t�z1d�rb�g�|��� ���L�Z㰂��Ry9d�7\�-�`B=�2�T�Y�G+c^���b��ХZF�'K5_A�<ȏ�%|� N�{���}6ؽbH�#_
\�i�ܴ��de�	ଵ��9Q]!��˧f�AF�k伆ȑ�\�}N'"�ŋक़���s킰ޑ�H��Fg.�Iİ{♈���g�k�g*��#W���Ү�:h�p&���<�"8Տ�w��)W������C�A�(���m-���~�� �x��g!�]L�3>�����	:9_�)�CF�R���=���yǧ=�W0>n����~�-Z��3���i/ޛ��� 6�����6x�;���xu�����gz��^��uG*�]W�Bc*GCV�rF �أ��m����;�2`�x1��N���������t!�@�i0hQ|y���w'��ٿ��X��ɡ��w����Mu��:�'H0�� QC���d2�W�BՎa�{ BY&�Q2���lL���khR�S�غl�4�ArqNٴ�̞�c����6����g~�o���+�'��Eo5Y���Pw0�N���/��॑��g#�x�d������F�i���hvq(7�В�������O�Z����ؖ�Y�H�/�k��s�s�)T�.+8n���9���D-uݒg�XKk[�w:i�ys�a��R`���~?��~�6i��;w��ˍA}"v��+�NQHҌjz�x﾿�^{�����0MK��8 I�*�p�N�!Ңw�hsMBH$���2�����=��Y��>x�u���%6v�&t�0���w~O�*0�U���{и�孶���.�&�R9�9}�wB~f�g�'��;���c5τu/����t2[\��R"<"a��:TG�Io� �=�G�<������
q-��DU�e!�ap��YN`�K,�O}����!�SK��S:�i��cO��C�RU+V�$�!x� �HW��v����F��k x�\��Uv*8V���]M�K��p��G�V���>u�8(k5�q�3P]�F@<�Yg@��z�{���l��{�\���XK�B# ��b/.)c�w����ۿ�(�T�$@쨩�}�Ѯ�<�n���܂�$�Ti~i?��n�G��]I��v����zD�Y�t>�nժ�����^ ���=����/�~��k��kPW܌C?��B�u��=�N�u���A:�:���C=�J׫�����%��}�#5�Re?��@.(�4&��.EF���V���/��RjR��N�XeOb"t��RD�K<��&�����ι}��i��c���Wy�
�L�{[g򼶎$�1�xd ��G
g,129�lVZo�J*� �p�F�W� ��=��d"a��P�brs�?<H����k&��qX�
i��n����]���J�0���l��b4�#���@B*�h6�A��5�Z�K3��U��t�{g�˖N����c�&���_K��С��N^�$́W[�H5q��;��5۟���$D��y	���՞���u��
rW�Z����(Jr(��m��Uvd�.��mA�X�꺛�� ��i1�ah�0��Շq#�KWp�U�`�'Ni/De��h(C���������S)o���ۘ�>g�X���O�qC��A��L�Z;5v��XrZ�C{���mv��ߢ�NI���ɴ;	���
X�����$�@v��3Βf�Tt���p�����W��uQ�VS�ģకkl<�8�#}h_
&�QS���dD!�IS[-u8Y9� 꿠��?���y�[�w��/3E}���uNr�̃XX�m����.����+?X|?��(�#��l�i�;p�9��ZZ7�[
����ח>?�b���+As>����SfK��S�����Y�Tׯ^�E$O���.��c\[�EoM�O��r׉� ���l4� *����	_o��	^ݱ��ԓ�B(��甕w�/5��V�\�[=�:���� ��6�cV�B�Q�@I��{A}�Sr��>JL��/��.-պ�\�6�>��o|9��DeO�Q�{饗h#,�}���#3����p,�}���w�-��Fb����_�}(p7]5�>c�����S����`{v��=;�����{8�L+�^3y�G���YR��jDT'���������FlgY{x���?��'��
�Mx���͵�{#�a������$㓓�L�����[�p2��c��>U>dhG��c���в�I8�"ĥR7�B�>�ٰ�D�ʀ�ڧ�O��狋��M�uhQ����
a�&C>j�7֜l�G~�����uHt��T��񏊎u����\�%-!H *Ƒ{��-�Z��d���N��V�Zo�0�I��)��G���/X�/w��èG���s��<�XHC~�Ҕ��z�� H;vX�Jub��f?x��3|���кC��M�#���C�}+��e�[?�I�-m�2���w��)�� C-�� �&'O�0ػ���@w��v�*e�|*�����n�����_{� �0�yI��:���՚�w)�){W��A�\10�]��6����t�ڗ?�A�ܛ���HI��s��c>���a�6�P��f,�:�;5$��cp0��~�G̚�H����Χ�	�C�W�7�g������wfI���w��Z���R:4�lt
S�s33;W�p�7�T�UMM�럇�(
����>Ck�e]he9�TD�좎+��s�P���R2�ϻ�IhO
�$��8��b��J��--.F4��Q-����|	��G��ȹ�AT,�?��L/����NKE� ~.�$~��7	���&.��-P2�%W+q1)�Cp A'���QCV���ǌ��I:��mi�ş���8_�'��\��]��GC��ɾ�k��3"��zE�<Y{�}��{^L���/�8�]�~9h�'��p;��Z��"� s�ܡ~w�9'�D��0|b�M(�����v���$<z���Xt�<�9|���i��Jy;��p݉a(�y��P��R\���g�w�vL��σș� ��3��]��O:좳��_��g�Я�����k�h��ű#G
Tg�W�p��!8Q�$�����k�F5������J�R�TK�&�N�H���pF�6���v��5�����z���b0F� {6�a��i8��Rv�G-/�u�۱s�]FKI!��z�T���8���6�A.Gdd��h%O��;���^�$8�~���`�f�����p$y��=/r�`/��gx���|���a�0x� ��nWTs����P�3q�3j�"+Z����`�Eضw�-8�]|�lE�����l�u®���a�!�p��dx"ش`�.��*�ѥ
%�,�E���y�H�f�z;�����/P/q��
��Iq+��C0,_������/��7 ǣ��,7�.a��3�<e�<�
C)��aY�Hb"�Q..�h�;AV���͇}]VHm� ���$ο�����vy�HN��T���9<�P�Hu�3�rٗw�1���d�(B`��X������fAL�F!���&���jr&{�g�YN�zҁZA��z@J����T���d���d�Z%�)'�ƺ�;w��7w&�(��W;�k��c�x�B�ػ�w/��0��w�Pפﭶu�7���0��b������^\R�AWb?�l����2^9���rz�����8v��\�fw������RE�>���3�y A� H����v�%�o�oβ�^}`��{~�bFb�����Yϔ��v��Bn,�/]{Mj���c��xlK�^�7����LW߻��Oz�^g��.�s�9���hg1g��e�l�y��%^i��ȥ�'�I�3�q�!QI�D��8�U���@:�#��� 	 w3jY�W?��y��»�^��J������=u�C;��8��{�F�( ��=o�\�x�o����O�GX��d�~��޵w��-[��]}�@��Pe��|N/FEy�Wģu����ـ�og�s&��t"I�#���� jLD�Y=!b~�I��r��N�V6��;���HWN=��E��Ќ��PO*.*p��Eݴ�7�>����F��������8)Q�鍞\�S��@��ce�I�;��L��|*#W��A?pY��R�h'M�r�y��*�Aokm8�hWi�����P���
�C�����B(L1����^� �V�^mv~d�;Ŧ�dr���L��'�8#I� �Q�!!LPs:��5��:4��\�h�M�1�4�`c�ӛa��ms�O����BС&�}��9	�&�z����7�ۿ�+�x�#�b0���gJ���'��y�!�y�2T'�Uk��o�*B��I�D�1�<���S�Gܳ���8�S����s��� �!�=v���RS8�Jճz�a-�&�D��W�RT�Uv������������+[�x�D���(�۫�2��eS��w�H�Nhdh��[C���~�anw:�7������]/��6^]�K��99�}�	�=�҉p��^���3���#�V|�z��{"�-�����\{T�k������PÕF���g��r�.lD0X�Pʰ��4itUhGQ ڵ@CxՌE$��%�����Z����6j�)3?t�=��3v��04e��m���c�L�Чe��?�`�K/����}�];��sI&��8�u�׬^��2������E��r`�^ǒh�&�i����
9��C�w2�z�8�?�kX��C�/�� ݻ�:o����3*rd'g(�^Ezv��I��+\�_�,>Ft?Պ�~�XLt�\h89�O�;�/j���W�g���;�jӪ���GM�P
k8�N)���2��N�e�2��F8�4p+�I��h�����M����GU�����55���Ҩ.�,<�8��"�����0{�3�\�\)�	&�=���J�&�ؗ���{��>5��E	v������&��PǍI0�+�EN��'�u���2�a�Y�fx{�^�Ȯ�v�q�kk�߻����DB�͛}����[�~< ?j��z�ϋԅ�DK��f��1w�V3�Q�L/^��.[:�v���e�.C��]�t��awu��Zk��;j�r����sëQ��6�ױ�_x�6�E���Ҋ3�#��>v���%S�N�n׶=6㫖A�k>-^��>x��}�֖/_�l����^|���]�d����J���L"'!���&�0hD��7�@�_�
�G��������N f�hY��W�6�;�ѻ��P�2�����1l)^F8��4�#�����´ng���Eg���^�Z���*�.[���H: ❺B@O�����9�.�}��z�=��8z����ȿ���S�KYn�ktk�N�l��]\� ���K�[�=N���8o��X��v�&��G0�� 8��C9$�ȃp
�'���J�`����E�g��Lq�� 5���P68~��g�s�6�U�'!V:�-�I�O ��|��P��Śa���W+<������+�3��,A{�g�
�u�9t`?2�c�����Oz�{4BJ	�}�1���k	�:!�1s��JN	�0{#���e+l7���}1�\U���^�}(�w��$5u"�
_��cĈJP��td��҄^�&I��@����!��}�w�R"�`"*$���He�}A�x�w�3�{���_�S���TCO�s`�#9�y=Y����@��
��Խ�ރ8B�C�e0��q�ꯎL��(yr^���n4�y�cƌ�����V+��B����c����h0`:d2<��S��ȳ��󘟬9��?�C(�4uT�Y�e��ng��:������=� bT�==�ll���>���'��o�nk>xB�[D��2��31�3I����C4���1	_��*�$Y!���]�����v�tK�)���R�}��'�W��ʒ,��SwXRi����+�m�JKo�w�`�jfj���QF�}�rt�O+�&�e�f#��>���|�}��S��+;-�\�[F�"���7���{����X�f�'�l��*���v��O٪e�-/-����%������#�̚*���*�N�s,q�6�299C��_׎U�"�1r�q]7��q�g�Nx��O�ܗGX@���\mb���l��Ɍ�-�F����|@o�QQo�����b�Ѣ%K��~cN)��ϥG��Q�WAO{�0oSS��L�l�z�����h}�ѧh�+��6����op���`���.���g&lcFz"�׹��L�½�(����N*�Ԥ��Ovр�(X�A�J��.B��5��
�a	t}�#�:�^�a�|I,F�[mvY�qp��]�7�!�Jc}�@�ԑ!g=�.��W~lk֬�/}�K�G��<��="�L��@`;�#-�.�������;���wi�_~��NT�-�(��X���0,����p�U�r�^�C�B�?n>�粧��?/�	��`�3�z��>!Ӎ�$�	�x��k�g�|�x��_x-�#2�@	0|?�E�#0�W�����3�O�?v��]�VZ��VWG�ނ��R�+Ƅ���h?�tֵ ��ꍝB/42����qz��ѫ&x��е7��L]@8,b���1c��=
C�v��f����G��oj�o���Z̼%�7�=���ߏ��Ye���K���e�Ə�C⡊�^L��h��,j��zߣ���	�°<�3c��(J�z2�K0~��)����Q?W�
DAr���a<&���M]U�1WJ�l0���qz�/f(�E͵=U#m��/�&�]x����@���
�5M�bW[S�+g���>m�m�Z������ǟ�e�¾��VA���}��CZ��F���7�y��6�� ���8��2$QZ>�q��P�[`����}����\NM>NC������%G�8�B�yid�$*�ຒx�q�X��P�
����Q"�g0�޽�r����Z��3���щ3�H�62�\��3P\k�O�y���9�0y>Aو�|���(�ߠ	�,�6�${W���A����.���}�����fO�j�ϙ��U{�@:��)(]��b��=�������&�ޠ{.�^��9N���
q��
�[{)�Þ�E���uJ̨}=>f"}+1�?�����(=/#�`J���`9Z�h��#\�fmY�}Ʒ�(荂���^[��5���᥋���>��Ws�U�l���s���ߎ���� n����Ι+�o@���K/C f�^}�pj+�y͜9�ϲR�+�@��O};�	mY�,��}q�W����$]I��� J$�;��oe('�C/"�.���P/�� I?ZI����ϩ��CxV�Pxp�=c�x��DA��[fn�<i¦�=�_�O��f�>f���;vm}���cc��"��ldwr���	fw%7�Tb�h��f�F@����ʶ�{�Y�T����C�v�ڀ�4�=#!��?�A�)v��7�j*a3c$��,m�RZA��_VJ��ũ�lv �.#2���L�����%��92�+��r��m��7��e
Tv*�q���i���������=�:�.�t�-�LD}���o�)�Ý�����ukA��}Q�O����u���O�y�v1�b���a�o��|��`�话⹞��r쪣J?@ل��8zo�� Vn�9�pۭ�����U�\�Bމ�F��	��5��\�h�w8�p��`��j>��jY�.��S���~�6�[o>��M�Pe�d�8R���l�B�R�C���3�}r@<TRP����d�U�2����I���[V�N�����$����G�aM��8�=V��Qu��1a�2xՊۻ��/��O���ӡ�>���<�(gIcj��(������Z�L�[����������O���\��/PAb+su���9�A�q)��y���琕d#��<��.�l ��cZ���T	��x)b�)v�31S����|��W�	�ʖ�7`w��D�Z1GZJ�U�킸*�Y�\蝟s9s^%� ]{ѧ��ITA��QҰ�?��x�����~�q�9c�-!Q`�G!�2�� s�����[9fcA�4�Q��$۬�V��ی31�?�Q�$6f��u�/i݆��.i����ÌuV@0�Q�q��o��t�= �v�:)�QK��;~��Hb	�ߟπ�h}4�A#������\������ÆV|�AS�~�m�G�����rGU+�������զ�ʭb�D��ѕ&��,f�Wv��fo��&5^$\�Ye.$u>�Q�Q���iˁ)#�`��U���M:WiN�������}�f��f���7��1��1m"(�8�>HjiT��6}Ya��~�1�k9�?�K�D8�7܇v����+q���a�6�����9�Y6�rD�U�⠆P��nL�4��uuA\k�M��kC����!TmCc=�b��i��tB2���P9b�΀���.I�익�����zk��UKf�e�.�e�m��z'z�l�Y��g��K����L�5�:~2����`U#�1=�:Dƛ�H��J�Ū�޶�ջ:>���2F���h`�[Nf>
~��;<�1�j�S'���{��_��f�c���G����zz�!+uw4yM~$�C��&{b�J����-N�Ս�L�@��m����
��$���h}]6&�W\Kt���O��� �|%������ú�ދ`x����د�zo�7� K$-wd�o!����x�~x��8��J?\vz��u���a���z^�P�)��?��魝:ڋ�\F6������y�vGQD���[��RF�#�\������"6r�o8�)Z�������v≈{��Lw�˽�깷Zɹ�S�z!]��M$� ���߄=N��F�"8Yr1���Q��ۑc�8F�u�s7ڱ�F�pMP��ә�3:����}#��Shߋ�᭱�����>��������O��fɉ'r`�V�F`�6{��g��tį�/7�l�g�V��_��[����~B�`���5�����idV �5�\0��ߞ}HŎ$�'8P�,�-Қg�q�F@ߴ�T)�I�RHh� �}/BA�?#/5���h%|�v�|A���)�aT ��?E
��l"���Wo�=cǌ��3�����or�D��6m���}�˃�f&��7!q!�D��@\C�[!���a:�R
��yJ��U��^O���M+G�i,i��:��o�%Ů�L���Ԙ ��m��g����}���a��!c`+�Z�� l��6Eɺ�<�0�2ҳ|d� a}:aɏ�NJh�F�z��*5r����u�ھ���(����qh�/���o����E�[C�%*�=�A�M5�&X��P��>�p���:�Y����hB#���r�?����_�!Li���>m��C�����mݧ���\w���T������Aa�I��Ȝ.dm5D�c1�U�Ec�����5җLj]":��,rS!-7�6e�
<D��pM��?�)��b�<���m�YWS��5�� 0Z�N5� ���x����ߏ�2�	�-��A��z���`�"������yv{�[;ǭo���}��ٔ��@�q��������g�A[`䫧���!nQ�
)R�Y 3�ԏk�{N�y+�L�`�*a����[N
�
L��(.���u="39��A�g�q�pF�[)43~3��0�#��>�%�Ū�N�<�w�l=�g���ӥh�"��Fy"� v��*x"���� uj�/<�ǰ��U
���5����!Ba��i-u.��V
�N�^e�w�]iO>���y�g}X�~�ۻN��M����Ԭ�!�2u��B;4X"�~~ȕW^I������� ���o�k=r  @߿��ە��v�u׺l��ݷk�s�%�������Р���v|�� �� q3���؇Ζ��]���/�����$:��D�L��,��A�g?�������|
ׯ_�lsS��iln�ep}CcdK�@v����#�L�f ]d18iGo۹׎l�P�D;� �S�`��}����q�n�}&�Sz}�>¡l�T��r79v�< XQ��[_e�����y�lƔ���+9������0_��7�����WͿE�C��I4�%
$'��]c�DDDr��d��\^18����6o�\V�e"RAv���Gn���8R@$A�r������D�]LPJ$����Ay��T�ʱ��Y�tp�o�ڿ�>q��v�m�����k����˖0�}��d�R��E*�5��Oo!䵻z�7�Renr��e�.R�c3������6�9��^�0	�p]RAÒ���X��?��"_���v=S�Əlu�GP΢�J�\����gᔆ�~����N�5aN�B�2eFq�%غPo0{X� E�^��>~�τ<�u�K=؊?�����o�jϼ��*�X�{�1�0��p�'���S�����4T�P����κV9V>YP����`�9�U�j�	�K�^3PL�
��?m�lJ����:�> ��$[gy�!)	~��G|���#?8)�����ǧdM+ Y��|D�E�
�T�R][�i�Kcd�:y��p"�)���TD]��P�Z��*Ѽ��s�j�˿��9�N|��S�L�p������>�[n�ѩ2[;]�J�\z9%�}�e���_�+^�Ќm׮����w��h�q�~���=x��-{�ο`!cp�8��3��+/W�n����qp_k�^�bx h¿B' l�O]Sr��;�>�r�r��ϺRS����s���ٯ��\��ɡ�jlL_�a��8Ꙓ�����[�QKLD��T���f������Ç�`�D�SD�����}�*cA���J��ͪ�T�\ CŬd��F�K�U���)��}P�g	r&������ߵMn���y�]p�v׭W�k������:]I.2�2ZB���Jӑ�`Oϖ�We��׻C�v9(#���QCk`&�-���F2\����'�ēO�o�Ә�Xu�d+
�IqV�����D'�Y��2~>C;�iA�]����{�w��P�>��\t�U|�.{�U��=g� N3���]i�@����Ϲ�;k�9�]>�g,�\���	��=�I� k�W��4�Rצ�j'�J�ѐ�Va*s������#g;~�t{��g��M�v�U����=MMp0
�_�!L&��J�2�U����%q&���YD���VX�`c�"�����=1H�IL��R) 6��^x�α�!�,�MC�"���`V��b��2U{:�L����md�@&B��ºv"�������C�Pe�T~��/R���_��x�\ �K�^`�_B;ϸ� @�M��w�i
3�   IDAT'��l�jd'p�wt���ha�o������ة�	�$�(g@�u1�-i,lݺ�1�3���B'|҄
��!b�g��_�?X�0����l��m����il_���L�f���"С�9�0�L3Ư��z����mH�j�� ̳��MSsw�D?��i
�Q9�׭1¥�'A�IK��з��P�,}߾}��~K���,�RD���_�Ġ(|�t��KBn󢑩.��������[.������$�;g͜��N�u����������>���y@����3!}]S$������ FhB���n�y����jD���]��<FQ��F�8�:�Q`��qK�Y�.�G ����1$��H�1��R����G���,E��������ޓ���~�nڴ�>��?���6kNA�zmS#X���Q6���)	�e7\\��5�w�P��Y`�l�2�;�찷��l�h3���O?��U�w��-�<�P��Ny�h�e��N4��{"y)v.�\TG�� �
��.�Lc������Wھ��q�7؍L�[�H�e/�h�З^�t1j]��z�y5�K���¦O���:;�����3g3�15��D����&�@
i�:���N��s����G�4͕�KtF5��\�o��o�kϽi_���vɢ)̟G��p50p}'�m�1Y�Hs�%���N��@�g�{�!�3�#�2=�:�F<4$f��*@���[�Yܦ�AT��A�� �:e �����Zr��s;����bŇ�`���� �i��B���d���O�u찡���$�#[�>bל�h�����,��^rB��ѳ�����P-����!���_��l��3r�Z3����^g��r� �SK֟A�$�z���;������)袮/-}�ێ�u��W 9H�(��P+�_�������X���̪�ei���;�
�E0L�'�}`�ԕQ�i�"��|���*Z^���>|D��|����z��KO����ι3��\54B�X��0��S���V"�y�0b��%�{h����{0�C���r[ ����2�@ !�*�	�^9�я�&��n��f�#�3��^PXp��)�>���?�������d5���T�զUk�ؚ��!��B�fu#뛽��A��\�-��+lƴ4;	���C�<xZ���_4R08���F]�g�Hv��b�b�f!��=��|�����l$�o z�j˰��Yn�A�21�#��bR�Zgd\���9[X����p2V�T݈+:��d��� S]����N�5۶��V_WK��0�6�l$|ᅽp��� ��T�ǁ�0�{�����U&f��'G�ӷT_����䕳m�Ⱦ�o2�6�6䶛�A���y�Ο�MEX&��L�C�t��{�dd|��G��~m��݅J�T�G�%�/�Dg�;o��P�gv��qB��lzo9����:�^��'.�ac��#߽�>zg�}�37P���vHH�tA���ɨf�ۯ��<�<�:�ikk7hx�F]y�5�r��*�&�����|�ݿ��D�޿/�_��w���{�))/�۾�i�����Y�b\B�$��������]�����4n����:�;�A�B�����=��̓�mҹ���h���wu��+`���Hz��m�7=8��''�Yw�}y��00PE�M[�z�9�w�ə+��U����v��+�]������΅�7�l�E��^�k���U�	����G�^Sjϡ<"�=���9
<��+��)����q�t	F���������&�X�+ߴi�-]�L�I�QG��$�U�/�I�KG"������3��xP%+J<��OA�~����S�竼�v�"_/w�����0�}��!��[5�:aÜ���8��)o|\��'�ث���`�N�+Fk��#>RdP�ѻki�i��[S��;�"���4�Q�À��y[�9sfؤ	�\��f��+�*Cu�?��%���sh�$2�YS[���j�#G��n=�#[���q�J�ߋ]~��=��-���U+����� �i�v���"���2N��kYd��8L�d�@�����¥��.�Hͭ�]�b[�~\em�M/�Ղ�N�z<`$q ̙�#����_� C���J0&�W�c��C�Mjc�8�&
�?~{�=~�Cփ������~���f����䙬���KZ���蔋#��a{��A� �}�UȠt}��u��d�P�r�tp8Z߭����{UOSp
m��Z�������t�T���� ѭ��hK�ůt H�����~!&Yp(�3�o�4��cIb�ݛg�a<i"�|]$ơ��w|a��:{��1�IL����l�v����g�|��_Ǝ�?��߱�ϝc8�NZ����_�k:��GN��&ڔUtpL!�Գ�l9��x��=�s*gDT`������jiL&��%����tx}W�re�����}M{5����ʙJ�p�򡜷TϺ���	�&�c� _ר���#;+g�.�$`�������$w�K�K�3�GV���"G/������;m,Zﭚ��Ek� D�.q�B|ͪ�K0J���G��ݷ?���^��L�.Nl����Mr���p��3:t�3�s�������#W7m����A�D<�$�|	���ńg���$�C�q�����Ǚ�=NZ�L�c�a Sҳcu�|`��Qמu�?i���|-15�W�����1��Zp��cE�n]�icCr	�Zx0�"jee�c�icc�Rݦ�Ȅ*L���Pi��P	9ۣ�'�>?A}L�^��d��'�1���N(�r)D�f��Lk����<�m�V}� �-���f���$?v�(ˣ��՝f[p0]���u�$�A��g�N����L� 99Y�v�����=���l�����l�7l�&E��UϞ�]��$G�Y���j��ೈ��Ia���5��XM��@��[�X��`Y Bwb�#�@}V����ꏬM�	r,�ik5/��;�Z�:Q�[C�.�lgج�S	Ph�#CΆ��=c�NͶ�o��|z4��f�#�8I��R&��/}���~Ϟx�Y���X����fvG+g��/�Z��֮�h�J��"�����t�]
R�a��?���YQz���kw�����a�9�1�G�� �O�P=���jo풟p��M�-$�^�$�H��� !82ς�q��\xF/��=;ԩ]��]�:����L��g `��܀F�K���4�G��J8]~�j�Ti�@3)#T|͍�3�}Pi�3�{���*��v�U{�+tKcF������R�T��3(���ٺ�ߓ���Y�Sz�l�ni�0����z���'���{T�G��A-i�s?:��H	&v�_�� ���Cg�k_+6y�Ć���>\I���j�Q���R*Y��/_�$�c�=i��~݋�/���x�E���&�@yjl��U>\e��INZ�ǹ��6RWK���Id�5�T�ʥ ��7՝p���h��̫�(.��iɻ�k�ȉ	�i��o+1ѿ��ً��^��E�n�#E��i���d'�
��������_e������� w�DEy��o4��>��>{3�w��Vj�N�V/(΅�؝��5�LK�w�e������%8���1�8e��h��1n�p+�#�4��^/å��a@�}� ]�\�4�%�)x\D�B^k
sǭA�B0r��8v��U�V(4AN�&3%"�õ2�"8	*vL�0u�|��S4�gQ�v�Tk����ʻ��w���-3��#�54�{q��Z�=���-d�2
b)+	�~�?VF��Ք�T���y^�*��4�LBư�@E��'Q�k�X�򚬫Z�	�S�����J����#Բז�`n�:��ҫm���FO�wW�a������2��E]75�lI�yg�-Z0�3�>,co��Rq@�hCk��Ńa}�V��x����^Lrcab������O!ےs�&ؓH�'���s�����W^zپ���l1e�y�̴�UsA[��Q�T9�H�2%%Eh���QaЈրŕ�Sir+ r��'=	��q�zFR�k��X8�{}#~�C���ݙȨ�K{I�� �sR�<z��@w�u(-$�*�
Y��¼���+�<�;����Ճ���8
���=�N��O��O)��G��{L��NIp���5���QMG�}���w���#������P����y�A:�㑣�	����wR^��/�g����hMT+���YJ3 �KCah]�-���}���m�=��Ӗ�������,w�1;�R&��ƌd�#�[=�z���"Mؤ����ҫ�E����6��5��G�m3\��G�Y9��6~W,[7n��h/�@^�2}���:U���s�މn>g��@r0�9�/i�k9u_�g� �$���I��;z4@I��gy �cuGm�r���ٵB�;y�M�6+
B�$i��F��L�ݹs�|�������� �x՘��pvf��h�N,�jHȢo[�Z�e�ZiǨ�1ᱚ����\G���Z�y|�4hqI���M>5���#�HA;X�MBm9���Є:4G��6"��cL�hT�L5�j�v~���k�&a��뜆qTF0�S�����. �>�zS����L�\Xak�[k��Ц� �k&�C��A(�����v�X�=@�z���V{��oTc�ҁ\��o!�(�O�[~y	
:);�=��`�Lc6�tZj���_`�pZzp�\�kWW�`�t��E!�h���[1t��D��aۺ�;wT�}��+-}�D��/����`��* ?k]�,EF8��-pD��r�9,�/�U��'�d{��
���P�j��=�����L��|�[v��>��	�{���fW�����L�^duW�Z�����%���m��d{� 'e��FRP��$D	��eT�vh^W//Z��$֗c\\��̃C�(ۍk�1ĭ���1�3ƕ¼&�B�C�8��*�p� ���q�0�24��>�D�he�/G��K!��+��P����y�Sr����B����Ro���s���(�^>�3%Y��<79��>�^�4!er��>]��߷��!�p)��y�ZC�^� ;	2���|�F�m7�v��Hun�۹�ؚἯJ5�s�[\>qTK�O����^�,dy/\�r�Ql�ʆ��Ł�D-N��ʋ33	_�������Y��y�p��Pd��x5a+e��jBTWx�g������b�ăM�U�$M��=Uc!�eg���)6��V*d�M�7`_fD�<���8�Q]A^�ug��y~���z�*�N���wo?~�������b���\Mk�Cl2���e8008ٲe�$����� �iC4"�
QsK��;�.#�YKz�G�֒}�oN]�Q���5���d�FV�EY_S��\J�-IQ���/���.rDړ>�z7��;�T�n
�F]��d���0\[v#x2Ē
JmՎ#��������5��s�b�AD7����A��#�T�3<�_-?C�jp��aF��z�"G�@F@��j�zU��T�=uz�%�q�q�m� �ry���Ȝ<F:�Χ����hړ2�S@�o,[i�m���]eK.��cb��Xf;?����V6t�u:�:��uI���&�?���x$���l;�Z]+�^)�d�@��F�p��Kx��]���yh��x�щ�N�g�(H2X�x��iO����;����!��M���'���#X������,��|��m�	�q�'N��{���;9���r�AF� K</]�i�h�g����LP���8�ߡ�~_*xܓ�(#�{�c���OW�jmF�>J�=���$铋��SV]��O+K  �$��<z}�U����"eۊ;��~U�Y�L�r��~m�G�_>ڵ�O��E�&
Fh�Sp� Ճ'����"`��8T��]*%�d��-[���L���I}���P�kފ^R����tq ����	�/���{����&�yP1b���Rb�3ǥ�b�0M��d�
ڦM���q��hohU���$a*�r�'kN���·X�~-��'��Z1o�w���b�%.WgFχﵢEp��Q�m�)l��N�;�ŧq���Q�+��`��M|ӵ����fĆ֞uggW q�Mz�B�&T=;a��y-�����*-F�q8I�8$ ��A��v�Hf��.I�}{������DXj�{����.�[D��meLF*\�/�U��O&�Q[M���J<EKp���2ow�b֪�,�OI�!��Θ�|Ԧ4�M:�:�R��GԂ�FA��
L����X6����k�S8�@��6���1�Ùƽ�qo���Q%��8�P��'xs�0i�SL��|�>�,����K �҃:	Mն�@:����rP' �=�T�)IY���^GvU1&O��1�(N�u�d���-��>n��}��Ͱ��ɲG���`¯y{�:u�Is���/gRRP�R�&��9d9�=d�745� G�����d�"��(��uHpD�;� �I_���r-�f=� 4�!/�|	}�?���^6��>�_:%H����7521���Ai��3�O-��=�׮���
�j�"�鉳X�쥲�W��3���;?-;���;nq/"�8��������Bb�����~ �y��I�=�|�F�+d��_IT���^"�/�k�����8pP���w�F��=�3��r���"�����`�u,$��J�����cQ�ٕ��2�q������P̤4	�L���
{�7��}Ѧ��lݚ�v��v�D�b�T�m^�s-ބ����S#Q�G��{�H�8��A���p�x{%Z&����F@���kh�=J9as D��" 9~'DL��GIZ*"���5��?#�b�LD-��W�
���	H��)3�E�f%C�:4��+Wr�Rlڌ��*���<�tm`���g�y�*��{���=~���e5ͧN^�y�ovv�|!��JX��'��e���FN�!�#]��\MU�i�k#g��6Po֬�eZ��v&79�'�*��LVvv#�IZWľ֨TШC�'\ ��A.7�r� 	�֐�F.��ȥjq�>��p܋��"�۾�`g�yN�3��Lm�YԂw"i�ŀ�4 ~}�_T0�k��#&���e�n��� $�-��?��W��cH�J���y��4��?`BU��㴪�'
 6cϧ ��L�3�?e^�Lv�_FK�"�"!MD'.��zg-Y��֠jw��T,Z:��#i���w��Σ����t�J)<CƢz�{TF(-C�� ����[6�E�K�a�5�Cq9l�F`���0�=�Rx��<p�`I{փ��D���05dHC��3�A�>��+�ޓ,��^z�a�����j�����@�Q_D*N��K�>c�G"��`!�d���_�S��
]`�_�f���78���Y�TD��}ND�Қ� �@T�	���U���5���p�Ո��"&��;hV���&��'����}��8�?T2���CZ?	�� %l�!$� �!'�����kՇֻ� �l�6^҈����j���NMFD=XQ�c�>n'��Nƞ��u�;�%��5pWJl�ıv U���˟B *)d��s%GݮVR�Z�G�/�g燎2�",Q�%��%2SY5�&�d�7h[%W������ҼtOL�y�~��+X�#N ���7���)���O����9'��y�&A�j��XLv1��]#�\�.��-_n�tL�̇����#*+oŮ�<��;�+�s�����/�8w��/�~�zs
�Y#��W���J�3ȉ�K�����{Z��}�y�Z`�#�I�z{O2�>`�� �f��in�`�֤����rz@� ��>�60H,2��m6��K��ٿQ�!:լ9𚉬y��a��P'�`ϾB-�� ٧Cf��f��t����O�E?;7�ڐM�Cf�!�b�bǪ���rT���L.�������֯�*�(���=TAx{�-L�R����e�.ݞz�Y�z�:��	V��Ɩn�&��0�S�8���Z�CFF�����Z�z�Dԯ`+Y̼f��à��u��}���wV��ɣ��;��1S��G^������	�%�Rv�R�����x�0I̿�������Qg�Ӹ߀^p�V��������u���zhN��B������6x����$�l]9u	o� ��T.��8G��+*�Hr��(H�d��4�cMqm�X�ǝ�#>qF�ᡶ���u���t\O�0")R��25}[�Y]��q6�Y��C�EL*mi��*;QF�U@����?���+۹�������Ԓ%���er��)�6P�6��|�O���Hb��y=�3�ڹ� 6
����@�%Y�I.��*�����Ҧ�c����,5"Gtr�n+���l�$��i�h
Ӳ��YU�6��Wi�|��'�rih9U�u�	x��K�������T�V�1oj>��(�M%h�f����Ƕ�ۙWPƬ�:rj�M'�+1Ԟ����b�+ tM�y�V�W�[���a���p`���ڛOB}�*&5��n)�qW$� �`���+�:��u��[��[����3f̼�̚�(#�sZa>��%�����&Jm;2k28�vF�n߱ӆ�bR58�x������0_�wS��s�!��5N�m�Qk�(�O
�5V4�O�������p�P�F�J�����|uE�(v�b�1r%��^0��?�f�m�]ck7��#D�Ɉ�t4ֺ�L��������d2�ة��$�>5UK�0Ғ���5K�j0��S�i:� GU%���h�S�l;:A{��C������:פ�3WICP�g��F�#�����<�n�3���.P�0Y�(Պ��Ae�ǯ�o;7m����̖\9��Ng�<�2���]v�����`� � �Du�6�!P���� ܁=&	j�&�M�`>������,k�0}l���NuW�ĩ��JrW�\�Ԇ�+A��x�QJ��:)"$��S��.R�ڧ��t�����8�Hu�z�!��a�GaҟH�͹a�:��;Q=�ș�ǃ!�Z�1��TvN��{��Դ����o��Mx��l���L�z�EN�齅.R(DpM| DD�_!����p2�	F�=�53A�9��2����#)y�v ��
����Z術 ���CTO�=�[���X�Gy�:�[|�BkR����
�ƺe��8S��M.&H��J��3�P�
���!2��bDL���~���~)"�j�>���l���ࡽ�W�Йo�q�^\�ܜ?S��;���g�!lׁ�G�Sh3���yh]��x�C@��7F��Ғ�i��'����K}2]7�T�h�{���l�9�@U��H⺺);�df�ͼٳ�h�U����
����8t�Q�4�o߶困�oK!���$�i��� ڙ񉼍C\āȂ�J���U��q=ҝ�-(˥�%�a�,�KiJ��G�>�g=]�Ԑw�SɅ�^YJ\^'Tf%�.e;i7��P��0a��1���ً%Υ��YD>��=r��8�j3s�-:o��<�
'�=���8�B�َ!��� �H�w�S���1�R}���Ԟ�a�D�F��p�r �JW���.�70�6��"��	vb�7;�BZ�9��Y��/�ko�`(��pa�b;�`Dr�m�a��k��G����p&<�?"~)��:��A�H�SC|R�'�~�^��\q�U��������f;����̧O�y��ԧdA;x�2 e�U�[6`�q��O�xj�J�A�ꪜ��ҌH�Z9\�*�T)��9j��X����lwJ��-G��A$+uVh�|4ｩ����C
Qݪf2]-�w��
�=�\C��:9����Z����:��h�o�=��C+b(�8GC�C�	(��?&z���`�L:~_�-i�HŁb�L�z"j����!qT��{��>�!ؔ���[-�0R�6��R�S��]��?�Z�vG�Q�%��L����B���!5
���o���Qi��^Ϣ�G+pJ���>�Ћ�����=�Km�:ɜ����<�>X�j�M�w�g��V���ΐ??���s�N�;�4�AA@?/aMC<t谳�%3{��ŜU���:e��awYCY�<��W_㊄�3"{��5&�j��}��N���04:�2���f��@�m�$'�[A��U��E�X�2�i���ގ̼�ߝ9}���:��+�Ӭ�/̡��
KD}�}�ƍ�՞��˴��H��1yiR��ݍ�&��g}�@K�F�׬	'�#���,���a8q�s2��bF�b�
�n�J����8zR��Y|�0\�Q�r�*�+��긲?�:iw넴�Q��1��""fZ��3p�5ntt��`�2�`?Ş{3�����λ�:ˡo��T��29�n�<Ԇ%;�2��!����d�>e���1�"ƥc<�U�À����4.H��6��Q���CY��E=M�5k>rG\�����V��}�QT�\� ��k��Jqp�O�UٯB���&�4O�#�Rɱ�@&���������m�j�\u�\�:��^zy�8�8�.��l���>�P%�.�������z������s0�Q�,��Xb�_����2��l�WY)z$���*����0�.f�KMeYm�'t��B��V9D�{<�։�du��;��ԗ�Q6��U�w>�2�֑�f�b��� �]]p��޷�(<\��Z�yCq���^���t�Z�3z�^a������3
�8Hh�����z���3�/��:�u�ґ��8���6�Vw�
�D.̀���>�e.�>:�9̛;����\:G����g����N�
U��Ѝ�t�a�?ϯ�� ?G*ǞlЂ8�s�����v�$�B�]=��C�:jF�A�ie���:ˢ��2e��@�� �'�!SB�X�.�#�+�M�hM���ڌ�ciS%;�}Y�f�;�"B���G�5p�8����y���r*!�:� ;	�I�P
�b"^��ZgG�t�G�ߎ�[!䎀��)�Ĳ	zz[lێ}t�l�ˮ����g
�XC�c $wM�4��Ɛ����+���:�x�Q��6��ڹs���IIs����<��8du�����%��7)�Ip����C��F4�Qcg-}�v���gX���9f��W����T�V6��C��z�����~�<��@b�IW��@-��QR\�5�,�ȑC8F2:���9���
7�t�����v��C��O���J m18�ݎcx_��ZaD��Z�>&R��ꥧ�S����kP��C��d�;��������9~�&{��0���UW���D�Du`e!q=8da��f���)�S��f�^Dgυ]x�'!ǯU����LYa� ���{�'�Y`�<��/�io��ܾ~�ޖ4�,:ǫ ��Y��8��k���AgØ݇�0�� �}�뗅��8��Ĺ�C���������^����C��k��]���VDwV���Ba�@E�ZS��B��&t��T]}�l�ƥy�x�@�R�F
n�L,κ����{L�<j�bcf�=��dv����{��$B�?�5�φk!+�S�3�%	��_[�4	Ԩ^���C���f6np�����!T�^Q)�	��
�����Ӻ��x��=�T���WP\t <�Ȃ��7�`P�5��$0�����&{�5�?r�x�0G�Q��H��,�3]q�y�axsiFx�^�6BqN�,�?�F�/$,]�5Μ���2�W��6���1J��Ϙg���Ĥϣ;Fl��}!?Q��	�
uN�MoK���]��Fjr��QJ� t��6~��;n�2��;
"����F~ۘѕ��=�qv~���8t]Ҋ�N����h�;�-ͷJ�x��J;��:��r�W��o������;vh�r���0��h�x�����Cl+���\�c�m������i��������5>�ۛ��㹠0�1���z^I���'��V��ٗ>`���{�햭z03f�a8�2���D�z�¥�P��}���qL��4�Z`rj�K�v�����e۷�W�|�v5n�Io����)=��%Jj�R~Dg>+{��=�@�T�"�7�8�)��P��?�	k${Ջ�ӫ^����^y��n�n��r�,�Ȫ	��:�4�S3�!2���])��u���>?��6�哷�[���_�ŋ�n��c�5�U���i���DAK6���!��v�w��'�.��ߑ�Z����j�oC��8�0�*�ax��j��\h �yr聦�������5വ��l���O>�q@�ɄzT�t��� -��R�6��i�~��恌�+�)R��,(Q��H{�j�L��[��Ǝ�� G�A�j���j�P�4*ރ�e�B6t��m��p'x�%Kq�]>�'�ƹ:��L�����䵬Al��LoIk�<Hq]%�V�޾�A�I��Te�ɪK��r����$�S�Se.IȊ(���a>�~*�"@�fA:�����Beee)�c}�	{,�bN��J��0=�z݄&<�C{�D�_ǘ7�b,�ќ���0+a%��4��W^����z���Q���6X��ُ�+�Z�����������P���� �֖Ɔ�$�`EQ�� [/.F����A8�$6~
S�2�pع�b�*�BX��g['��G�3��!�[�$�z�9�m�6��1c�ۄ�Cp�!�$�G��E��r�:|��O��$)�ٿ��Jy ��wk��b��J�:՛ak����s?�`����ƻ�
$:�?̞��c�osfL��CNA���"��ܗ���6� �T��+*q��L�k��5���� 28%�
���v�u�45�"��3s��9¸K0m��W!v=-pQ��
������Ba"(|��Vʍ)�U�s��Q��w�w���U��u�,�E14�&N�!i�|�ú�&�̐��v���Y�h��.�&�Ǹ����5y��S�Z@����*���ڲ;�(�����]F6��ƻ�|w�4W@=�bs����C��lz��О5d�p�ko�P�� �=AʎV��GL�;�4��E
mq�<�Ɵ�,N���u�����-����Q�1�.�C4�tx�4��hhPN��K�?�[�P��N�j���a�&�ʧ\�3��-�f � 6#R��e��0�ao��v'nD�(*���g'^���U��͜1���~�L��,ңZ�:E�D6�;��y�߶ێ��gE�FZ}� ��I�(0��׶m��5�����(g2�WH��j�]/,.��	
W5n�;�Ľs��<m�c� /���{oC���ATi;�	���I� ���e#m��s�/��J�h�	{���E����$Gzx-��GƏ����3?�)���O��T�_Ԕ)S�=�܎�S����=nl�5�R8hI8Ф����O!�J�J�i;�~h�9��+)���@��ja�����ic���E�rt��-���ۮ3��ЅOơ'ɱ�	�4�P�X
��a��u'���-�`n�@!S�M��u��^s��	$Qq�ҳ��o��zժq�ͮ�e˞x�I{�����[����䖎"^&��A�+�lL�8H2m���`P�i���^j�8�'�Q�vN�</e�N��P�3��m���!�PY+mxd;i�2��e
�O�SM7�.��ˡF�.v��0���TK%1 �����|k��{!�Qho��.��G�m��Cݺ����.�c��~���4���H���6�����w����jm�{�u_
$4>UR�1�-#�(io��;������J ��X@��YhX�dh��
P��#+�#��]?��.�މ�vq����b'��D��ڎ��8{N<��f�}�sq�y��q��w�5D�y�>����9Ew�A��3J�W];��*G�����]�����,WǴ<�^w�кYOp�uU��:�zЙ���M ��if"}���d��Zڧ�P�43����Q�d���Q�b����wшxSÖ����L�R�Iq�v����J�<�&��r��|�\C
�\���?��CxU�T�RA$��m�L����9�'��Zx+&��p�1�|Y~�+����y+�}�@���J�gRh=�Tg/���>��]x�����K���<��ٷ��������V����ym@�{�1|ٮM������4 �Q����`�m�EO&�p�����}jc�f_��ZkC���>�z�mob�t��f��-���x0�� �Y~:caZ�>I�����S�v�X�p�pu2�A "d���	$��w>�]ZM�����N/l)����1D����z]=ϊ�E�Wv"u1��h��\~��������
�4��֓V�#������/<a�?XM���i,ݲ�묮�ىt=r�~��n����x�J��S۔�Ek|/���x�\�]���z�-�D~�gO�g�ъ�:^;�� �ސ$k Np��<��#̡��EI��6�TeÌ�<J`� 
w�̞K}�yv�-��=j�h��t�<2��B���|�p�&k�bD��$CCZ$���/ؾ}��+�N��ˠ1�E��N@��~/A �3�+�h�����t#ҙV̵�Ez,s}��Ѕ�\)cO��e#xS��?�0-�f<kF~���%g��Ńx��s���U{2@��L.��u�~=3� !@޿��%������N~�#B��0X�1,�b#2�yҳ�-�D�������
�*���g�\����Z�._��{��좋/A��!~DQ��p^G-�B��eϭ�ʞ���ե��F2|}]"09(��9ڶ13!�s%T,��Y z}s�zH�?X���ɏ�o\������&8���/�]�s��E�qv�5������z�?����9���ٵ}�M�tw��!�)��|��<�y��^VA����e����s���3"`cH0ph��������/^��o�]��b����-��P�wlٴ�պS�����SVչS'#	{X��28ȭd�Id����\g�W�õ�l�4Zi�q�Mv��y>��X����� >����d��ad0�q��T�4� _e?�n���wp��G8ĪS�Y��ř�0'�;�A�Zi0��		v�G$/Y/'���a$;���777�zVa�1Pյd�������_���.��.;JV^3^c4��'���܎1ԇ���U�p�3몱HVv�Ϻ�-uj)i3�����q1��A1���i3�Cj�b7K��d�1	~�x�P���D��-�l�!p*^�KW�|׶"Ρ�V#�r���S�����o��]v�B:��*����!Kme_�=EO{��i�.�>����(4��?.�Dsԗ��Sݵ��1�Ό���[���������r��x{}�%N#����[���}�ۜ)+�5���$��n 9�p1�2��+�E���~&.w��q	$��l�I]��{�'�����]'���H��w"�_]r��N�'�O��B��rH��l�jǪ!oř��<V�ЊZ Gn�H�8EX��v����:�@�
��o.G��M�5�W��`�n	��YHC��������Ì�X�Q�#�&C��J#�h�'��];�� bG�� ��q��Y��G�`3��ë���S�3����h�U���5}Q@�{(P��q�TH���R�wvM��ךvioDA��1)�;|(&�t�p��+ �h߾����/�pa~Ⱦ��վ��U��]�:�]LjK�jfGW5�֟�8q�+gl۳�<�?�
��:���'O������ܳ��@���'#�������z��F]-�������nT�v~���W����>	�P^����G�0���$ұv�x�P?+'�M�A�C-_.G%ֻ2e���qKh"M�9�)+��Q���90�j���`}���%F�A�+��8�0���[iv�؄>{�f��)���uͶ���,73���@�yi��L�p]��d�R��Q�ޫobv�o0��C�n����hg�fxƷ��)���
� 	�����ӷۚ?rt#�]M�� Ve9�s\FM���X{���8��>b7�RG���}�ۂ���ŗY�]wڏ���{�|�fM�aW]�r�-��Rk�π�xU���,Bf���D�r�H��޶�O��i9���y�Qm���wZ�=�Ń�[|9�&���	���S|
i��ҝQW�|moqcYX�@��`<�%H����t��b��S!�S���'Nĵ�8;�Y�B[b����
���l��I-o����p����ۑ�ȑ��3j�R�7���;@�NRNn����+8��X�x��)lI���A��W�0�э����0��w���g�>�"JV��|�aۿ��*��Iv钋�XG��b�J97E�߆-V�t�N[J{Vf�Md�y �i�B0lRP1y�Tߣ�w�t��մ�!��m�����=�K_�zu��v�t� �5��~��1c#�j��"��ˮ��&��'�Rn�m�[G���c����,��_:�?a~%���oW�SS_�Z{�/f�6��iZ��0<|�C_{�����kw[���>h�u��r�8 �&�!Ds��:w�:LBr���.��XW�JWլ_��X��=�(U�mi��{4���X���K#>�	g���!^������ ��;Y+�]�C3��z�;B߷e�x�}̿�S&�P���� �l{��R+*+��S�l$����Y�1�4gq���{9�PT�eХ���G���=ѐ�0��Yi]�2�m��mv� �"z�;y-����\~
9�m����oܲ�kU�v�����5j8E�ځ�#��٤c$;�d���OP~������|�@����n�+/�g���K��w���]u͕6f*5�"��"20�����n�f����<h!*)$��&1�^u�}�І��P&*E;ݷ����N>�-m~���p��hVzZĊ��ѷ���shW hP7𺏳��!�S=Jf�[m`�V;?A.(8e�j�J�<���{	����Ͻ��}���O��g����r�q�BL��|������3%��"��$��]V�:��K��; _��.D���މ�"u�CC-g)��N��5`Eg͵��J����W�����M�dњ;/(��^�� O\�����މ_�-pu�W2�ƈ�$� �N��l4���d�G�&pϴ+.���#?������<r��K�\��sf[	�/�xwX_-���`�{�R#q��9��H�k9ٵma��!�г���3����'�#��w��k�@��^Lϟ�W�Lb��8�=RXuv��h����ƛ�͐��~�׽o����?=lXš�^��
�<W�Wơ� �O���[��ˀ����*�,�v��VuTEA��>T��ˠ�YCK�5~��ƩH�@.�M����ӭ�mj��a��1~.-J�v23����ءc�sOQo�wv�
�N#�����{�}���4 �|�?N��� ���G	�W�LM�Eҟ�{,���Hi������1�Aģ����Mj^S�X|y��q�Ў30]K?4�ja�G�CY�H����ԭ��������օ��k~�Md�Tt ���P7ɤ&���h�b�Sh�QK���zM����"�W�cXCV�HH��7����{�m>p��W\bþx����F��������.�,����a0����/��k+&9T���Zf��	���H��-mt!i�]��ݪ���&����2�l����O"��� a�`@rb��k��1���ՠM�s! T�Bh\Cܝ�c��Cv����Ƥ̐����iMu����ޕӊ~�oM�@�����~���,=�@���ܯWLs�2J�̙��8���u����^\�pe�s��v�^_��Ⱦ��b�c%�?����[�QL�y_��$(Z������~���\�V �tᶮ[�g��$�.��JX�{RR�gJ�A����^��<�>���G�P�{���_^	A����H���a�\���wJ���J:����x҉�T�f�(t�y�GÆ� Ð x0�*�-�5,Y��*=�~V��g�ǮD0F-��<�n�˥$?:jt�]��%-?OC~��ή�V�WʡǏdҤI?:v������=���5����\�Yw �%3B����f$���4Z�L�M�62�k,r����]�g�@Yl�Ɖf*���vJ>#���l�U��\Ϻd��ཞ)��gU�z��#ߎ!��V����K�5���  ×|��C�>w:z��e�xJ�&���T��޿�ڠ�Dͣ���1���a�F^F�3g�Y���*���S&[=��;+>��P��-r��	�(c���H�Q���'NA6�z�����	L�s�#��B�y�����mY̅Wf����{������˙7m�=������W\h3f��GK��՟9AA��(]��א��)���G�:rr��cǥ9>g�L�漟)&?gwR�!S�`-5��r��o_���"���߸��b���*'-���[�������vK�4j�C��q��(TぇĒX!
���(��j�!�T6^1��B'�mΆ��`Jh�K�-�q�P��ʶ��zv�^տD�;�����;}��Ϋ�$�����x��H���y��u�`%�W�/�(8��u&Qcn�a�X�e�icȚ�GV�^�a(�)ە|��ݻ���؜�����:Xk�A��u����z�3�h*lؼ��t� ���r/#�d���`[���@i5D�0���Lx�B��m�cFW�&ҳ_\�����S-?%�[Mf�:�Tym��Ŝ�Ŵ�%����t���|�y�~�يg�|v��+�+��uW}l'3\�gǎo3d��>�Q'����9�����m�4N7Y�KE}��}ȚZm4��
����7���t`h���gbD������-�̮�ǁ͚�^��xի(�sw�G�[~b������L�x&�U��2��₽Q�V91�cK�n��J{���j{1z�,�#���YM�!�;	ý�2��A�C�KSİ��{CO����O'[O��fg�گ��M3�iS���_�ĜL��?o����Ȅ�;�H����4S���E�N$�!x[���!_�ۑ	_q,C�AD�7��:!!�K��{�����EH��������������ī�o�����&�S��LA�'��.�T��S]�� ����)��c�o�1<���Z��K$�� ����=�+ܿ���1�Ӽ�!���C�)�'RlQ˚P$��j���牙yh�
}�r2�^,����� h6�'��VKJ�Y�D:��r9v�:�<-�����6s�Ϙ�����WZ�`���0aP� =��V��۶��@�]�b��^�����V�vZP�u�7\Am�L���Z��?H� �"8A�N�Y�� ܍#��):���Ɨ�2���o��&;Jg��4�Xߴ'��>bDM�r'g�+U�*pF5RWg�G*������5<7!?��TC�D�~���6�j����ȅw��gO'�l�3��k�l��	6u�4��m�z���CW�͘1�������]�a~e��97/�t�>E�웵���@��p$�.�H��>Ȍujѩ襷bԺe@ ̩Y�x������,#������&/����I`�I��q�4W<%�����Fk�}�1��Q�ʷ!|Hԋ�+���q(��a�P�����a�W��WkY퉺�.�F�ԯZ������(p�o<��v�"�������Y�����Pr��cØ_K�Q3�0�ʎc�]�2@���J�Oƕ��۲}����5nB d��u���t&�rC�Ĩt:\���zy^_�]��kjj�_�}��DV����u>��� �z]RKRA�%��Ȭʱ&#4����@�������3��O\m�-�	��ʞx�Y������|�E6y�����Ψ�"YY���&��R���� ���Qׂ��>�[���z&9�Xs4:$���N�,�C�.����wwC��_0lBm�	�hffHL%�⬕2ɠp:�Mb* 1|(���^^�	
!�3���#>k@e�P3�U�����{8Ppz��v���Ԓ&%2u;DK�P�Z0� �:�y2��p`�kw-_������r�����Ș+��%�3�u
�Ŝe�ߋ��u���{5ע�N�P�AH��ڪ�dД6�,�L�~���njk?R���R�HH���4�4�7D�cƌ���h�!0�u��u���[D�m'^j?1HǦM��_l�\H����'О_�z�s���1/��@���+���R�y̠����5ik;YZZ�'N|��':������0���S�����X5�r>M�tA��gf�4z@9(�w��!2�)�*�y� �c�y�&;U{�[�z���pc�8�s�B`�\�p�G�a���%�l���ߋA�*��h4N��7c�Uխe�\*u2����Fҷ.e-���h|h��{�W��]{��o��Oڨ��v�ճ�O_�^|��@�����t�FY�^Km32�{�u�����^s�@���#�!a��ͶK/��a�7Y���+/B�4���� ��Ӈ��V[��C�aɻ�q8��L���B!���~��;��=�q�ٰ֙0h�@���2���B
x;�3���o�cO>��U����|�N;w�v�c����S�6�,qwЇ�Z�d��ͥX&���R����y!3�Fݏ�?���g"B�O��׊z�E���(;V.��Z+D�Sh�wS:)��]��U��V������R������;�v����+�>����c(>��A�Euq�5�$o��?��h96�sQ��\��t��9�4 ���|n:���[�)H��5H?����bC�w�6�Ғ��e�H��T�8��@AA�T2����G\���˱��%G��k�w�C碼���Ƒ�rF`���e�\E���h�ޏ��I��ɯ�;X"p���_J�%��(scƎ�b#4DA�����ǐ�ݰ~��,�4S��Uu�fϞ���F�� ^�{��d
�Q���-�`�e6�VZj�p/���f��9���5'����[V�W:CO���!�v��4.޳wߟ6���arZ_�XV�e�Brrƕv"�#%S#��^zַ��e�n�UM���<k�oFe(�F^�lP�M�:ŧS��؊#�% �e�C;*�"2o�(��72 �[rf���S�"~��"�l�9t���NF�TO�:���u�R��5۾n��|k�M�;ϪАO%�o�(&3�*�LAuM]}$~���43#ڧ�,�4�/C�F��Ҋa��L���d�|����[wZ�qmm���CV��]���2�nt��!����u`xe�2�>�6v��&��!����v0��'��K9C�!�>֢����l��mv��B��eS��w{�����_}��n��s.���h�E�ܱ�PC�><�Xߡr���O)���Dbֿ��H�>�*�:ʂyyWZS�EN]=�w���ؕ��6|b9m�L�F������#׭������{�g�y\���ݧs�iz�'g�Ld$�1S��'Y�s����l+�r�?ٺ���`+=�&%�ҥH1G� A�4�&����	�շw��� � ��;`sf��١��Z������S�	��3�$��]��������f�%�[������ڗx�T̶3U���F�	� �M��jG��z	,�@�<�&�)�4>ʮ�_ nh�9��v��ސ���.|«X^�N/O�L��3��T����$�1�Jd:1�Y��{7C�`����N�S+����t,a�uI�ɵ+��Zz�7�p��:G�B��T��G�#7���\7U�?�����`�c�a���I�f�_���Ï~�Q�voO��fе8��a�����%�9�p����P��	̞�� �[|o��ˉ�%�:���y���'N����?��*߾��f���*dH����eZRMO��9��de���T��b��k?>�`m���� ,�̒X�h�@����z+Jg�x���?yj���0��=�E�N�ڦ5��n��n������X�]���Ѥ>���}`Z�z,bs�B�}��sv���=o?b�1�]IƷ���L3�~/`����7���G�/y��w(A���#��z�f虷�����=~�I�=��������]���a�x8��U��L;��<���Z��Z�g�E��);[s�%��OxQ�E�F� :@\AJ���]��C��E�0���Waמx�n#����c���'>�Y�c��G�c�`i�`Q|�ɸ��/�<��f\)���P�� >�W�/��F�*�<�#@Pl�Ъ⁯�,	��r���P�&|c��óLL@�[����:i$��_ �0�.��+��j�#�����]��X�?���1�V��m�a�۔=«��wp� �7y���N|	'}�J���2�C�.��B.0��ݽ������?�������<YSy�pNB[
"�{���9/����/Y�1��+��X�tÍv��6��*�#fؓŦ8����K~�u�O>��K�^u��.;�]����-Lk�`iL�]U)�y!"L"h]���P��u��@6"B��Z.�>��9�H{�������S��=i�|��XcȏR;�y�ݲ���]�A*�b^�\R���dk�}��n>z��/[ZxO�f���=1�0Y�2��Z��R�f�Xsy��G觑��,58��Z^�[��A�^ee��X�vz�M�y���N#;� � ��J�r�r T���S��V��å\C����z���P��8 J��$ 3i��8;g�U���,4��6g%���/���=�yWtSv���J����@Sߏc(G�+C9��	1�ɲ�9���a��� �qGO3;�9��qC��O���O3�F�&�3�_�U���o$5���܁P�Կ��,`�Ԯ�9=N�}�K2�P��`��%<uA���2�O���3�{;�,�)t�o��=v��W�V�O����7�����;��b7B&(�M
��E/gZ̈8�١��I�x�j�d9�2��L�f	ȯ����g�A`E��\���d���R$� 2�d}��w]���׊�n�!�W�8�!S��0�|Tٰ�ߡ��Ҭ2�a�ۙ��I)R��Y���B�9�$�01�1:e��:͐�?z�[7�t�k����t��_��΄w�c�&IJ��Q��������on�k�8�E����s��	����d�a$�%*pU�Yf!QE���+�
��g*to�n��p��3N؎��h]P�xUM�"*�
���Z!�1����X��s�Bֶn�{1کe1"e8-%U�,�\��c}�����sL�4������EZ��:~�*�&�bk������	F?�}���������+j��~������W��w#p^.I@��򄄜���G��������n�捌�;^��ड़*F�~qU>>t�F�Z���TN?s
���3㶁�{+Y`�\-��:���Ӓ�u����)t�)�B�K}CeYz��r�j+z�ez"�={��6t}�A$D廝0����3k=�g��؂M~��,.xhT���ƌ����(���'�:�;��8�,���%d1 ����Y����7���(�!���_!cyю��.}�!S�.A���F�.��~�//�;�'#qI�QqN�<�/�G_+��}ޡ_�܊�S���k���g���l����淿���?��}�����E��1�y����C>�$#j!����Ӣ=��7��2�󾯑�$�K?���{Ү�������F�k��m�Q��:z�ZQ l&{s�1����q��
�Xm��A������E���<���ԫ�?�:��p;���䁧}����4�t�訴��b@��be+�u΃_�}�k[<��QL�mU5�G�ZGi�ɫ$E����#��ju��E��K��t����"��03��jW�)KTq�d�'>	(�򬋪�x�PO&�9�"���w��oGW�^����t��\�������u�������x��C@�#�4����b"����gN"-�M�����o������m~��zP������뮸�_G��x�"pI��^(8W^y�oo��van��T�zq�"Y� �rK9,�:D�3�D+~�և��cj��po�Z��q������N߬��]%���V,&{���ぉ�t4�._��/�NƋ<��fbp6�{Wx����ݰ`��d<N�����q��d����1,�{ z��%*��!L�N��W�T)���"�������}�*Y \�n��d�RE�����8ۛ�1NٷJ�M,w��Ͱ�N�RoVF$I��8{u�T����z��t�Z?+�*���y�/������c�t-�T�ӏ=`���;w�{�n�]~��c��`S}�s�eA=�LuE�w���4Ctz��ص2�z�.�ڋ�U�Jz�)H�ǜ΄�~_���4Ui h%vR�Tp
�P4B99:���; �<�5� ��x�|�Y��<�A3�*���������j[^��l��^�f���`a��G�o��}Б�ˆ>�^���"۩�� ��Az}��OJ0L��)2��(����u_>F��MR�wr_r�(�әoS��S���f�>q���.;���@���@Y�*6AB#gaQ(����c6�)����U����
�t�J�/|\�	i�^�l��[*5� jbe⟈��\�}�.s�4�nWp�iDn�6�g��˔���w��E6�.i�/秺Z��N��
��~�\�z�%�ܿ�����-G�����ŏWCVڵ}r��lxb�V�xHX�Y��(%�¬��O<l[a�����4l���@2����
J�r	#6�y��WQA��z}���
 Moؾ%�4�G�,1����c��v�dٺ�J7�MML�Xf2��S��G���n�_f0�SW'�{�E���>��2C�Q����j���8���v��O������w��@<�(��R{[ױ)�f�U�I�1y �)-m]���dT�����oga�,Ki����΃;)�����u(R��ϐn�!* ���7h����e�q߻������[�G �.��ZZ�*��*q9`�ҭ	�$�ߢ�G(�'��Պ�s�q=����X�C*"�1/��?��� ��eb�C0(���C�B�������O�m��;�(�\G��� �P9�L[�>�\���s,&``���H�^����3����f��뼖���}_��i͐�\�J��t_�?K߻�3:SI��/]Bx�ms�s��Q~'���yo\`���/r�(O����T;�����k<�_`����	]�'t+ky�k�u���/A�P*�k����+6���G�����+!�����-�u�]�s+m=�<�]Z\xvÆy���{'�����x] �B���2�?��O}mzn�?Wf�6�U\G~`�O���sU�{-�e�����ǭ-k�(@���)������u7SƆ�̃��^��X;�-ǲ*J�����:E�|�	�xhH�M��f����Z��3����[��h��-��6�|d�j͛�+���22>�z0%�15�|6[D�by`��ob'{�5c�83�k�}�Y�b��K��!��,���z�>��՗ۅ."��&���]yK��Zi�g:���C>�1MQ��~]�Yh�d�����ud�2ȑ-�7��ЂKb,��Q�>�J�!{�=�����u���|)�s=\e��8��z�a���1��z��j�� �6���.=/��hA�dA�կ	�{� ��;�Ŵ�{�-Aa�ϡ��,���Q{{�s�����U��NJ�l�	��*1��U�)a�O=}���9�0&��l�{N6���w3�,��	�Z?r1., ��[qF�*Dz(��hq��0�Y}z��Ň�kU����"];�T��)|zX�^v�5~��^X$���,�|�O�� ��9*J:ά	,����m�ΰ�J� I�\1�F��|�2��n8ÿ����BEO���<�Տ}{��y�r�0ϗ��5������m���a�N,ظq�G`�/�a�{��k�����پ?>}z���>ɨ��@�	�C�L�3�t��+Kr�����8&-��l�k�Mu��K�̄T�j!��l���l<aY��Wd���l���a2<ҳe���R��֐���'�Izr��r�q� �t�c�B�,�X�S%�jԳ
�9W'���_ �|^��||.[aO<��m���|�}�k߱�j!֕U6��[�Λ�d-U��'6��By]~ީ����E���}��w����[\��[B"�.�#�<�}|J])�i�1�Y�z��/�k���[�J�s�Ry��c��f�u��8(N�o]�t�+�'w�^zz���?�H���e�dlQ'�ڧM�D٨�Bi�Чu�62��V��71�62R�$�6ʇ>j� ���WnG����4-
���K���,���B�qQ�5�<�)�7K� ����¹͌�_�x����R|ð:-z�,o��{ƞ�f�l��{'ɮ�9���81�޾};�dAZ�^
1Ք�D��×��1<$a;��]�o-R�!�������>�畆5ρt�-�%UD���ӻ�96{����m�'Kva�{�d'v�=T�V���0����w����������#�>�;@�	2#{`bj���ǎ���yu�۽��!;���WLs�v-1*�Xg�y䁇l3���8���z)�Y����J�� 8� ��y�$&i��S�?wv�e8��}6;0�K鉆Wx��,١[Ie<�X���V�+���,�GP	[˾�\�ƒtti��z;7��70F�qZ��CnA'��E��+�?Oò����3�Z��(y7�I����=��k������A*r[��$��¶�C^x.��1J���BP�h��XHq�>�8�a{�mo���/�Y��Y#�_X�'�O��%9>���K��/w?��"����q%�t�Yb}'��Z��u�r!bJ���"-9�)�6�土L~ q�N`닀�L<t9D�SN)y�F�"�)��)m��=�9�C�K���3 ���ă+[q�!���1�5��ғd���{n��E����S,��$�޼K����N�1	�s��	6�ry[�]O%�u�ɚe;}��ڱë �[��Ҁ����ҩ{__�	���A���"�X�@��j�GA��3��믾����>���1{�?ꤹ弄j�^����-[6�����8��R~��{^��.]�knl��i|���??21��0Hh�`~TJnC�#�;θ�G)e��J���S�N:b2=�f(Wg����v�\[��\�OS��3��9�z1]��Ӈ��g����W��x��<a�C�q���y�Z�� Op��˽��9U<D҇�g*^*\˰��EŚ�J��7a�gg��Zc[��ֶځ�?i����

p�2͡j��;��U>��u����^|7�Y����%l^���/i	8�~�Z����P��/tɫ�F�D2�,>EZf��X�V��s�I$k��󟶪/������s��ֻl��ݗ{^�HLs�Ƀ���YR�U�!��W֓��R�����1�rp8?�4��e�*�!��\�L�F�t��X��w�YTrq䤡.g�F�T4b5::��U*+d ��9d��θ�:�Wk���j<NZD�OZ%����c��\k1��̻�=�K�����~K��9���S���g��PQl�b�Q<ɮ��b&⪷�t';]swx��k"��isjҾ�{��]�ԉ��Uy�k�sM{�����
,�1�I����c����
�X�4&F!�^u�����Ǿ��x�=�:��iS�D�ӿ������y7u�G��E��-���ݹg�;u�Է�~*�������>;~���"��@+(�f��B��sCh����Lp%�=����1���Av)Ne�F��ռ_@$�eۀJ�)׎Wf,��iN���d�:��z���1f����z	`  #3��0SʻzX��5)�**�_��d]���cdu���"���$3��u�\������ࣁ��R���fZ5vI_f��s(ͮ1�C�w~�]��eΤ��	��X�<T(|+���/�y1����P���XF2�2���Ӝ�b!� �URF	{Q��fM����}ڮ<s��ۭ���g��!A�T �+Q-�ڒ��*��kվtp�mP��>�WҌ��P|�$K�z(m��;/���^p���2O����/a�t�2禲����%^�Hj�>�߸	U�����5���W؍7]���u�wΉ�*���1^�9+��W�ܴ`�A��t\)P�ew�����TI/$�k�\�d�/��}��gO+E3�ȓ�G��O#�sZ�h�Jn�-�����}�g�5������h��*�7�z�=�ēԦ,�W�5�]�� 5�T�<ո>�%]�2�c��ٹ�Sv�m�ہ'fn/�Ѣ�O�E��#�c�V��"��`7����X�K�rՖ��iq���/���ɳ;F��s"�t�1�'�������Co����ܵm+�~�NA<Ӭz��x����d��	�ѷ����f�~d�lj�`a���1o\�ͨt��aj�����Z�b��CV�S[K��(uGh=V��q�('`�GW�R�'����ܘş�Fe����X�vw�ﱶ�z��ۑ�;���,��##VG@�%�i��>��� �Z��
���i҃^���5e����k��ex������z%K�(�|���x�������������M$vA2��Z�>� o��.�߹��,�(�k���W��FƟ�"2�,!L��!(��=#R0rU���s^ߒH�!�'��(�������ʍ�ʹ��1ǁ���h���;�X؆���׵0/-�挷I��W�w�S׵S�@���W1�񥫖P�y��B���7�����s�}�1K�����r���{[��M����f�_~���;�%��U���9�ꋈ�A^%{��*�������Bv?k7�x>���cl�e��[�Ԅ>D��Z� ��/}�ef���ְ�`�(�G����۵��/vğ���Xcļ�G�*�ĩ+.��c��U_��&Y�oG�f���ۘa�/8#+��̙3�^���"�Cd��=���*!'-W�`��ՠ2�6�umm����RF}����5��EG���<�k�x�d}�I�.W��ô��&����^���&�Ck,�&JZ �x�=����V8��7�ͯ�c�~�*�!!c��w�l�µ���ˉ|u����-�Xp- ��%��Ҳs�X*7�����ů璬��<!�%킠�db���X<LZ�J����bF���3xȯ��]����>�&�]�s�>�g��'��_�k[=Aeb��4� �����4��)| ]]�����):��i(��x������)�>�{q�^d�E2�eq�hAp|j����#9<��o��O���1�p�hka����4�Ct����phѤ����s�uM�[���zo����Wدvr�0�؍�/��H���T�կ��R�=-Nt��&R��$>�[�l�8E#�~ӆ~��C�9A�]���s��O~Ҏ��~��+街ؑ�g�o�3�p_�x�����ӈ���g>c�[���oz�=2|&b�Jx����-̟�
��_LxCd��߽{�'N<���_,�O�oBI�r�E� 39�J=�|VR�����Zu��nرF&�K=���Đ��Dk`�.ef����>��w�PEPd\'���X�������bϭ]�D}���\����g߯E�{��*��1qd_��Uَ��g�+쫏�'��}��'�mo��EǄu�m�7]����ѧ)�ŰPN�r@h.���z���5i?��M� ��⦫�)R^1>��A�τ��굗~$���w���}��$t�!ѯ�l�f����!kI�T��'����k��	���s{���ڑ����t����C�x��xD�?4$�2+�nRJ��/h�)8g�ii�xDO�H��~{k�P;�Q�Y���rg����淾�~�' ��V���=��i�å�� FҶ�N�{"d��bW�]�%��]-����1�m���E��-����=y��U.��k�J�������E��R�V�"����H���!E�z��Um�,���O0���%W��<�[�}hp	픃�b�3��%Bx��Qtݯ�#ǎ3��l7�|�I�{����U�Ƴ��_�?�i�m,���I���o�����z'_�<��c.��� ]A���}��-ǎ����/m�=��ϡ�6��)~.�����`Ԩ��F}�i{��l۾�d��6�vf��3C��0�F����2y9���M$(���Z�~c,���2�1$;u���Ѐ�9��i��R��2qe�<]�0�@�Y�,��z�kN]�хe$`�~��c�>n��]��滬q��E���	�K�����Y]N+�*ִ�m�w���֔�_��] d_N$���ZY�1��a�x?cY��X���H]�����+R�J{��
�i��*�gh�]��tyo�@RD]��Ƀ������a�f4�ń�TK���ᗐ���d���B�ȓ�A�x�����+|_����T��CU,�,�9)���~���ko�΅b�yK ;�Y�QJ�.�J���^z:�{5��~W[���|���<3N\�8�p����=uG��{HO�qI>�{ڂПr�M�k5�A��Lk�ܳ����F+�'�aĐ��<���o�sQ���R{JxR�[]\x�C%AQ��+_�����;���5~_΄QL�s�-7{�C', ׾��8e���w�w��}t�ł/���p���?��њ���w���\�xC�.�J���#�������ߪ�.m�l����ggP��T��+al�2��'��	����ͻl f@�����t��N1�ޞ-��-����*����f�ǃ��RrsK��̬C�Qf�a���2$����)��8��y�(SЃN���Z�aJүC�����+�<k���˕�y���|��zW���G��z�N`S�Rs�<�Ha����tgګ ��5�cǎ�V҇��n��x1�CI;d��\�,ź��}8Xu:p��-}�e��9Ff)_��+0.���j�#�3��$��>�&q���7�gev��a�,���n�I��)�Bt�t��B�*���*j�&ǯ�kQ`]I{=g�x�t�~t)�=e����}��h�T�jG4�N��uv�O7�X����i��!8-�2�]�J��rm���>���U��x�R`�=z_���TuTr���P�N��6���}�'���\q�.�K%կ;qK�w$�Y��Н��<������F���6˖��� i�k�_��G"�`��)!|o󇑍���R���^T�g~��k���r��=1Sް��^�m۷������Ν�sطW6�'Z����P����0)��@�����
�W��Icz'�2�
Htd�Y��hf�6k�M�Sf_ ��q���6���l�����c��!�16�ٺ`֙�k%`w������&��J���t��Y �,���Q����H�ҞX��?��u�fDG��lS
w^�'�]-�"�d��=cϡ����t�h��V���ӻ$��C�K�g�V��؀��U�ٛ�<>�2->����$�q��Ve��i�p�o>˵�1�	�ŉʹJ�l�F��׀̐���9������m8e��t�Պ	�D���p��e�_�5p�f=^����� �T\��m���,���)�Cƕ�D+�t�_��$�|��e2t�R>���'"1?��z2��
��ϓ����*�Ƀ�Mhs�qρ��.��D�h5�{��AF�n���߻a#Ğ?��u�?�b3r�����}�+H�؛n�����#G)�ov���}�{vvh�>�Ꮲ���<Q]D٩�����j��Q�,n;F�G���G��Kd�8TU?~��f���L�'8��I>z�%b��Lrd�9���s�Yl}��&Da�V����L3a�9z�<�f���
���쌗gg���!e:�P�4U��-�n�^�Ǻg�����6��̪�>3�w�Yl9�N��Ov���d�fj�{�&-�ht��q%��S��vr�/���T6}0�e;譻�I56� r�B'd`��f��+�ݻ���X��˔���C�A�sp��_�̣��%x�qeV���S�ֱ����C2U��eA��2v�^���DN�c����w�B�޺ϸ����R���D(�ǵJU���p�Y�(��*�/������P�i�;GBٸ�t0੾h��ן>_�R{��yWD1N_�E?]�VK�E�I���V ��Wz���y�����!K2h����|^�-�����a�����q_�����3gΜ�&�H(�3g>6��
V-�G��Ss����<�����g�)�ٵs�} ���07�x��޹�������4x��+_�:DČ�y�]^9��r�Tsc��\�ϗ�h�G��%�7|��^+������G�026�G������^�m��8y�3� �������v�c�͐���8f�[)����N͌�p^�^H8%+��!�%���J<�˙_���-ͥv�쬍��1-��jkcc�D&	h(��%��릞f��>�9�Uin����43��/
�d���Ϝk8d��G��PL�qMn���ʷan:-yz&��1�+�V�"����ł΂Ő��.@J�%������۽ݶn�A��j��0� \���ƴ�R����(�Jo��P	q�>@%�:SdR���f}Q��\��K��8������-'/�"��圏���Ffw*?kS_��m=��]�[������{�[Y_)3�j{8�z�;�y�6Tt�~1��	���! -�����t�$?��z ��Ѫ��*��*��8�d��<x������\B�8P��9�0Y\h�*%�E�9�$xK��AJXK�g�>5��S�!$��u�+�"d�����P�j87�~8��~�Wd�R��a���g�W�BB�w�ŝ� �ۢ[s�A�{��C�����`Ϟ8joA��[߼����w��������A����/|G��厷�¨�	����c�]�?�{����г;j��s"}]H�o�����C�ы��L���M�_�g�>~���T S&˔r�k0t��X3��Ɣ�ڽC�j�\-6BF?��eOc9�8)��hz��ì���^SJo��b����B�f�mW;�Ml�d�!N����
���N���؄	H9�G\��h�V��������r%{�XWA���?�5A��Y�!��,[`���o���Ҷ.�򠒁�|RV_a����i�L��XO%�����B(lnk��X�ޢ���	���|�ј]���|�h_�W� G&����}F�s��?�r��Hه16ޫŀo�(�aCz�� �nD �u��w��	����W]i�����j�Y(N5��m H�J�	����pr������D� ��y�c�M�:�,���c�u~+3�([�����l���}}��O�k���� ���s�I��cX�b����rZ�%Q���+	�q�n��6��f�v��`Ky>�M��-Pt��f�!�ܞ�6�Y��4[cs�]v�>�MTŨv@Zݿw���g�q��g?�Y��7���[҇�}��o�����Ǌ8�b.�D@��������o{���Q���*���m�~�U�&�qx��'��PM�m����߿�Ѷ+!��d����Bg<_�X���|��yv�L"����W3:'��3��dHx^v�>dΒ����li�[�q���z�F�d��4�̲��z���r�C�3n�-B�K�hh5�JJ�wu^��O|B\J�=h�+��`:^�<l��\F������E��.��9�R�������J<9?tI�'��Io�����[�Rz;��T88gi�g��N�drd{:�,��0��Z��ܘsǍ���	����肍L��A�ܔ}��߂Hx�n��N<��%Z�lOq�hXXaL.!�y����V>Y�PzW�C��5.	�~9$-i����Y2��\�5��d�b �|��d���
 y�����s[I���U�"�]ҎP�8��˼��	T~/�Z��lOO\���� �B��m(U]������x��߅w���0�q���NU�*;v�b���u�����h���f��X�w�.+��qߖ-?���+j�_�8�>�@��.߻�ߜ>u����x1��у!F�2�1Ș�!!�լ�ri��Զ�C�'���M����I�t�����@Oc���&�����Ar�Mn��+J�g}pp�L{�^�J��xS/��'}~v�'�HE�������f}g�7����H�4 IT�Q B'ݏ_��p�eR@�:���N;��s�/�z�`��BW5��>�6�����>`���@YO��G�~�v��/'C/�3gN�Z.��İơ@��=u�(6C�[B�o~�r�#cqTUQGvK�^���<8�_>w�����,�	?���#��1��bch�����e9{*��m�����ʮ��M���k�ȢU�|-PT�#b��VD8���b ��u��Ǌ52�X��#i��o�����ꓫ<$��_�^i����:���/p/ȋ�)z_��M����8��Yk�[+�?��ɷ��'�?�p��y��&�!�|��eۏ<N��z�ۤ���U�zQ�]#����!ޔ�f�d�T'%Gݣ�ã���m׮�v��\�Ml�eeI-4�#���}����|�u1�!�yU�*2+���o�?.����K6�_���m����O�:�	J�o�1��-d눼�2�À���
l���O��Sƾ{��[�l0Ɏ��Ȃmom�z����^xf�斱�Ԩ�SSXAS/���Q�R�c�[��F���Y�!��j6	%k�\�R֚��ٳt���)G;��㢈q����gRn�>j���IH�x���GѴ��^�����´�E2�uȔbiY�b-�6?6�����������9�lW�u�CF�݇ԫ�iߧ���,����Qv�Pf_���mjl��=�q}xA����>ʬ����Y�f@9e�y�=~��!6PQ���>*A����l���^M�Ʀ1BYp%g߿�k����n��Z�7����������X�f��e�k�'��T-XT��jE��*2s����fW�d��Tev}���5������Ck� ����n�4����������d����JXT�e� ފK
�a��p��e�Ӫ�0��2�v��1{�;���T{D3����2��Yq�<��{﵏~���0�xc!��Ï0[~��,n��z&"�)g��	2�*AO����#��(���O��\�瘊������?]�O�x�1���/��hnm�mw?}��ώO��fUeu]wk# dvK֕rdá���'s瓐�z�ۿ}�5!8���Ll�=;��mMKVS6k嘱,�@��K����9K��}uJ�Xe�a�;<<��D�@��}5C�(�q�og�=ʗ�Fɹ��,�'iL2@��ON���Jy.l;|"���R�HH	!��5
�VW�dM�.Xwk��Bx��I��F,K	<?�(��pv�ng��ܳpz��X��:{��'�P�(��9�L�M"2O�:v�Đm'�����R���֝�8%J�d\��x��O:J��C[]��p��"���u�#�C�j #�����f�W��4��L-��s{��>e_��_�5���
�x5 ����ʿ]�6��E�3�tQ���U���*;r_S�W/��r$o+d��W�Z&1����%�ߵ�K��ѯ�u��>�����e�y]K׶�v�qL��8r%�R��:�;�]H�����Ͻ':.�`�_e5�g��v��7�gL�U�t��g6N�=�������?�s��.��	���~��D�X�..�5�V��5�]�g/��>�%F���@����޵��N������'	��]͔�y��;�y�Y�d�<�5��%|�чl*tw�A���\����I�Z�Z�_U��	����N������;�c����]����9�(c��3e��	��f��`]Y��JҐ�dt�f(2�����$������y!�����'!��0)��7����jk����:�\���l<�=�,ŵj��~�i�&�0�z��|oǰ��tg?YYΆf�2�ό~y���$��'�9,���Cjv�>��/P�F_��N�%���7��c� �/��m�.o���	!�Ş9|�h�p������S+%�g�&P¯%[��<툳l��۹��2}z�Ŀ��ľ����Sv��o���n7�)��E���Xe�V�*��誨 �R�e��>~K3]1�UA�v�Į6��&1_ƫċ3�t�����}"����Bǝ�XT�Ci1��ԩ��Rܵ�iM����'�0O���O�����d�^{��h�aav���UZ[�䙳n�����"o_��W-������K�_h��ܹ�����|��Ͽ�pƏ�\����^��ޞ����t�̙���/vS�mon&Su!�|I�P���pY!;;z��-�Q��*ˠ6]�a��~��0z���S��ku�z��s�}J�O�2J���<;j��y��$L�Ef��/w�����ٌ�T������˲Uҩ^@9N���!;N�q����<��J�z��J����.kZ�����|ɚ̩��e6;)�O��%�H�"S�`��Ы���ώۙ�>`��>��c������ 2�۶n���ǢQ:� �U��ͷ�I$<��o~���`W?�{�=l�����v�5�1~��QS�ѝa�8��,y��}631�3�]���ZDI[�"Sτs�'��F����[8�
J�d��N�7�:�z�}[� D�J��'�w��餷�m������QD>I�
�+�er1e���-�n0�Y��Ѳ����t}���n_�r� �//)�?o���y����6��(�{��Ps�9=M!��^�g��j�8]X��������Vx!�a������:������������Ҁ��/��׬���;o��:�$g�����=?�}ۦG^,^��1�r�;�z)�ͫt��������K55���%󳶽�&�g�d5bUE�������(���{�~[���.����^�e'f���t9%�>�� [�܊U�(��R��-W��쵍�m6v���u``�&����ًg��;(�1�R���^&Fۜ��c�mYsۡ��Y�&��X��k��֌��^eY�m����{����()E*�����ib
)�9�M�H�g�C����f ����& �-P�?�ȳV�z�Xϭ���[mna�N��s���?��+b*�m�,P�gJ�	�ހY��И����VV�dc�r;|z�3m1�#S���mm���~��ޅ@Д;�u�l��h�,�����"��n��i�#���� �t �
�=J^Z?�����>g��CV���%t��מ����MR4���ԯGV=����U�q<1��y����i,����9�Z�h[�I�\h��]׮x�=헯��2��&~g�+1k�)?�?�|�Ň��$_�8.Q�|�$����b�u����H�o.E@M+�^�}���}��<��d�,�0^��~���m�!jI@�4�@+G�%�Y�����L-|�3_��Un��I)Y$U~?���������1��5�@��_F�w����3g�\{nh�K��;��`���f'aw��Lx�O4*u��(1.���#�<wj���\��-7:e� x5�eD2���i]l��Ô���w�,��f�ϝaƽd��1������w�@K�ڿ��UA>T/φx0�Lt�_8kz0a>Z�c�Ĩ�r><�!'-�/X�p�l,��}���-L�R�_���[�N	����uY�yb Ô[�@+�� ������u����7S���^�$F5r"�`6��[�[�dO=u�v�鷍�730�c�;��!��Q'�� �|fǦ^DD�(�3�AO�MۜF��`ؒ[,���:�u؞��&�z�T?*)d�=��B�,,f�๳H��ێ=���^��;2|22�͐K�U׫ ����Wp▩��D8ٿ�?��2näT�v-�Y����9qϛ��r�/�_b?ϫ���\�O�p��ҩ	-6�'�*�>�{Q%
�Ы���Sj/�z�����y�n��6'j�P�:�.�B����7_�~��9�=,�;��̔}��o��{z�q!�b^����2/��$Hq灃��˹l�W�%߶��2�JmЁ��:���:)������ݻ�����_�	1�Ҏ�Y[����� �ZK[��9;���;�~'��MAr;wn��L"�:JK)�0X؁�z�nI�;���I=�<emW[�K!٤�%+�"Ki#��h�{�N������$\,.!����5i���[�ӗ����]�� ���+o�/���5h�GP��A齽����ZYc�]y���/|���es�]y�V:��j��$;:�쮮}�H�+=}��8�r��Dn��p��{�W�1*�;���{[Ms�<�8]��N�<c�K�M4,-JK�+թ�*���
e�R�{��o#Wz�.��zι�eJ�e�U#��Y��r��0�B�c���s�'�.�g߉�yz�����]�̻����~��j�?���"����/��	�ۘ$�\�E�	��<�2���g*�ة^^/!V�L������w�?���}HE�
�"�}��9�Ҿiw�����X|��TV����^�s?��ŏ�\����
]��{v�Ƒ�G���}��;7�n�����OA���K �Ze�����ON٣���.��JI>Yء�a��m�ӂ�	��Dv��ۯakѦ y�/6Q:��G=dgO�z�e�ӈ4'�K����z������I�r�Lb�sC��*D, v���[�*�Z������� X���v����Z-�J�H���k����4�[3�泥YJ�S^��݌(QIhmԃ�G3�8{@��rw;'k���c��+��}�Ȃs����_<�jZ�E��h+ac�ދU�`��~�Q?�ݪ�����-�.��R�{�����D��������.ƿ���e��baQU����V���i���T��o�=1�A>V��lX��r��r�3���(&s�4R�ӗGy z!6�y������0](�}a�}���d_�q9qPD6?�C~�P ��}�9�&�'?���f<���3��8�/���z׻l���̼��!P�E�}��G�Ǟ��C~���׮\����/_͕��N;~8F��@�W�m۾�����N��Ӆ|��&DVvn߁��)�-'�ha��,'�n D���~�\�vZG����no;=:d ��Z� ����l�2��h�h-l���3#�Id���h�F�	��ʞ��[V�h[��B��4J��e`�n��;�쳫��n��2�^����w}�Bee�sq�6�)UJ�yx/�D���̯$�昧�@0��y�����-g�mn���\�j�Ʀ����5�t[W3Ûm�N��Ϟ��'N[������׺d��»�+�%=��\5X�����{� 8+9�
I��w�4�� �1�e��9�����
E�:�q�$U(�IF֫�h@N�"Lbe��tW�c�?�<p�v\v%<�F�ƩP�[%�tn��E:�ny�+���W�t�\HOMjRw����L�g˓�=��/DB �y���N�[������Kw@�t���p��X�� �1�%���%��թ^!��J�g>�Y���v�UW�n�$-��kﲓ���������V��l���]�؞8n��Gp-��u5����+���+�k7#p�D �+|�::�4���G�8���QS^�l�Fa�yt��:f��P���%��Oǎu�v�"U��� V`<�8%�n ����Db(���F6^�gk0y��d_ǌ� �>A����e�g�`-���e�T��2n�6K2�b7�@f
�z�Ho��f@��+ʛ�TTsv�U���vJ�m�4�{;O\�/��Uoƾ��E�/0zƑ���?�����t�ێm؆B4[A��L��^�@����FI����Ĝ�{��0���Ygs3���?I�.��Z�׵�~~~ŪUކ��j��9"���iWw7a�ʸ�Ш=��1놫0:4�⤂������Y7L�R�i��t��!ɋ�|k]����Y��MpP�a_F��h��
�� UOS���s�b�u~���������{x���K]$����~�2�A�A��b�5p~�-��o�wv��vǝofA(�ga)2"o��hy�a��[�~X���o~�&h=}����@�W�S�����=;��
�,n&F���@��%��=�~���/�MM�	p�cSG+Y`���X5�����Ƨ�K�n�����pՊ���
lyV�8�s��5@�Ä��R|^^f2��I����jf�G �I�dͳK�4p��hE�he�, |V��� q���5-w�����q{����u��3�ҳSz �q�`YWVJ"5~Q#{�E �<i�L3V4�nAnu��rWS���"g6����6>2��uKc�����Ƕ䇾��IS��J�t2�%���]��ΒaOCj[��r�$�7�,:tƝd�NT�ȟBe��k=��}y1�>
���>��P�c�PB4���GbNS�(���@KW����w[#cp��9f�k�Х1�2t4^��r)��Z�^��o��z13���M_*������1G�ĩHH��f����s⽏O
핉O"��������`�c|ķ���m��Sv��W[_W���}�_����o�ہ߽�
��t���έ�O�b�7#p	F ���mۺ��ё��N��C2��t����w����/�e�E�[`L������m�.63�z��'}-<�P��,t��V�x���U�V��0̫���a?���A�E��X�I�E�n�*ܝL]O(ӺQ�)��0�d~����[������)��+HmR�/������:ܔ糰ʳ̎����8%�<d�e|]��6t 3h��=cKx��q��|��~[eu���#?c=�coB4$#)P�����[�1 ��  �
S�n��'�Glk�*�YM��@ �֝0�.������7���v���һ�~%���/�>!rA6s� �Αcڰy���a��|-��Z�#W8��ņ�u���W䵝�7��f��x�/�=�{�7k�
ޟZ <�tw~ƾ~�}����SL�K��a�w�_���J�󾿌�J�l������JHfB�����m��N<�����')���mݻ���d�M}�B���7m�����3�`��b.�D@�_���.���O|����~��<S�s�&��O/��z� #K�\����9q����������3=6����p��u FS�$��L�1e��<�-�^���ş97iã���e�� {����<��X,�S��"�1I�J\],y�on��cM���ui�����}��3c���0��=p3��g�l\}�R-J���R��/���l��[��Ŷ>k�w�'�_�G��� #ph���R	x�1�]��t�R�
a���+6r%S�V��t[����	�.�x`���n�7�FG}�O�*�
����o�3um������p��=o߲�6t��V�`Y�m�7,��"U=J�9�+T#�;��{?����i7 J>����*�e���N{܀�~�j~k��*~9�aU�Fh';��Ac�����d��=�`P�L��e�ȼ"���CI<,��+̑KQ0, .�CO�Y�r��W|���4w�"z~�\4�0�śF�D, �G�y�~�g�
�I0	���N�i�dde�8k���K_�n���V�ͭt���Om�������fF2�bb"��J���=����S_9;2�ǥ+KWv�5�G�EL��k�G��M�g�5�a��#<�߳�:[m
��ٹyL*
d�yی�wM	ٺ@���,�)����j%��@쪪�3�s�/}8'�	ܒYta.)��Ürw�^۾k����`@���ݏW�(�]��-6|9��G��F���6�mc���	�T7�,���k�k�nʧv��#69z��R;~�<x���r���<o%b�S�V�@`���\��չy�2a��<`.p�t( �Ly^.]�/<W!d�b,.������T�j������_�]�ȿs� ������zFNu������ŶU��6w�<�z�ك:����P�V�y���b#ij���Y[�pOލP�v���]^͖P�	�lސ��J]�R���������?�S�ņ�҈��Ȣ+�:J;Z�R���S��T�H�m�[Z �TE���="��3g���K{�;�em�]#��\��J��k���W��7�&F���@�W�2m���������O��m�+���̬�#Sc��Pi�<�j[�
�����-�6[*g%u�P'ƭ����&LQ���]YGyr�0#R��2��k(W�Na:��DP�d��]_�-_�X`�ˢu9�u��ۿ˺{�0����s�l=U�%���Н��:��Ӳbď�!���XDp>�0���][%�&��v�Gm�$���)F猇7nYX�Ճ���̨ﶇ���75x�$rB�@"#�S_s�d�di��z�Z�`y���Ċ��NX��d`��N�Ve���E����zN�,��o.1j�vG���_D(g��	�_q	;�����3�)c-�4Z��؋2�����9����^����ymk�����_� =}ye�g��@�ݢ;���.��FJ�Z�(�.6�)��_h���ƴ^�X�B��B�00��ٳ���ʉ'BD�%���o�;�q���>�R�#�����|���`UEſ���+~���<�<F������hk�g�?���_����OKK];�?��>2����l�T�����SH��ٶ����{�S�~��}�"�]�
Ӱ�ˬ��RY�M��P&�2�e�z쑓 Z��\��Զ���U��0܄F��W�bT���P�y\˶0Rw��a[D5k}��0�3���%J�Ӆ1�l鰕, EF>���
m���d���/ڽ���M��Ѐ}�[ߵ���C�F�����ֻ�i�/~񋶩��g�5�'�WY�ʁ�Kԡ��2�*g��?�
}���Hȝ�<�)���_צ*��s�&�=G������s��U���
�ܗ'���i7�|�ghe���z!�jji�5��,
&7���zW��ݮ鵧��T���܆�d(Q{I��b��^$8�
���d������5^�k�nwE;)&�=߾C!d���&=�jb��t�B �'s_b��{����	̏Ô�^���Q���a���~�kF���5�V���]��^�ŏ�y�E �kt�wo��Ɂ�����~r!���	bUu�&;58�?��-@�R�] $��v��ԃ����;����F`��k�,��S��-㖦HZ���\�oӲ����l�8��^ C-�"K�an�ٮ�r$2(zd��e�+�4�(�jxPϏ�6@���1�G;n}���� ��M��Ȟ���}��0~w��;��7,˘Z;���[;$�A��2*��}�ڛ���i۵�:���o����Ȑ��>�x(@!�w��M��eEZ��*;N��t�PX!R����9qe����N0F��D.�����bZ��SB0�h��#c;o`����S�����dA�<�Չc]괦[*���l\�H{�봏��Ӟ3^�ܷ��`u.\����g�r���,��Q
H�e� �8|�EI;��Q��J���I�M����6�(;o��Ӟ{0r�=�2Ծ�į���`/�ߎF��O?�o~�m��\A'k_��7l��}��R�9 ��lgS�O�ݻ�;�ѯl�m��E���%���=5==s����
W�@��== ˨[~��]Y&�Z��*4����6o�����Ε�C����5na^�=�2ɰbRC��!dbe{���J�4k�<sc�ِc���k�ߊ��F���$�ge�d�<�����̡1�WBx��?k��p+�|������S�����8��������F[����߷S�Y�� ���cOr#����k��tv���6@�޽���U��ە��L H�~�}e@��t�+������>7��2f�ݯ��M����vqR/�>�������JHr2U�$���nɻ\LvMU�׭}ka�qc���,��iH���|���h̎�K���̉	�#zzcij`��J��;xY��䞺�=I<�Շ>��y�`��O���G~�c�ؐ�]uEC d�#b��;�����u�A0�O��3����Z(��J�^�z�Q������z�j���}�X��]���CtF|����{;;?�sۖ�/+h��1��D@�/pCC��[��ȉ�_Z�����b���}r2���Q�
K �,��Ͱ�j��)�t��#��jzꥭ�����q�(X%�
2K��^wÍ(p���s���ѓ̺���^��kM�d� ��bIr�)#ۯ����9��fx�.v�o�_i�����V�B�4nk�����6<�	+mh��d�ff� ��O`Y�Pc���ia|i�-Ly��Ajۈ��3�`̲�*pa�KZ�^`���ܻ�G�v����� sK�H��K��:��,�4��rz�yƠVX9�$ �`��: P ,�X8�i֝��{fR��WW��	e�vٯ����sU��A~#q�6�/�^�$I_�P]w�c��'�=�w�"�k��H��M���I����� �)Urb�,�ƴ�J�:>)򩯞���H|�O#�pԏ� �D�-%�hU2��m����4֔2E1�������6ȓ7\#��Y���@�3�7|�C_d���Ϫ���?�/�k������48:�I�B�-on��Vc'��j6�k������Sc��C�S�߉�H7%�FW����S���Qc��et�<����ط�v�]�-�q�ǔ�)�/3#����f���Ȣ�Hy�����Q����њe^���Fe�e����&;y�8�U�>(������4�sn�HMM-��¸W3z�gN��	攀���[��
m"�)��"�d�*ե�z#�ֺJ싰�+0Q�M�)�0���n�~6?���}ZWjs�9��	WO�]N�!/�'+?�I�@�3.�
��<��B��q�ↇ:Z�>���.1ӂ`53-���/�MK�~N/�J:~�'�k� 7��%es�;�����xC�,��R���Y�0���s�4�������c����VPp�Αw��C9����	ټ�.kLp�>�7_�n�Ŷ�V�YS\����Ol���]�]/�/q��.�Èx�"������������ܛN�9�-,d�f�&�熇]�m)�w��#Y<tss3����o�uo��m�J��L��3gl;Yd{�g̞W������z@!��B���4�ky�F��@���T֔-�y�.�}+KI�%��1Fwy�.��@��m�@I��zɦ��n�u쩇����c���*���ZPa������au�� �$YR����۷���ag@Y7�P��}����=��h�m�}�ɀJ�T��)�sʑQW@���@�c����myT��{%;�4l``�򳣍�h��q�;z��oا�"��*�;ˆ�鎍k�Vk�ϟm�g�S� �Ņ3��9,�����)(�4Y�@�[��W�FH��^%� ��sk�Ţ��'��m�� ����y�-/�?��=H��]�����W�g`-�CH�ǭ��S)?��+������S1"��}����@\��e���ϳتc�'�Z��j <�F�_������ZOO��gd�c�u�7��E��%F࢏@��5�Ւ&�/<{��'��~��,�U�Ӆ�˴C��g}�u����
5v������ff=��Dd��� n`��l�f�����,V�G��0/0�h�٢<�2, �x&�6��Ȗs29���c�}��ey�����R�OK��g�� ������������
wl{��-��Y� ���<��N��v��;vo�Zƾ���Ń
��
�@�[����TM8{��2�.��˺�ˮ�{�1���s�f����;��>_^��2��(��N��1�����0�L ,Qq�"c�Ty��|�{Zuc�m��&F֤����ԍ[B&��z�{Yy fun�'���L����y��u��zR�y�����`��x���'��ɂ� �3lo{�[q�;m;wwy������-\H�N�]t�������H��U{BNk��p�ze�bD��#�%��}߹����H���P���3�����o����W3N��E���%ڱeӧ�F�38:��+���%DC	~`p�r;sШ�e0D� �u ����=��wm%˦�NC���}+�!���)��׎�jY*�4���Z[��L���xK�G�g�
,�iJ��[]"�e����w�J�����r�Y}3�T�Գ���aH��=��!���~�m̬��h2F��3�=����[8�j��^-����z��Q��癝�&B�J���IK�nh��;3�B~���J�ln`�2�+d��g�s�VN�^����x	چ�S���������?}�:J��M�X,@v�_�˗�'��ϭw�Fk��壜=��ǭ:%�#��J��-����.B�r=b:�[�h}�=ғ��|aQ��S���Xt?�f}+~���0�wQ�(����m���['����\�׺�K���:�V��",�!�tJ���Ȕ��1�*�N�4�$�����~�*�n�%��隚ꟹ��}_|ig�##P�������vfjv���g���\���R����b9���_�̼B9���~Y�>p�6mZ�����ȧ*[)���W����M�@���%C$����*����f�M6�2�Z�ㅊۃ��TvҞ��3_���ܱͮؽ�=�,f*�x�W1^��L��0_ކ�{�_�G~����߆P�����f䌯*�����w�Mٳ�q :E� �*2��������������c�F�;�9�X7���z�붫�76*T�h/�eh��r�fD{fr�<�I܂]�{'d��}�/�`?�w�6�e��{�EG�)�S�4��vϴ��'�h��iV^��L 6�H�z�^�'�� �:��oДq��~,]�_���]J:�.�i%EX���Z�N��\:��{���N���W������ܝ9�̹���Қ�v4��_f�[�"o9(��&���U$��F=0�&_�O��b��N�0v�8Qc�R�F��@}΢����X�
��~�\����h�Ϯ+x*�tr�}��ŭ�C�i�n2�`2��L��W�406�oUnYZ����3W�C���?4}�cd�r�o���n�o�4�{�>��ζc�K��}Z��oLS����<'%vHG�Ê���E�ѕ��Ű��G�t�t9).�l\q`��?�P�;�D���s���nEy?R�eɼ��4�;�-�g7A!<`�H�� B�U{w؇58�U�i��ENÍH��#�7�|aXқo�&���ɸ�lجX��D��c^lg.�������x��DΑ�.�׀�E�3[�Y$dRǱ�*�4�/�g��m����F� �#�}��v���Ʀ~Qq�7:���u��oG��.��g��ۺϝ�u�����`0v�Us�F�
Ƀ0�o#�����^����(����3��*�,��I��/Gx�L~l�����Ck�R�!ũ�)C�L{��/�������ɥ+��s�A���e�y���Zz�eMY��=���Qʃ4۹^��'<!�:So
jv�v�g��F�b6���>$~�I>|%B��8�_�[b�]��_�o��6����Q'NnA�t ���VR�sb;B^����2;�O��o�v뱳a�W	E�8�8���$N�����]���"�|�4���ӹo`�#(�x��
Y�,ା�B0p�`Ț�肷�`DN.Ȣ|b�n �H�U�G�P�P��%���$Ƅz9=�����R���H�De�)A@����D�S
o�����F�����^@{Z�5��̬^��I�}�_l#_�Җb�M��M�0/���f��~G�f99�%2"�*��]��+]=?[m�z�݆|,o'��G��9��KI;�bQ�os<Q�},>cq��w߃Jh��C��$#:�������`�O<�0ϲ7}�t�w�cǎ�R�m晎p?��Δ׵���'��;t���Q&�O�Ob>�f~��o�F��Ȫ��,�^j���.1��R�4K�K�r��}~�|�he�`�h}|�6��$��=nĞ+݂(��/�~ݷ���@�4So�-?T�Ѹl����� �j��	�&�\�0���dA^$?�p�+�"����4\ �j�}��0�%�Z��G���/�'��iN�gr�g��y[��m'S�
��k^#����HϻJAd�+���k`��$EO�G��k>�[���j���l%��i�t����^=���ywf&G#�p�/<~���u�:c�|~�ܠ0=<��>A�G�ըrVb^�ؔ��r�R��n~��h!�8)B+��H�j�͸8����P������<"w�����@k�h�_��M���8AN%[��,�S�&��i���J��;��*�������[�qE-�ث�XL<�v��\�3p�P�·�����밌$��� QI��m���[oF��x��M��]��2.���֖>^Q���0�<�V�MNM35���'SBt��ϛBIc����q[�j�H�G���|��s��X��GhF��ٍ��Y��Z����[�`���y/���7���^�uN��_h^P���_N l�ߛ��w��`R���R�Ʌl�X�N��kW�d鰩4?r`��(�[��Ղ�mZ �e���S*|��iJ�8�o�5f)�[ǋ�e�/j���:V5t��5�A��G���qP~�E�Q_lA���`�b'�������oZ�ׅ�a�u����ib���uw�!�z�S*q�Q�Q�p���V����^����'6ޭ�3�j�L���́Ac�W����q�ޭ�Ћ�����`P��[�o��h��0�M�����x4f���]�z�_����tb�df�.�B�B�4��v �1S�R���Z�͗p�vh�a_"��-<��w^�>�K>�`����M��wn���.�|3�3�٣���.�Ѝ���9GBz�;&�]%`?'aq7�wB1=U"%-��q*3~(\��(	dN�^L�5kp˒�$J��o2alm/P��O�j��]̢�d.ܔƿ�^Ld$5�bӋø��٢G�؆�C=`�JVѽn�ˮ�/�����ɥ�b:I�����K�C�����I#��3����)e�E��+�?��Rtd\ض�1�}�u���syf���>�*&�L���F���k�SI�jXoW8��N��kC����]~d��&�V{gq�e��q���ecy��t��.θ�D+8��C"NT���i�'����z;O����H��z��WJ�T�\w���H���?	����N{�N�]M��������C�\0lBhl�?E3ᔔ�������H�2�ÝCK[�C^�P_��%"q�hpd�	�L\-��&�w`����F�U�:��{r���=o��c!�l�r+����כ���ɞb���!xm���B7�~�ɟK���pk,�� |�恭��ᯚ�&Tx������G�T�\Aƃ�Iҟ\���S	U���t�]��
d>m�p��]�(��垷3=J��,��`�X�A.�\ݪY����΍x�y�nҼ�V�JkI���ie�c�'zk�{����}О���-��{&�b�F�C�����**,��'���	�Z�c���7�0��C�)���8UH_]��������d���'����ez�c��7"����}�{�2IO�������C5s�Kf��4��"wq`F�1�D��:�I��`�5�spj��y�T�2�*�@��) �t���EX��B��?Vq������j���tb�}���ɻ���x���C��C�#n�G�;5�a|�m�Č����4�[<~ƽ���J&��{L������Bi�����������rP��J�����l�$0�X|� �Ox��U`4[�B��x����	��!�0��d�L�,k�������g_v���Hw�z�
w.y����3���!��";����'�����MVH�n�rT]b��87?H\_;{�7����}�g�s~��@u�(��5�t���sG�L���E��Tk١�md��n-wʹ��E���$n~�jE��.�1V�炑�\�$\���D��?-���Z*i��{C7�ֲs�)"�َ�����Vg���V�-	9n����/��}�W��:K? C<��yB	h�I�C��w��B�����zTfƌE�Y�\WAU��-Y6�d�����ũ����&W���:��qɃ�����v��T�-o7�����)���(l��c������w� J�t��U�~���\�ۨq��L�Jyd*�b>�>ԛ���qxaսfs����}CLߕ[j7���ɔ��ʵ��b��2=�F�G���L�g�V6�^g�b2����&ccam3V	b�M�<���RҬM��
5ٙ����4]�� F��1�Ɩ��wl՘i�|[�p3�9�
;G�>���=�ךwOi!��5�-�B�!ɳ����3Z�����i���}��늖�����9���@�^j�wȫ>���ą���k�1�{���`K�o��.%6�?�%�xj����7��n� ��.c3Mͺ|��"�m����KT�s,�)因}�a�U*��=�r҅���x=M8��6a=����}�nd1�Ū��u�Zb9͎�mP��|@��	��Ӌ�빍�3�&�����3�+_��V��9	c��U��N�5��M?%��qe�Q:`ܱDX��8���4XTL*�z��T��u��1�:�<:��}/�b'��F��=C��
#��^$��R5���䢇\9���`kՋ����n��5P�ɪd�s`Pn0��X������@��Y�$��6������]�-���)�ÊsEV[-&x/��V�m�
��J���2]�8��옘��N�_�%�$H�)��M^0)� �P�dzљ��0���{��'[ul'9�*#5�㮪M�s�"�0�{�B9��QW_�	Q�2��/ ��E�'�R�2ֺ�3mܛ<bz��$�x)Kp�E�G�*��V�(jO<vp2ٛmG	*�����$3Ҋui�H'��9��۸¬��~X�$�Ԉ;����/ef�j�a�EA���b�*�l�X�&�ݒ��*�l]�C�e}u4]n&�>f�!_:��,O��5��#�@�T�[�M�Vasמi��=1�6��;��fu7��[r�}��_��pSO�_�w�Kx���j5���6�{�
<����؍���%����#$'���B��Z{�)	d�p\Xkc��0����=A�F�$�4F�d�A0��"�rӄK���u���kXr*~:�C�Wt�k-Ě�Ϋ��L��g'�%��}e��29S	1i��;|_��X�v�˟4��潫����sk5�^��,福�w_����e�sq%�X���yQ@��؏jf��f��K�-y?|�M��:92�$I|�����sُ&��	g�`��sR���C����qe�p`%|[�����a�j��26�~�G�4��K�62~�=�f.kHv��(MNX���xЈ^A�e{�ϙ�o3ePt�Q��D���+�L���߆�v�NW��/n��b鏉Ғ�+AСޮ͟i�|R�D����j��	��w�j�zy/���|��:f�5<�\�4AZ�%<��hNh&�=#L�AoF<��n�#�m�xU:���f�>�ac��K��c�C�h������i8�]�3���_���<=���ټ)l/�9�5��Z�n�Nv�?�O���Z�$����d��_N�~�(�	!���b�T�J���[�����T1�O>*��d>���U!fi��$.��~�}�gf�j��I�eoz᱑��'��C���1�L��`��?�U��VO��rS��Q��
߂�ˆ���*~J�=�#�a���N�?�z`f{�m/S�'�ez�P^uR��}�]��=�G�Y�3W��͘���}Rw�f�_�%\+�8Q�tG{��]����/G��K��p�kpc�^�'9�T��I��5Qiv�ri�)����<�ń�3*���5��M�?	���"�g���/����	p��7�2Av/7��X�9�Y�H4]|�ȅ��W����j]� )C��Ɔ淙��*xK*��~`��S7뇕�>�C����Ǜ���kcY%��2��\O5��+�s�'���g9�Y79��W��xε�\lx���4�,��N�~��D�MGpirRי�t2�8ݬ<��!3�����C��U#*e�]|�!����Mx�14�K��;�<!���8U;��Ӕ�
�a�A����90|���!�eʑ��v��$�O��ܟ4S�����q:��$F=���朊��Ť �b�N�S2R%�n���V%HS���������@�j�N��݊�-�����z��ĝ�yI��o��×i&-A��Nk�>��E�'������n�������#/D��]_�S�^QV��Y�mk��ڴ.�����t�n
}�C�m�jm]NS?[�6kb@[|:K�#��.�[��䤌���07��j9T�� �IUj��˲R��XlzD抶���Gfͧ���W��oE�{sq��w��e��HU(u�|�C@�6~��~lSp�21���6���"ЭQ@�M}�W�R���)���uJ}�}lW\��e���ȱ�贈s�tp(�4�m�MA��0>������;1�t�s�y&2_L���񢀅�/��ms�*1
�%����":\E-���ei��?\�^~�2�@�K������⧛�Z��>���׿�,mS��j�D`c���P�,��`'g���.��I��xu�����"E_cX3xL�e�]��m�����,�!�⍬8�A���ۇ�Y�S1�.��{\�+r�����q��΂��8��N>����}c #��E'Ot�%��]�7�)}�+6ν>���_���8�O��,�c�c���,��ʓ�=�9=~	kc���ɟk���X�K=�:�SV�q�</���}���t�����ں$C�~���i�b��hM9R�'sY��p8L��j�X+�U��8���s�.��b�-$�^&Ie��W����EZ)J�D��0�� ׾�E>����u����������GN�oI{��c6Է�]�׿��:�Tr�f���ۤ�F��BA-��^����X���zc~��5A���!�I�+�:���!���7��so��5xnCצcw�Q��KU�,��_ս��/O�T��ƌk�,j��m#�&��.K'$<r]���4� �3s�)���$��4�ʺ������^��ǳBc�������"�C�yC�)�&[��8]
�X��&�=�d?�ް��)-l�¬��@�U��&�*�D5�I��%6��5~�{x�� �Kr�a�9Ba�H48��J��������sK��������¹�;ᩐ��ڟ�� ���é�];�������^h��3�K����w�'a�~!)}v]�=� ���'i��?)�c����}�E�a�v��1K0)jU��Bu���g�~��a���%G��	���(1#�;�_���b)f�)C&jӣr�SF�f�I��=Zkԛ$���Uh1�C��X}i�EQ�u���v���v4J����]��׋�D��RW����N�Y	�KF\��\�{�ޙ+WՖP���7�҈x�fRJm���Ls4F�YU�З:QsH]���D��*��h��o~fzB�_e���~���1��M`"�i𛅼�:���mmo�c*ӭ��tn����LV�d��
�vU�~���}�ռ2I"X���81iÀ':���~��w>d=�!��ȵOW���Ocn�Ӓd;N�$�!M�U 7ܧL��$K�5���#X���Ц�Nj2�s���1QD|R������b�jD�[�Ӏ�ԋ�rKO�.����o��0�h̓nΡ����=�y�nΤ(T�u-A�9^��V?AB���A��7�d[�i�W"aqAV��Q��c9��SK�&��"q�IA���:2�p�o���"�e�'8�������\qW�mg�Y������;{�s����L�,�h���e^�{s�����S�Z��5�[�{z�<-q��R���C���pt&뽼���H�����ݏ&�����[��x������R�T�����(Sx-f���C��+�����^oSS����>����RC�#ѹV�ǖw�{��8�>�4�S<g��Pw�'~�����7��V�j�x̸�5�$��p\|@��{�)����ޟ�e��&ʳ�ɾ�|����ߌ�kI�#����1,|6P�M�$$��/�\@�q�@V�"c��,���n����Z#e�~�wn���bb�Ug�p�^wL�"{e��!ܧW>--�-ci�#�.��3�l��iW��ë���̖�=}/X��:�L���Jn�eM�k>�k�^�^����>J�#�jU�(_�"����b��/}�}����T�H*yͷ_�r�}��+�q��3���$��sBI7w��9�t�U&�nV�����-�G�Q��y��~:����2�*\�cАL�~�<� r�����"�ʷ����}ƹ4�we��qdv�,a�(��xc�\�ǚ�����'�_����ౘ]���a���v�f�L����.�QCzn˦�}����D�:�� W+�J��3M��"�Z�4��m��֜*{(iprT� �Oai�a�_Qz�b����XGP�[/�ȗ�7�>z��^:{����=}����-�ӿ��*0����f{h�����U߯W�)y2���L��Ԫ_4�m�S��*���Y��2q?���Q�]�CuGڷ?�%�cE��@Շ��6��0�թ�r'���e@�ft�a8���3�������ǞΌCt�:����[K��J���1	g?��G���Ξ��4�M�2�wB>?�����їo��׬	Z�Hi��T�4Q�!Z��G"�Є�3~M��w�M�X�Ȓ��4q������k�z뛘��k�j|}8�q342�R��.��hi�ԛ��"�ϳb�>:��u��-wf2�Pdc)��A�*����pē��p����r��+�!X,�ߦ�m�2���o�-���Q���^z��=\� ه�t���8���i����"��JQ���b���03Q+sdj��M�G�	���Cy�"������У�~�����j�U4r�{+v*����)�������Ӈ��k��T��F�C�}[����l�Ƭ��?"������o�S^V�V��؂���%���d�gdsI��ƞ�D�GH�L����)Q��EiY��cF3D-S3��"g���){��3o��y"�}���5���5��*�9�-��3�6�@T<{G��E�WG�M��Y�՜ �n����x���;�&�ִ��3�[���jXU/���+� ��V��˹ry�C\�43����=f����}/�kK�G	#�s5�wm�c�\⩦[�&�r���YSWLLL~�ڭ����G�/��:l��:�-�}}}ݦ��/
Og1��<S��U�M�˳���FL�N��wyRzY|��!u�  g[`��j���9I�\�<�ی�D1U�M+���g:�"ه��o�,�NQ��i��p�5�Eo�i�ܞ�j��\���:�	{��c��.h��W���N�ϗ�s��+�����Ѧ���~��L��Dh���D�3M��:�|J�a�3������)���vsH�f��.�.�)�F��]�fk�����������2ٙ<'<'<�����Pv�i��H4�v��o2G�o�)b1�e�۠#�sS8�'�A]E��N �Z-��1���j����{JqM�Hr�P�ܼ��o<�S�^�b��f�T�n�]r�+aT?-}
ae^j�A�8�E���_��3�+�J�b�n� mf[+Xwv>_���"\���z&�Ũ��wg�.�(��7Ճ	�`7�h��gxy�.��0��-����غ��_�h�`~���gވ�A�B�/ٞ��kK���Yѭ�lt|]�B�7���8C[�\y����G���mO�-�j �(EQ���&�l�9"@�k����ђj�ID�%$�g*+����IH�e�0�p#�y����{+!�:�!����YGL����>χ���|ـ�ڟ�_�؟��+���ʺ!����<�{M�Ԝ/b�#��ǫ��͖�ծ�y.�16��Z���;���~��U�r���%�'�O���]�]�۴��9��~�^ L��eF�R���6_V���C�ĸ�x-h�P�9"G�� }CnNX�K�Xf@�A���@��4k-i�P��m�fm[�mZ	�i19'�g�����hV�.�nސKj0;�=ǒ�R�����@�]��bsjhk���n=�ڂ���A�і�����K��zA˴]��Y���Ɏ��U��}|���pon��g����K�������*��0�!��EH�x�g\�v�g���-JO�#�6��	��p>�D����/���M�`H�/M�qzz���I��RRbr͆������x9�d�wr���M�IW	�)�ul�f��e�ުf�T	�̴�V�U"!oW��M�¶v�"ސ��U»Fp5m�&)���l�i���3!_7�����M�ש���q�6�J��n	�*�t�>�2:��a^<�xGG@$��i��:�g�:�<\�ļJ%4+b�!i� �
�(�{������a��[o~y"��Kj�Z�'A<�+���
?]�Y�𽪔��5ܴc��nv9�.֏����|�}F�e��s�B,Nb�����I��G�g���3���۟ [���q�	�m
�k�'���Yc����P-&
�X9�j>@���tֹ�g�	�z]�}�u��qR�휱/�T�*v�/�X�qs�]HD��em
fJ��v������eX#��-�<��i	׳o��̺h�m{%��|���G�1y�z�6O����64
�u��B��W$�|��/��,�y���Na��c�>���ܐ��,�y`�aﭗ��I��r�	z�M��
|� ��Q���O�C���vE��i!�(ۚ��r5�ߙ�te ���!WJ!���E�w�&�C�!�]*���^H�!P�fw)������y�$ɵ/o :LN\\�x5�Yz ;�:��f���T�B����͟$^>�-׎�x�)(X>2�΄i �WZ|�.G�ƵJB������_��k�����b��t�&;(h��%�md�᪑�f&���}p`��^�`��(ȹΫ@�͈�blL�#�^qX�^4���p�_uT����f�r���g�Y.P�|��(��o\i�f��l�9��㳲i�Ȇ|�F�0݀������/L�"��uL������n�4�Y�m�q��M�%�������0�HH���1XS��bcm�����.�٬6���n����*�.����$�'p.V�,�K����؈���2գ���۩���ਜ��Z�U���I��mYP������yX-�P�*��r;O�(K'}�\��&�j	ff���y:�WU�ۑ;��B��.���w��%��x��r����&����n�
X�\��x�HQ����K�/]��
7|�v��uzq�J�o��3��/֌��_�Y,+�ZX���� ������zZ`5�t��a-Ph�5���b�C}Cp]��Ǧ��w
򱟪�+���JK

`$��\����׻u<�����j��@�A������ִ��[�y~�a@��\�vqN�
W�tм�N^�`\S(k��S���	�(�*s��2&�Ps�S^���p�4C?{Ws��6��@z�'�1*2���������⦚���G�������őx���E���������g�Ө׍��l1(M��)��9��d�s����ؼ�$�׹�9&�tWf��YYU1�����B�"�C����
z칥ˠ���Y1+��E��z�Ɨ�*޴"�!�����x ��i��H����^</pF!_�H/���d�Óq-3�����IX�*� �n��u������]N4Ĝ��Z�s�A�v�*�����﹮����pVmB��5u��N���@�����'�^Z�W�V�.�׾YW�/���;��/�������}�-���	�0� ���c<���6����ĭh��Mq�D��q%@*Q]�n�[NJb*{����K7���2F����-�N��4�8
w�0������� 8��1�^��LRx:������%�S�l��>�7�����Z�ә�N��s{��&������[�B��K�Wҵ�b�u��6��A�V����r��ό�~ϧd��Uhf':�����hֱ�ģ9���j^5TGh*Ubc1�t=�ekU�1l
	��"�Њ�"�l� �R���1v�;�I,-���3܉I�D�<�?�i��6v��=�g��4�˞��<�U+k,Sw��t��J���F�>Bee쟥��Ӷ'c)��	�~�b)V�[�ˮ �d�����Pd��Sz&ER�;^�����P��I���+��z��i��Rk]�Uj���/��e9������G;oy�6\��YDE�T�xo@�V;��]l��Hv`TZ�
���,��%3#v���.K���?/I�<�r�ү���&d�؄�}m�ؐS������3�9�ͭ��~;��*zl�.S��	J���	�}/Ɣ�D��{ �`��0�M�G&�n�Q�����BTM����u�uGۤ����6{���i�n�0���8v�3n2з;��vz�S���+S�$�d�K(5�7�coS�q�"�P�Aw?4��ń�u'�恤�kx�&I(� ������\�:[.5�r��H�1�[��P��y3�E6{���;t��"�\ప�!��%x�(��P�6 2}�-���̳��g�A7}�݅�����%�/��ϑTU�مJьjC�/��7l�f4�=���VxZ�GnתF�y_�vfٕ�)�E?
����4���-���
�нv����	 ;��i�=Q��R��s �ȧ�%�Ɍ�in�����U��Yjv��x��vA_j�?����G�H��)`#l�*-ZN/�"� ��f��4�8�ws��*1�4���h8���\��l�,*:/�.�!�^�eWq`7��Ir���`8r>� /?ͮ�|4�r��~�L�?b���A�|����~�6v�{@���Uf?F���P!��	4<-ݎt�U��Ջblvv���K�bj�H�%y����WTϤ�!a��l�k�U��ѡú)��a|.��G2��!F��/|-y�L�y�\<�a��Z��q:U�����M@�7��$t��FhLҧѶd���O�Fa)c{	��$a�ײ�&���n�^�*�uX��}2)��q!3�C�Ko�+?9{��;�7pS$�
yn/��ʈj����I3R����t�n������/ .��Wח���c/��~��~]�]��v@�ލ5|	ZͳЯ=�ʹ"���C���x�;b��`#^8���0T!ۚ��"����HVW���T�k��1�Ě)�,��s�jf�Pހ8�н����j�!gp�`7�1oM��<n�O�û���M��}~�H/*o�΀������6Ig���N����
�o�~Ykˢ�?Ϭ�X��x����y`�^H�)�2ogG8�@?��$���T��3����	vkG��'��\9Oi*����0)o�ܹ�N��J7�P���Y���.*���/�@�H�K�һ�Ҁ�z�-ro2�R���0�O\��黁4?��[5�/�����w&�k�<�P�a3X�]���|��mU��s�{/�j߿S�:��y��k�����:���W9��Վ;�i6��,�r�����Tq�רͪ��12[��D+U��U͕�n�a���V��P�i�li(�uCKb�����W���Ɗ; 7�����X�ͩ �l�L�-<�ǑVL��v��$y9�����B���փR��:±؝�-�\�	�ጱFl_Y��6v�o�SÚ�B(9CN���z�dY�=��i�����澝�r��R��k�I��Id|�54��Y�����+z��G��~J-�̹7D
���~_�����~��ö��KJ�x�S��T�#et�y�YVr�r��5���=)���
���Ӥ�-�^��&�3�U�}��z���Aa��\ۭ\�k�t�G'^���z?9eӍpn1��?����j��,�|?���M�;���{���x5Ab�J��fS=�]:��o夥�<SB/z:C^'�J���j�_dg�� ��;���^Z�A�RX��	���-������]~��ć��E:�jY�qkUse����C�8��i��g,jB ��S3y(S����|b�������d�%�s��q���M�hr���W��gV��W��6�P\oS֧e�2p3OOa��c��H��U�()fB��*���~������ZD�ԠW�\�#�a�/�D{�C�=R��F��ۮ_&pd��̀�U����eP	�2ol�Nďa!�;2X��W�@1�q>+���G��5ª�K�i��G���������xt~��q{rM;7=hm���?������N�5�z=����][�N,�ù1}�м@�+���N>;�;R��ǲIh����W�o�V����|�ᕩo}yoYߚ��=��G3֚��h�^��=�7�͋��@U`k�����nsq[t�>w���Cgdm���q��E���{_�Α�V��v��r�Y���PG�4��3È���J!.��ᘘ1���;#�����D��$_EO �$C�C������5�x�iC�i�4�F��F&p>�}CI��������צo�`�+��|-�1�ƶMo�>�_3��	<�$Ջ���Y��9��zא�o�]W�j�T3	�Y9"��Q���'��Ih.W[��K�#ޓY�,�e����$�f�^w�8	�6,F2�f���o}>���`�*։|5f�N���n;��+ ���U��ٰ�䥂Qq�*����m�f���Smӥ���,����y�3rwĿ�0�]��ʜ	J":/<�Gp�݉#	oKUna��L���2&1�[��,ɫ�z�$���ق{|s 4^����I�r-�6z�LL�1�"/o��*�ᎯA�VQ�S�d��hG���/\����=�/���� ����J0������t�u*{�<�p��> ��u� ��^���F�&�aSK��;�ҫ��Q̡K�=`�>����t�	���o��S��}R��J��,�z4����o1,9�w����i������Д`/b�JR�J%�Ë��?�߁J�^��ʬ�k����ܸ��g�3^�������f�I��rl��	��H�|#r��/�O��-wNs���O'�O��w�.|���Ψ�Z]����/���x��E��222���9�)r�����5Ơkm�|��I��(��N�I�k�Ņy#h�W��0�N�^��=<V�;�{���VǕEW��}�֑0Zd�t��#v[��=�<�.6Yފ�&�}+�-F�˔;�M��hVƽʦs�(V�=i:�Y�3g*�ob��p{9���>kf�^�EQ�ؙ=�Q6H��6UfP�`"��I�[G����͈h��ޛ�D�	<\�+ RO�q��`���D�Si`�tτj�Ye�Qbe������	�N*Z����L��1,����@J�1�E�yĪ�-��.l�������kH�˞��(]6ϼ�������8E�]��דx%��j-��-�gL�����|�L-���~e �������:��[�J*Z���d�Y ����O^\C���
�䟤>O�ߍ��Y1�փLM����z�������^�t�Ы`�I!�RCmw:������ley3�DM���]�2?�х0Q�=���w-X��/��>�1m�9�kI�����p�<��v��A��=mڰ��z�8%9U�6�o�^�����Sr�$��lxEn�]N�.��C�$�����l���"�~:DcI�B��|_�`{�=_et�-�n���>��m��Ħ��7qH�d��r�'�i��p563U�x�/*f��(���Saz�]x�Ό���P�%�We�v:�����K��j��=�(6b�:�����^"P�mo?���_���g~�F�n�6��ɑ�	�T|�:�==��6p�|�*dh_������c���M�햖�)�����5��C�W�㰮�O��x��;�܊O������*j�j��~�W��`ǔ�V��=A�<Wa�Zt�=�=F� ���k5��S8c�nC�v����mDh�>T������״�	�aPM��Z���	��.��[M�5e_2a{�`r+'/*����/����W���KΟ������][�&�>����D:C�(�^),'���!�S`���&-�/X�sX�\��akH��ˠ�/?l
�M�g�� �N[:%���ٟx�^�؞�'u&O5�0��-�͖�*��VSr��%i��M�o8Bͼ��ߓTr���**m(ܧ\q��l���0|�$�~e�&x{Ns����-�w�h���3K&�LpF)��;zq?#�$�*�g��b<w�}p�PIQ���2�E�+�M#8��l �5݈\�;C��E͊��4:��}��M�%��X����s���������" �-:��/<,쑑{�Ϭ��q��H����b��ߗM�ќ��k.7��l[]�r�!M�4������^S}��X�ʜ_U=i��Bv�!B�ݽ�Օ��fxJŏ����AI5�!{zBYD)�^�a�C��gY����b��ˡ��^Z@^S@��d�.�}:�j��6x��*�k�F=hs%����	@��K�i0{��"�
�����^/��u#����`����^_�"�[�����[/5��fd�.ȑ�w5������ɠ��s`��C7J)�%�rJ,͌0v�����R�~�����;�?HO�&��{Xu�qŸ`W�m����#ɦs�2��Ԣ�t�Ԝ0��	JP�WO�l���=��X+��r����q��J)�-�q�j�A���
-^�K�k��毃�߄l�̄�'K/k�z����0�=jn����&��A�_nh������	ËG��I�ƹ�s�Y�I~�������Eۦ��[����e����8	#��>����S��2�4ٺ�@��=�4ܥr!��Q�E�l�ߺCNU3��}x[1hV�U����� �O��ۣ�>F��	ᯂ�o��o_�6��&�F�9mO��H�R�˫a*.������p2�Gs�~� V�U.�7<=IE*�o�%�]��~�fb�W�`��'օ���)��&��w����;?��]6=6�xXib��SK?ߋ���ru:c��s�/��S�<��S���۞�+?���%|'�������U��^�Ff�y;ӳ������^l��jE����S�7'��/��x���}ʳ�o���=�j�uwi��	��eA]�W��V��?�8�������O�>ϤRV����z��ɥ��/B�l�?|�+�|��s��]�t���U�()���λ��/w�jf���v��KgO
��3gjf5���&e�_ ����3���ߤ��(�W35���/��G�yK�|�ڳ��3^P���Q��������_�/?k~�A�s�hzd"x{G�㣇1wn�ϳ�~�x3��ɶw����?o���w�㋻;F�( �\�t���ᙧ�c�@�����҇���%_�>f�t�sY�� PK   �cW��cH�1 &7 /   images/4657de38-a294-4f46-8901-aa5929bd88a8.png�{�_���J�H)ҵt)H�ҍ4K���(��(�% ]�҈ KI-ݹ4�_��{�p�|���e�93���̜����H�O�  ��^�� А��K\��_��RL �e���J��L��.6�N� �OFb2���e�d�/�^����w#��ph�=P�ɱ��6���G��d&?r�^V3M�Dr�Z��~�p5|ww�-�?����y�	x0 (�i0+E�Fz|]F��n�as<�9�@{�)��"��{������ ���3P�������eR�p ��@���a� ��!�@���yy��X�D5��yN �/!�@�M.�y���6`�O"K��O^-���]�H�2�Ut��pt�*Z��ay���R�G������o�}���>�<���U�|U�W/�|�N7�Ĥ^��7��,��4@�[tSߢ��$�%�`&�N�f��%�h�5w*�X'��x��ʚ�"�$%_�ؠk���61��ض���>�c\idv2�@Wcޖ�NF�#R	d��tA���[9���Ӧۏ��o���H��D�Y�5��<o�� b6�2f���)��2OߑV����8jo�k�nMN}�H'����G4����o_���cri��&�E���j��!k��̫�x��|�~l��h�G~�-�.��^�|���O�R��zu�rci r��`�_�ڿ������x�q����M�q�V����}0�`�ɲDb�1~&d9�2�'�(�t��I�
�X���x��`�>ծ�J)��>Bbjq�-��]���w�LV�d5�q�k8�e�5� �򖯰�"&e
4�_�!Cvr�r�G|��a�G���n�R+�x�B���VE4:��K����H��n��+�?�s�p��Rs] ާ��w�9�Z��>��������K�5^	ݛ0��<1�z-�_v�i�
sS�8��b��o�׎p��$nal�y�_
7QJF߆�C���D)ɣ���wSX��ե��D�4�B�?hO�4�
�:=S����0R��{dg�+P-��A�qu���e�A�����!pNQ�2���ju�����.�Av�t0#�&^7�������̴���)�g/t�p���(��1	?�!c$]����=�ҋ~�7q�q��~Jٽ%o	�#$��?�d?`�~����@����EY�5�&K[�Q�W���:5�+��t��y*�t^ۯ@USX׆��5\�[O��_�7R9'MS�5�k�G�/~����t�u���i�k���x�Q�$�D�NӫrkB��ͫՑ�4 KrV���.8�<U��J+I�7�"��Ս;�c��X����R�����q�������:#�lzG�JC�-$��/t#8.(b/�(5)�h`74aXV���79BxIxN}M�*��!r4��p�_(0��P�c�Q̫5���q�O���ڧ���L�*�z��`�J�*Ė�
/3�	D�՝a�Y_BN���T���	i�hɈg	#bN�mh�DJD��Uym���\�yo�-Ȭj&�ά5�?��.�~��x>Pֽ+:�a�e�6~]��������['�Fa��K���-�#Qk�!�Y�p��T�B�T�������Mw/ۂM�ZĐ����l �����g�\�6�>A�� 5��uE��0ԓBl�}�-Otl��k�tb��`gnIb�r��RM�:Cߪ����p�P�.�~�74�Ճ�6k���o��3�=̟ɚQ碛�3l�)b.~;u�qVg�����o��uXq�`�^�31]���U��_�u�	���jCkcm�,	�
LԸ&���ٽ���@O�� �������3�|��5�̔��P�cm)r�����cq�3�{93��iV�E����E"���𯼸���s%��Ȏ��#̏^�E�0n�7>>�H0Hx^�e(��irA��RC�[���q����-�!�����t�+���h�l�;�L�;$d;�����/Ô��S���-/{�x���p���|�Z>�p^��i!�=�N{�k����w������p��v�B���"��<���_�v~����_�w�Y��
R�Q�w���A
�7�r(���y�} �&��(i�F~����}땕��ە�d�n�Q╛�銕���dc3�j�϶LV������� "i�Ǭ��ҕ�8��3TJ���bg��W�*�At�ò�:��Yf���� ���㥈K�f��ֺ}�Ҡw�յӹ>��z2پ	�ٱ�1�݋݊۷�:]V���ήU�O��>V�l�j8�����/�����4�G�L�z?�\P�c�e��-��q���x�&z����x�p,Y�o��,4Ӕx���J<B�ϐWw-����/�^�{]^6V� ������!�H/n//�:�o��ga�M���*ao:���I]_�׺x�{2I!��^e�GG��v��i9�j�CO����*�e�g�4�nvou.�J�K3\�}
�gZj�l�l��ٳ�~���ދ#=f�y��Z������{f�5Lܚݏ��:�m:�MeVd_mדg�3�D���s��3���A�J�M���6��&b^Ի�)�	�?�����T�{v��Y�N>�	�C�D�wP����E�u��xk[�T��D�t��"��� [++�d��d}P��H��F�/ϥ��i,�Û���X=��ػ�������۩�)+���	����f�����9~�}��>Y;̗��@�#�������^ъ�ʊ,+Ad?'����F� ؉�1�����1ӮqR��}j6��PYL����.�RaY}��$�1�vb�|W�۫�/o�����s�a@�ky6����m����� �c��6��s  ��B�����N�[]��63�ML�C��T�@��p�N�ȫ�w"{�7�pMB�{261�m�����c��QR?P�e�щ;�KenC՝�z-�>����4N�����L|�Ɇ�Hm�����-�����S������ˢȕ����<5�}{:ry�=�� ��(� "!Qs�KGcꞩ3O��w�F�K��muw_�&�f.����kk�'��ttDi:�Fa([����f�fi�7�w7S����..w(������������֖��;wЎx�jP�3q�6���)9�'��9�6��3���ӊsWT�Ǩ�����'uwwK]��}���~=��E��cvc6�D���ξ;!�~���ؖ�ѣ6�����[��D�z��Ukk�lss����I�Q�x���;��]/��R�S��*O�վ��v�	8�幹`��sP���*���d�4�L�������u9�iۊZ8j�>{cv��hvRRי�u���Z!Ϧ�蹻`�~�}5�HGC�7����ypp����4� &������E&V�.�Y%�}~��wm��]�fR�_
����	+VV j���u��qvff�]l|�-ͳ�zL��Y����Lf�q~�3&�0V_O�����@Ou�r��vd۶S�氬5)]���[���T�T^���� �wU�������%�(���(��f�� n��66
	
�~	�Q�xu�NYg�	�o��og��""�D��,�q����m P����ty����J%[�p�)��ؼ����Ԑ�9լ&���e���)��<���m�p��}�� �����i��͉Ā}���<蔾�D,����0�;9n�g_n��(.���ϩn�K$�Ǌ��ϯo?��k��ON>�y�:yC��>&qp����QQ^~��x�x��5�ZCG���T,b����j�S��6N?���)��s;^�pէ��I�b�g�p �|�v~9j����H1m4Vac�w���r9���Qu�Ow�SwW.������P3����j� +o۞�G�pґ�ڒ6���z��i0U�����ӿ&D)�vQ[���� x#�N+�Ҿ��s���t�玷�$w�e�B�� ������� �!F�f�גeO�`I�E�Rj�f	
>F!g��T:���9�RM��L�Vrq��0�0�ޯ��O�q;IѼ(������V�>�Bq6��y��g�����<-zܣ��h�f:]ϯ�Ӭϖ��y�o����я�D��ֈ=E��
G�	Yv�5q��M<66���0d���ȁv$���A-��q�d���!x��TOeX�|�w���n��%'����o�4������8!�"s=6�43�K`sSK��1��"ΤS��w듂:";��k��kf�Me;�R��_?T����[HV�766UxZO� sW�`t$��}q�_��L���,�4����_� 9�o����3�������I��[�+��=��8,!`���>^Ǵ�E0�����)�i����£������±�t�'��	��He��|ѣ	�햿'�*�{�����Y�]Y�[��O�"��w�(s�=&��w0�@���[=hL�Zz�Z�n���l��~�^N�h�I�������v43Ә�ɻ��9���?�9��jl�khi���Z��W(�4�������pq��5E99�B��ԉ9C���J� Z���rͷ�iqFo�B�Q.s��.� ��:�К��"�5K�F�#�훃� {G��w�/�3GqH���4�W����99����08HVڿ��,$.\t�$�c�fG��W�pu�#�4��,B�Q�{w��$��^���vz�}hg�Q�qw{3D,$�"]�BV$XQY�,uw"��tP`8�P���} !��8������E�����u���a��<.R^��D���ߦ����'�M�����A���:��<-���3���v-��lfC��}�����d�Q���3;�o7������+(3�F(��k$���F���̊���ʾĝX�I~��N�:+�H�:!�b���	f����{���}� �~��C+b�J���A)��|F���)�A����ax��S�h�:{����F�`�B�D\�V�(�� �⯌5��0!!��`�㶱� >W��B��FP=BpR���8(��S�\ý0�����'��q��o���]b���-�$��RA>��ӵx�4u&�l1�A1)�I��S� (fk��Љe�Ϧ��^Ϳ�yy���!^�̜�������(1RB��}w+��M3^-�S��2p�Ry�kQۏ�à3�Ȟ588��8�����\1t�L�t�T��x�d���m��A	0}�M'ZWmX&��WݣI�(�.�ÃAk�,do��P!��]�رv��H��^�=C��[�ӚAq���sV���Tޖhoi�#/O�Ǳ����{���
$s�s�_W��p���/6�],�Xru�%�v���)n4�a�ⳑj��s������ۈ/(�яn��
Ǿ��������E,?�W)����9��=[Xƴu�$K!��2����v��A�����ѝ��cRu_<�":]�H����9���a���_5Ŧ��-8#�OY���;CRK2����|@{C�ʹ�a�s����ߊ�Lq\�>n�pz��9l���[�%�>臋,��8'`{��޳}g)�K.�w�@�l�K�s������郵�9��jGT�8}��;I��F��=��iB�tTn�x>=[;�r�P�f���!_?�>���d�lM�j�	���R�R �Sv��'@K��s��-��`����L�j��>�0�l��������&U�@f���W�Y�����Ր�:D�{���J̙��'~�j�~X'�D� ���[SfV�RO� iGZBF<����P�o�,�̽���P1���gfg#<��q�fi��j
3��C��葋|2#lQ^�jG��t���Bt=�^HЗ5�)�à� -m�����o�9bF�&�"��r��e&3u~_�G@�!��_�捺��n~���6��=+*�9�Ӈ�1��j�.S�l���鄺}�S\������e��*�tn΁ӄq���%��b�n�����V[m���d�F���uL%Z(7�ŭE�}�E�
	w�v���~�o�R�^�n����0!�<�m�z��ͱ�y��h�)���X�(eߟJ��n(T�s$.k��%��(���%'~�I�����̳�L��e��N~�֋�2��{�����@���v�
	����sn�����G�9��B@f�!ӻ+�p?̏9��lG�nK�+SY:�[�2�l����Ȝv[��A܄�R���~?���Q�~ ��x�H�$�N{��89l�x�}�˗�(.��H{`���o��@/��/g���ƪ�dp����I*,�%ad�_b��Q���ē?�Iں1��x����'7��P�q?�����fЭQ|��\���.�EN�Ԁ��'55~����1�a=q�?�K�s�8{�}���[���K)O�`m��W����\UE}�h�b҄E��%2y���9#''�j��z謢vu�:�~8dV���Ktr��k{���m▵�ց��$�� MՓ|~�(I����0"	=�� ��q��i�c��G�b��ə���IX���A�����e�����e�����rE�B�^#�m��e����l+j֏�@fd�/��>��T�-g�}�,��_�|B��PI`p�LR�yx�V�n�<چL2�-t����%�;�HJ� 4�:�[`���3+0y�{�a��N�yj��m��X�i8p~ݺ|N������M!c����[;U��ZB�q@���K�m�r-%�#2�TQ�����ނ��>
UY]�6i�fVyTk	?����Z�ʘi�WG�����dӦĎԍO��F��S^ɀ;�g�K�����ĉ��ivS�WV��s�p�d�%���䆳�����I���L�Q�K����ي�ɥ=C}V(d��}�p9�#���w2��]�巯�?X���ʷ�OB��xv+�tʗ�� M�y�diE����D$ْ�ɟwv�\B����!#`���D^<�g��I� )&]x豧�l�)Ht]E��?i�^g�(�k�*�_����݃�5	����y���>d��?J�_6�c}��K0��A�ؘ[�R8����L<u'�?ev�"j����Ve�W��[��	�4%|̇ߪ����j����zZ[�I���\w���$4k�������+�~��b1s�_j���-��3b��P,lo c����,�2�`n�=�Vn��"Y��V��Ɔa�A��Ȏd�h��
&oR�K<%F��W����i��s��Y����E61+<��&a�5/�r<������}�~�K��������W�; ��R�"��mM�
�먞��r��\,C�B���2�S=Z���?1��Dԁ<���ސK�ۜR8�Î�����Y���î��V��7������Gǐ��d�>�x7+Φ���g�N�9NAC(���s�],P�e�Z�^	�65�(�G~���u*���a��W�i��b3�pnґv���jW�v���f��HK�������(Y�A�w6y�u2��"��@Ӥ��'˹)/�	��`v+
����r,����Ue�(�U���B&21Qg���?���$#��̅�c��Ut>�{B#���:����¸q�X�D��>��ڷB�J@��<�po�i�d;�?�ㄭ�(�����.&�xu(����0�������騱667���%�N����eb҂���΂vޘ�,��ف'Cۦ⒭���<�/^M~GL��|m�<Z��짩s�/#+V^傸��@��|���`�]���&�u���C����*i���H��`�,��Y��wq�Xj�[�ǎp�EM��;RB`W�c?�a��OZ����~�ݫ}�������x����2= o�"�i(3�R2��aA��i.,̈�O5<f�ށ+�f�Ǡ`*zz�FUŘ]̈́�u����͘��b�s���,T]+��od�N�d�q듾�r!�w��Z&�5dō���~0�H�Y_B����X)'�e/�_�o���s�FƤɒ�װ������x�JCI<Gt�?>g�`��n�k���-6�m�z����;r�^5*'�ɖ�p��h�=�j�>c?�8�X�CC����t���&,�9�A؊�Z=�!���UV8B�/�!��ܮ��_Aը�}���j��jA���ٽ>�-�d`7�A�~�'�2��F�Z!Oh�½�Ս�3�1񼭩�6&98xED��3D�z�K�z,�Eda%=��g�3?O�UD����(�\�°����N���HrԒV�Ɍ$5�d����%\��um�Vi2���p����+B�bѧ���ڝb����O$��w7�G�>ʉ+��"���`�==��Q���ʷ�ɜ���HK�V5��#o,����c�4,Ӭ[����ɉG����MEF�݂/�k�in_M�#�qS.�6�4�?o ���~Ͳ�ۿL������r ���,4�o��6��Hz~�����bQ?�Y]���+}�Q�q���+P�����cz}}��R�?��G� n\���ڠ�?����{JD�GF��d�v;g\Q �Qw5���t=R��jw��m���Ӕ�ĩ�)���/��'(�$��?����ۨrZ]��INp��}1Rx����ʣ��}d���؃���w[G���\)H�k�����:Q�t���?��a)Nj������=��k��6�Lm�m��xf�5���F�)o<>��u.?`�W1N2wV=�Zݏ	T����.�WC��2Fb�-���n%�
�lߑ�z%�� ��ҏ=��:�LS�����^�/�O�?lw5�X���2��C���􋨜���7������gB2�F���F�i
R71�) �$�m�.!����f,��$�=:ʇ1�*�Kqxc��̺�u8���F0����F��(چ1��ۄ���h�佉$(��[�W�xU��oH5��GE�#��b��HSI�M;��O��q3�:+YH�������Y��h��t�Ź+����zF�=�14���eu�տ���$��{��;�Q	������A{��Dg(m��T��/�L�����1	i���V�|b̛�gУ)Ͻ�I��UV��@nMɞ�����?I3�sk�Yn�_��W
��v��ҍ6`����bo���Q2�rN��,�O㡜"%=�`��{�U� B�6P3��yP���^��-5?�"+� �X�CƢ!EZ�cp��LC�[�v�
g�`�?i���z��͖�K��I��95{1}��f(���c��ĸ�N`P�O�Go<dW{t�aΠ���a���M������r�,։W9�2�Bꐾ3�/��Ze�vs`�w6���a �����צcN_��	�d�o/����̞�u�7�nB�R�/s���
�fl�b8����{|t�J-���uy[l-sw�e�xCg��:�� !��kF"湳�
�0u=����z�� ܫ����A��J`�8�q��s����B3J?�҉R��qN]�I�D.-C�w��WB �&0IB�M��"sD��:�%Ф��c�'r�^�X~�������@YW:B�E�(@�T��`&����.(3�`@�ef�<%���ҍ����r�\#iDv� �s��o@����PY]U�X�y�kj���`:�fͥ7�[�E���!10�j�Vш� �>��)��8-l�k��
���"F�A���]p
=�Qۅ�=}s�+-��	�$uz������@ߗ��Z�/�:ՙ�-���G��5��w���e�zuKZ|��O�C��J�
��;�b0���'��D���Qv���L�o��<|QE������� {{Q�|zi�B��	�w�En���Bl��|�4�������Ğ�2_	�\^��p�Cߘ?�l}"sE�s�MG��b�m����̓�������_��\�I8�qa����������%���b�с���� +if��V��P�l�j��M�q��l^LE, 4�,F9p��=�WlE������>��V��eL��:�ں)8�#�-�^O����< ̏��鉵&4�a(��({���:�v��w���m�{��x>�XZ]�K�%���f���)��Rye�g���Y�'Н���&+���ӛ��	��}����0J�lt ��\c���_�pB�1�n���,׏���ZI>>���>"^+'�^��\�� Sӷ�%�c��1��z��E�H����4�`��8�	ao-�(gDrR27Zp�����;�m��GG�h�2ޖ�o9]��x���1|(�Y���Mxqj� ,3�{3��.w��]�W=��!��Ӭ��u�O����k�́������@�<�l:���ʞs���6��c{_���7@�Y���$<#5�>�F��爘f������ӈ�#�'�:�
2�.M�#��Z��Z��\����'D��^Z���L*"���Yqy������_�I�^����+���(ۗ��	�?um�p,�7!��0N(7�-:���7������M��Ⱥ/���⎿ c"���-�aՙ�tǺ�M�֒���"n2�?8�ě�5���ǁ�|97gfwg����̃��rg鹛-ޒD�ڤ��U]L8�fU_T�7rb�-.�1�h�؄+�����LM�@���6�Ϡ߃r�[.�!���=�s�� Y:ÔQz�l�ڱF���b�3!�N�!hv���֯��i6�#��{HF�����nϓ�6���!,i���C�f���k�+��Up��9���Jή^��T�.�d�'�E���� $4�m,��q:(��o�h����A0�I���m�E�y���*��3'Lg4P�p��Jl�����F�v�뵎��[W[_%�y������E&��@Qo���4�@?�����\���IF�R�Lj*���&�T���3����<$�s�j�@C[no��QԖ�VWSr�4�vq�-͗��m��tN�Ա���0���Ր��2^��E�IY]h�������:�66�h��q RV,���.�F#t�2y�H��~kw��[vܱkz�#�@������Gݢ�^�j���~,���v_�M�2��n r;��.�?�G���Ғ��,L���Q���B�,��\B�\At�qv?5���"Hݼ(b�}��Y�O�l�M���7���#K��$����S��R�Ⱥ��7"ݡ󴪊w���A5�����,��9�����v��_,����V��3�>���HT�Ǻ�IY�a?0��ծ���ցNrf^��E�N���69i~�
"���ⅿ9�������]Y0w�����J�ܾ5�-2u���>>�`�#�p�ko�y-���n���������h�9���F\s��+rV�^U�w�a���:�-T��w��3 ����3R1B������]ybRR�^r�8���ǁ7�6�&͓IY�{�ر��xW��3�� 0���}�{��c��M\�:���bQ���߱0���I::f��B�" �!D���m�p��dU� .+?�.̔ij��{���M�\�	h��r�Y�Q88
A�{d�6��gG��z��U
����n�f���c�������_��D<��qP���K�i��N�>�3k�GX�!Zs���C�Pl2�\����1g�oR:�f>�I8����
OAI���,�#�6��3R���?�i߳��O�e�G�䫨LY`�࿑��&�%����(�J�ˏ��tY����ij���������b.�%	Z�'K�T���{����»s+lĄ5\ �Qu8|�d��?��_*��?84LT^�<�G�\�e�������|������՗G9����j���F�
{���b�����"E�HN��P�eP�j�dxA�~��q��{}����_w\3%���5�1��:8V]k�����
�Rt�)�0��� э��?;�z�G�IJ�P�$���mcc
�J��p&8W�ң%&��C �?�&"�ē'�߼�t�Gͨ�����/^�ڭE���h��Tw+�f2$'f����I!��|���x<���ݟV<����S���IB�^S��<UH��?BGQ HzN��i��ćU���MO	�E��p|o_[[{k���z��N�(�c�3R�un�|����:)�d���v�cff��]?N��RQW9���uŤHI͔e��U�i�8�|y��^��o��yP� ��9c�a����D?�Z��j>d
�˄���	�l��4J����Ƿ�oy�Y�y�Q_p|;%?����+�G�pY�����gy��h���.��&v����QO��WF�Pl;C�r�]19Ґ��""i@�-�e���Klf����[2�zN�"�?tԓk�YD�����T�Lõ<R	���ù�m�QE6���ro7�"�-��Ϋދ����1'��z�l2Ca��e}s�X�����K���@��^V�E,z����R`��|X8��.����f橗I�ۡ����D���������P12(_<8̴3�L|�ʂ����ԛLnyѲ=�1Ʈ��{�����2�?��)��U'Џ��Q�V�s�d����h��!?g�}��C�nov�a��WT��
~��˟�oy��ڟ�_��<=�į#�������|ڎ��nd�n�E�)u�u��dUq����\j�d���hI'R�J�^�������^5��tn��t��/�槞��mL�>���D/��G]��?T���q���c���R婬Q�I!����UB��<%��>��ғ�ΣRX�u\|ڪ���j��Q�6		��9sd?��w[���L*�",췲E$���_7{����dF����2��)!�?�;t>�N5Y?M�ɰ��h�/�$99�FLw�6�>hy��ϟj����P���Å������p�����r���*H�^����C��&�zO�u�*e�w�j3۟i�g�{l������t�g �pj+��@���j��2W;��]�5�����k�7W�x�?/ p"�Vtn�(D:�&S~���åI����gd_q~Yv�-�˯�6�;�ޓ6�1	x��j�>�f�'��T�Kංa�hP�bq��d�l)m��sso�2�@.�p�Ŀ��{��JIB��'J�̣)�C�j/Z����m$24��Bړ�Ϭ��B�������*4�����NA�N���iCֺl�D�a��_��n�s?����)U��J��c���$��ۃ��Ց�2����8�}��K�[xV�o�T+�2��G��s�O�4����z�'��h��G�	1���,��G�C���g��=|��~V��B�D{���w?&[��Vj/�,��673#����N�id;1�xod|�O��l�V��s@�2�&P�_-C�e��Ž�YF�1�5@�\�
�RʚV0���Y?�ߵ߽���	���HI�'<S<Y�9Q��a����!'޷����}�~䫁^F���zJ.C(^�� �.��J,=:M�7C�U���p6�$bY.GDtx����J�u�xvNw`w�y3��E@�x_*=2�	 uh�{����8���iol��[�\y	�E��0���麞��?~�D?~�m`b(�ü�4D>��%Z�QV��B���!̮6o���)GgƓ���f���j���x���3� *�����Ԟ�Š��~��B�SR.?i��)���
I�6�Y+��z��r��V��5�T*,,�Z%͜Я�K��ߖT皛G�^ W��zzz<�G��	�3��ٟ��)�B��^�x�~�M�d�Y*)&�eS�<��S.L�a�Ust�(?��j9�1PB�Yo9�)�V�<��q�O�C%L(F������Q�0S��+�b@�s����@��=���t��W�]z��r$ܺ)���fĈ{���܇���?�΁Gr� WݎtW����їO�9�R �bI1�YU�w��VQ:澾�T�#�2���)��=t��ϒ������tE��<\͗PF��0)E���z��=n3l������k�=���a��p)Z�V
/g{B�'��R�\�澷@����B�Q$��[�px> �QYV�nQ�����}Z趰��^����%y���~�uYW\�7�����:۝�M
l���$e*�����"ImU�3td>����98�k�J�=�m ��%]�fJ
.�oƶ�������¡C���Y��9<���v��n#2�ڨv�����p�O�UcὅѺ���W+�A..׷7���y�N�7��h׻��@}ųmӚ�(~C�!;�O²Y�>L��>G��H��G��1� ��4�L�P��zH��j.�cH��ho\X��t�@��m�{�a1A"r�DW2FrIcxj���h4�C�vxoJm�k����i��C_�FU)��2�{ʝ�2�}��
���=����X#"�O�蟆v(����\0��-W`�s�~m6Y����@�:�C_� �-��O��ܲ��4M�6�׎`�׋6��ǳ��q�Cl��)���p�5�2�݄�{��5"<y����� ������Ҭ��7���Hո����<@�+m�<i֪	|;�7������ܻ��b��'#�ư�eܣ��e; A��F��9������F��_�X6���}Gi�ף���9��δ���&fF���kC"��j�1<M�Xj�4�Sn�J_��%C=���g��pk�:��;,��nVi������F@(:`�sAA-`uA�Y����8+/�ٻ�Z�6��:�C�U��%V�գp��7tr:@qm��h�]�Q!r_ka[�ٯ�!D���c�ʫ��/cf���K�����LW��e��0�י���_�xE�Om{3(`h�Q�#>�؟rL��j��-���gP�}�o�+��9��S�on��iX�R����4�['#���aZ��/�@e�����6��;;n����|F�s��fυ4�A`	[+��}�M�q���NF(k�����q���v�R~���g���?Ӭ��pe����<�3V��}�\t=	�>��C�U�"�����Ve��{f�9����#�9N7^��`���&���VwyC'��(�Ŀj��"%3�vzf��ڽ�G�z'���Z������o��p��:��fM�OCPn^���Ð6�Xk$�Z7D�r
2&C0�1��,o\ƦէΜ�?ޣl�_R��m%$(��;b��O�U1�i)�uICS��z7�� 6[s�:u�d�]�~B�L!�{�!�69e�i�ż��.���b�,((��C��13`ٚ9F<�L�"p��d���d�IY�SYv/;3;~���~.�����I	��V�#N.4݆y������/������n�(��z:���*��1QN!��bV��f��{U84�p`ә�� !99�>TЊ������yq����OW��; tm_'�n e3�܍�>o+;�'����~?�qي􀾏��VJ�i��B�'�54f�h5�c�'���m(�/�/�T�;�5,�d�7>����p�ZX�$+������p&I��iy!s�5'�z#�o�	�%g㙎7��Y��5�M���Rp��5�[���^l{ ��'��JV��z_5�ǋ��騨�����-���I��<�S��W�3�C��[-�EN�.���cE�KK��z��z��/�q�N���#����>.�o�n*4;#Z������F'a$�c������䦰Z��^?_�d��1�*$z�~\�r7eɱ���EE�\�E�ʹ'b�s�(儆5O*E�څr[��7nN&1�hG�����E�\>��8�J-Kț��UKvW����s������ee�X�18S~T]��ED	Vi�����=~Y#S�#��>f#%:#?
�����=շ�WP��������l�~�� �kG��aX����a<��4U�,a8V�����N�����7����/�Y#Y8^�~DP�]Oی���"�{�N���_[�� ���mQ�"�~���׹G\�s���L=8���Hy,_��=�;���_����־��3�TslmȦ���9��5ŉ���T���)yT�@]�����פ�	2�A8שy�d� �|8e<��J=��:���~�1l���Qɧ�Sln����ܼ:�@�qk��B:��������{�-���	�_��"��AA�vnn�n��5�r����7㚯O����bΟ�ڻ��F?L�o�iJ��x�ᆚ����d���!��q��!�,�cU
�:q$i���Ʌ�iSʙ��`��xN@T��������Zg($�j2D��ج��JE܍u7zl:����W�!G���y��{md�鹴F{	�ڕ�˦��j��-p��gw؛=�����Y����&�D"�����<�H1/<�b͙�_�XY���4�gR��h����&Y�/��Dv��k ��)��
�D�z�}��,D��yٺL��ʼt��i.0[ht��������3Y4�0l�9�����Zu� �wM��8��5z���!'0$C���)��W�J�kMٓ��L�C�S
�p��w{+��m����~ۜdin\���:L\@䩀�&{��tqX����_��3~��/]�Q�?�z�N7����Y0����J&�>�+��zȟf�x�w��2Sk+��J�"��V]n&]fB�� uު�nn
��;Mu����C�WGE�}_���H�tJwH�(�J1t��"��"��!�!1�4R���~����o֬�Ľ'�>g���7�~"B������'����4���%8�%��؈�,��+�Q	U���{)���h���
dl�{$�~<{7b�s(��lu�ď. ͖�C��g}h��Z�����T� �.$1;�_�%��J��s�*Sƣj�b�$��}9�b�^U �맓�sk��s�徺����������H�_u��&L �ٮ�R��v�|;���;���U5f����\�v-���os��c[\�ZW������P�,s��v�:���И2;aV'4�k7�xX�hy�{�fr\==/KJ��=���L98P�%��"�SQr����Lv���%�G���9[Y	�x���-6�	R��§�.���k�����x6	�鰒2�o��RN�?���'�o,�ܳ\Am�/��4�Cx����o��(��{ǡM�'OC�;��j�y�fƐ�#6�CG��vz�(B� �����������5�#vv5t��%��ur����*��}w��O�է�_��A�"?^ijϷ��s�r�t�m��c�F�����-��L2=:��WU?�K��XlM/��!��]�[|�\�ӭU�B����@��o�͹����^�	���LN�2���0��Q`	`��77q�/(p���H�G4����')sW7��rFG���}m/S?�&�z����ejgB{f��J^����I(�GI��2Z��[+�k�L�]^�����N`_!5�#p5�`�����36�a:�Nmc�]&��ܗ[\�k�����D��>�O�(�]HXOMϟ��V�~_��zZY��V���J�_���P�	���(�>'��u����aB��'�{�J��E��b�;��:�@"���L�(�P5���4����F�f��0�[k��/����5Q��&S��$��CF����5$\d?�>��$�c�畽���;����|��7�%�-�i�(�}��>(��GX����r:9>�2�\F!��(Z2�&K;�F������d0��.�oU�pe����kn-�Snݥ$�R6P���H���b����~�sQ=���A�-A$zų0��t& �S�x�0�-�����Bwa�L���ׯ1��J�����%7�$ ������qvw��[1|dp�i���LM����66���3����$�<��'-�@�۩���YNrXL���'f����f�����/U�V�L}���.o�p�5���t��5���9�8J��32���5s>��S�_�^oq����U�J�*�
��ӽ�[H��/��"B^�^���
��މ�	�=����$��t��*`��-����h;���_-��z��{��퐥���P�r�뫟+��N�'�='N4��V��m�<�#t$)�Z�M��h.�OMJ���z�Wm~Sr�"!�ҋ�Hu ԉn(���e����þ8tP�����o�ék0&oKU�8O��m�h�E&E��w�R���7G5BbaA
���Ƹ�mB�`Ţ��
/-�>�P�Gh��^l������[���ր�b\$�5�b�Q��!tם��spp@�p�-��:�{�ϧ��·}+�;t#S���3i�L�;��"F4h�����RC�gmJ�ą�wޗ/s�B.Ps�d��hD���74�L�40�0)���S��z��־x�5j��+�|�����?�Q�0?����g`�ԉe����1����&�gZb�74� h�L}#�C�n��.���ܬ]���U��U���xk
H��u��+�B^ilu�8�4"��vF�y�?��I���:H�1���s�-���B�:�̓��X��������������Ri�@�k��Γ�z0�����+�g�Q7m*��48NE��#ް��^�0q{0z�������*�ϱ��4���բPz6���;�v�aR���"�dZ+��t�|ffƗG��f�ge��䌅����q�&#���$`BZ~,5�Qf���cV1N���}s�"h��c���E?��V\&RLLFU��*4]
f�@�ۺ�.�3����^��.�ǰ��F77ń�"�/���l@��,�vW����oJJ��u���q`;9ã�����SAǷAy�BK�a�mZ�P�.���y!�#���׊L�#�C�>J�����vN��.5??�<��jlsG��9{MR���ri|��u�az�E��߻6ᚣg�,���ړ	��� ��������%ݸKR�A���/�+s��i%�����z7�ko@�YI�������Bo`�	�өK�)�$$E�9�Q�Ze�¦�� &r���d���kj���E��yweUQN�;a6l�=~�����4j,���hҍ��m�<��!:9�;��A�<��ꑈ]2���@�����d�x���g�2�G����[�,B����Q��r1�ѡ�>3@��4N�b1b!�BzauM�5/ˣ����aڄ�{Wo=�ͦ�����3	��D�dͫ�H׬Vh$ÞB��6I�����9Z��?�z�咭!�
`Uc��u�\��n�i�%�2�9`�~Y�Kf�m^2���7T�վI�嬘�3�1X����]\.��F����,Qҧ���D�1��]�a��h �B��mlpjQ�aa��=�iiȟ�8\,��z��w!T$~%b��5�98�֜���5ʨ�tKn��ʳ0���B`9���-w�.�璞�ݲh>̥/��5�(n�����iq2h�e�b��=n�{��06��E娩��A	/�����K�0It� ���^�K$�(f��k�Q��2)�,���割}�z��a�ű�`7
���y>z���~#}���=;����rT<��E��
[����Ԋ졊Ftm�rׂ�ÊL�����F �~�Bk驒�!�j��;��9X���@n�ɻS�MЩ9�u��I���5�A�)�7�:��J��o�]�^E#��"����O��⹩�5�� |�S�����B�!�J<��ޔ�35��S�7UG����/o��zw��K�+��������qqq�+K��V.��c�#���}��M����g��)���y�+w���$8::�%��9'���~���D�V�:���H"M������Ǐ�0ٷc�K����ᰲ�L���p+���+���F�>P�(L��c���\�6}���!LESӑG����+D�3N��#&��/�H9C!�d��5	`�;�]����7-[G��o�lrGn�5���O����?M��Sս����a��^��[g�˝I$��O�0��R����vT{F"�AZ�7U�1�l��:+�;b�g!LD�&#�����K%l��Q��EnUBܳ/���v��q>��E��^a稫�s���>LlL,jv���n����JT�>1*2�\�B��W�b8�7�^)�!�q�{@�N-�66�tޑ�_n���TF�`�=9rp�~`����&�x�A[���HL��3l�\P6-0s�����i��1� �/4-Hy|�x2��{��.����ʅpu־��0�^I����v���8����<�t��Cg�N�`��dD�o�0v);_���/�@!��Э_ؾƒɇ��J]�_��(����/��{��W�����R9티�~.��L���̭W�j�- ʹ�O�Z����Y���6Q����٫k��]��l/���7YO_�U��uM�OuΥM%(���\L!�-#�<�M?��k�̣�NQ�k�f\�j��@��i(�?{~?!hr�y���d��LL�ŋ��oN�I?�|��$}�<�C��>
0�Rm���{ǃ�Hvǂm�10*��S�a�T�H�Am�ߺ�o�w������#=&���MN�>|S���?"ҩ0+�Ap������p7M�Q���T�Ŕ��sȭ绊<���ɪ�:�=8��򚴴��1�ge��`>��6oy��H����j��d"=�`�v�d�'��O������~�B�Ϊ{]�jv:vC�,�|�t����E���OOד�6�9���<��4xb���5�ciHѣ0>fgB��]��w�:�=&%'JኼD��h���q�x]r:,���1�H�K�6�[{!�	<�&�.�(Hl���}�T�d�Knb���ܳ�E�3�]�;q=�s�	��-u�Y�!����BD \��G&�E"a_`�$�%�դ[�U#Zݳ�0�b��v2Fa78S��U���rNN�e{I=�/��t����xq��I����A99��<3){�_p!�8��Ag�>Qؖ�9^�&��ExKG&��Y�R~�:�5[޺z���
|p� ��f�IS�o��^ן���x��i�jƦ��"�;VOT�zLJb=A��u<��h�(�;J,�=�Ԃj�:Tcr@�&��V��Ć�(�#��0C��m�l0�^�E'��?x���bW�J�Y��#�Ez����a��d,w��eH�7�y���d��Y2��z�e���3x�|d+�o��?\�~�'-d��Z; b�.�����m�&D1s���W����X����|��a_ڽc��>�oU�DOƼL�$.311yך����l��qo�Ir(k|�QjR�@|Fpth؞�GX�8ֿ���/O���Ix�ad��ܢs�X�"�{9'�fJ���%�/F�8M��s��~�9���?�_��ro�Y�[��,E�m2����y�^��ͻ��]�]�4��<MR��yw�m����m���}�fY��(Z����I)��
ҋ�hW���C�&��  &�'��	݄��v�~�W�D5�f]�[tʼ�c6�e0ª{m-��� ��!w���E
	?//��e_���o���莦���i�hS��	��gi�5�p);��Ė��#0ʙ5�S[�~�'��5Z"�WٍE�	ʃ8x���w�JKK�c�;؛$�\ IP�/;F	T)�뵫��q���`�7Z�	EF���6F@C��~�`J��e����Uȟ�>�b���+~N*�A6�*i�H�,��E�sԵ��	H����k�[q�n���4���ô̋�E\Y��{4�8G���%�χuT���.�hN��;��&��Z�~#��ɺ��鶤��9O��W�K
1��{�3��
���c֛�j@���}Tm8*�jyTo�M+:������z	�PӬK�ݤ�K��Ę(�LG�&6q�k����H�t���P��� 1]�}�d&�[YS<��l���(�P����i�rf(���$/l7H��MԬ� �&�;�U�pVc�ǽ�-!uVw�_���E���o�Q�+k��V���yx�f��ۜį��l��4�����+%���`�KM5��x�4�&�w6a��M�.|Kӻޙ�S���u�2��������\�K��R�-����zy_��-�;��n*�pbrE��%H���"�1��af��!ᚿ��~�����܉Z����#��$���<�����t[��S��H1��p�~#=��� \��X,<�]�a]d=6%]��^�w�l}oJ��̌|e����s��)s
�n>��SqO��wT9����6@8��T����{��Ni`m��'|��W��f{N�J3ia'�a��{�o�@�*�@6JM%ì�(̠\�IG���$.�;������B�Y��O����Я�t�)P��O0������q��������dA;��S->*�"(Ɗk�z�(��������ch<//+K5��N���Z�������	Ϋȗ�HM��DK���9��V�Jx;UP�e�o�����U��,�./��a�B|^�v"+�&Q��vN�3�Vף����I���AK&��Y���"-�"Q
��~�D��K��ݛƙ��'b�,��k-*�o[�L�0s�bi�Mh��V(9zڗ�4�p5V[˦q}@�`��v�P�:�r3��B�1�,tmi�J����Ӡ��h2q��Qk�zRN[̻�K<J6�(������Fb@�+~�zaq?�N�����L���0���mN��?��yg���k�clC��U��!0GA�����2)�;ʇP��3ww�֣F�<��9ru��;�{�,P�{-�?��Ν��h�kK��������I`�/�����ht�;��Qa�x¼���r T��l�f�k����X��,�p�
����.7���z��N>�k���N��C���ED�+�$��]�L�+���C)�{�;q�Б�;I��'D�A�n�E�"�z�I�����wk#ߩ�Ycn�C��ikuy���zL�$� 0��T�:�ט��4����� -��a��8�X'LG8��L�WI^��_Օ�l���:Z$��z�cǙ����l�	v�%�x�ߺ]G�ifC�x�:0��:Y�F���'���i�
M^�g��C�{S,w�t�lN��V�в7x�%$�_������PU8Uu�0u�F>Ȋ<Ym��ﻮiq������̈́Y~׸=�CO`t(�����X�9���뚪��.�C=���ᗗO�v�8j�ΖP�)Q��k��U
���5�
Pzϒ���\*H��H���v�f�P $�2D��Z�p����5&m��B1]�z�ys���8�f�`�H��������HC�)۝���<T�2�@G�7M��4�a����^H@���VKr������K�����2�HqjAu�4�:�����%(d?�Q��}�+�jT]�~S���		���<8z
n�q����y��@�-b����4�m�u��a����R�쀨n���-lqQ��j�G�c�H`j�V�+� }��)N)�Ћ��l�#�_NOO׬���.Sj-^I��-��g�y)T$^&F��IQ���9�g�9&��P�h�W��#�E��f�Q�]�@熉���d��fe9�,""bc���LuV�SZ@�9�|�㼣��y`��q�@.�!LD ���,7'G}�*Z�/w��4h�!j%����Ш�~�O���d��� I�w|:++�M�3�Ƭ3 D��e���+���G��B|⍉����!Q�{{S�
JJ��6@��g"�Jyyy�s|cÏ�[�!t���W u�Q���(~�
`pit�
,��6Ɨ@�Z��9"Z�
·��]�#_܌�]���EW��U��'�h�C;�?�o�I�� :S�����E��?4����HN�k�f֝�����>� 8�t7SS���G�#S��P���b_�L�}]�����++�s]{���fu�1dQ+�p%_��	 ��L�7;Z)���1�F]����~�t����e�O���=Ā*�q4����i!��MB	���wp8�{�J�� ��DV	��zWfp� �c�kU�`:�
�\����O���m]ɅJ0�^����[�Hק���k80��@f&��j�,�b{$L�_�s6��Y��4��4G���'o�;~��G���*��#�u�C\.�G �̧܍
�^|r�o������A̚oI�3�3H:ċ<�bn�  F!}����ӗ}OGXGvђ9|�%g<�S�k"K���w��A!3YL�ۛ-�^+��0e4�溪tEh?�r#Ou�%���͝��R����f.�jck;T_�K�X���W��������(�ɖ�>�Ҋ�Z�l;�eY��t	=8BFq�� �"u��`�e�`[�~T]ى�<¢r�h�'X�"O=�����@�-/QhG,� �U��]:.�#XR�9����ׄ��Q\�2μ��z�~����v5�.����~��IE��������dq6I��Q����:��6r�w�.[+^���ͬ�Ø���R��N`�iS�~{�Lp��W�Z4>l1�"�~�{��(ۋ;��DˆF=���|��X�!�H:�w��<!o�[�M��t0�Q�[��94�j#��!���X�#drX-gd��r���v�Z����Mr��4Y�����!j":�H�ݐ�I-_�-��1SQ}5������rވ�PsI�]�TF�s�*dꔑ���5��
�,*��^�P,�X4N(�|S�F'IXG��[��bY��='�=@7��dY������tZ1"i�Z�>[��'Ms{N��?R�  :�E.-� :_�1��dLB[�L��{(����I���I�ߑ���N4~�eS_�H�[�H��y0&�Uy1�ږ����&ס�2Z
%�OIX�2�#c'}�8�2�_���
?�M_J���0���ҷ��O�Y(�m� �O��2�O���ؠs�[K�s˓�\]^�x\�0���X��W�=H�a�jʄNY�n
����R��%���p-��۷&�)�;GXe�_��a,|'.WY�x�tU,��I.�Q+��p�Q��p�&$x1fQ`!�ox��-�T��-TP�E��q����q��tns������hۂ�����ħ5�zf��	R�^�J��� ����1���H������{ϥ�W	��&��ѳR�wr�uF�2ﺬ�pDe�A�]����,��u�t�g�L�p=}a����H�L�٥�|��N��||䍾�fb4B���9�~h�-[*�0��n@���˦2�OL�M3wpS�a�goi�*4-��:����~��bw���ˉ�^|:���\1t4?����jov��)uߛ��XU�k//o���R4�f/4Yc��L
&[Z3(\����?;�O3�e�^��ʦ��_��%���H�K	>`�c�?	�m�q��hl��z��T�1�����w��w��8��&������4RS���w�lS�}bjA�!�%=��3�^P����h}����?�xde�1���wDl�j81���U}� &X�ap��!���6�P���g)i��I,�y�n����܃b�'��ƨ��C���W&V��j�h@��8��"C_��3V<�l/��WN)�9��͂�M#B��3V
@c�^[v��i��G�x����V�uC�;����V��f)���oTG5ͶG_�G/*Mb�Q��wp�>z���p��EKə�]�$����2�]-W���L��U��I1Q��CO 3/�y�_�P�tZ��K�͕��Z	�=)#Y+ |A�߅�V*d�B�pr+*8"ǌ#�Lq3���Ls�����e��]S�&]���'��f`|�JM� ؋S�2��Ӯ����bϘ�Dѻ��.d�(�E?�O�����dv�Vi�9Z�0J>�C�.*���C�;;���|-]��Փ��D�zq�^趭�Z���M����ޤ�2�,힞�D��|/Dh���� 
d�R�d.w)�i��coq(s2%̺R��D�
�[���Χ3x�(j�ǔ�R�5C�+D���X�r�4,qz]�̓�:�ǽ|���b�e���]�\m�٘U}���?�-U�ş��tv���Bn`���E#ۮ���.�5�G;?��,�^����x�W��,���&�Oa��R�ź�	P�lk�;$��ʎx�3��ͪ��.(��ب�5iU#d� �������
�|�@ZJ's9�9��~����e+���Q{	0\l�bm�D���?$�".�`DYr�3�#�Y��f���?t*�/7k˛ŏ�c$?%cU}$D����E�����?v�xk.�sθ۪����a�[YQ�1���8��`��7�;�_���aq��J
�)/eT�7n`��mr�Ɇ@���g�uZ%�[W��%��iJ�����#����YRx	4;��jgj��ZʣΩؔٚE��re`7��?�y!x���� ۳?7���p�����+�*ug��\���M~�̗m����$�N�=�-ѷ���V(;PT=��=mu�?`Y�����I4b�KZ�ˍ9�,��)r��e���Y]�¯h�)��Y�;��N�V����w�xkث?�D��)�w>�_�\��־êZ���J4B*�����(뿮�q�S��#B��:�l�z�خ��:Ϗ%.�ɿ���D���֊����Br���]؞�#�z�Q�f�t���%��'���d����d��T��?t�x�d�WҒ�
��ȵ����]���<��'�\����ˆ)�y��?��m��|}�M���m�^*��6�����fs����� )I����Ǐ�͘��ܓ�o�Z�4����O�~���&���c���s�&�h��� �NO����PG�܈L��i6�f���{{{����y�Z�Oc`�% ���̷�-��VZ|��j���,�[���~*���#�t�涷�y�?�}�NO�{H�����qz]���N��F�FQ`I�Y�O�L�Z�n��;�SqO�m����g�)�h��89kў[��[`���3����ʊ��s�Z�����7��"���]�@8׸�e���}P�,��EPP��i���cٰ��n"k(i��~�j�@?�
c���ҽ\��ڨf�#�f>�w�z�4�� �Tg��s�h�	\+ݠ�S�}����i�#�|��]Çw}��NZ�r��2�/kk���w�8MV�K\,�`����s��[g�cq�V���.�0�d@A�{�շyna�W�).w����Z�	�5YN��h�!d��,�t@�M�HTddJY���zh֝`�!I1�9Qߏ�������h�t
��:�%�M�W�����Ĳ����Al��[�^�
�|�I����v��$���2К�6�)!*Z'����=Y�<�Y��)��^OLT1�b8�R�V����zN��bW�\µ�L��?I�`���K���CW��w�⹟�s�U�ߋ�� K�BbW�ٯkss%�����l�BB�z��~���\G��#ۃ�J3��ň�<���G�=s�>�yI�����$Ѡ���v�O����rs�lo����&�3rF�,�Jt	�\=סU��EcQ� �⦵�B��Ԯ���<���n/�t��m��N⢟���읋e�u,lm�)ֶ^@����$������ ;0��lh�����v5�ӺΎ`2���>��$�*�9N3�k����J#]^6��T�!Eێ~�x�y�d[����&*ee��F�����g���!����k
	�����u�����yx�ی�������i��W��]g���K3#��U�v������5G��Ud�󂮖l�};^�|���=�I3�/i�����\A�:�^�,-U��9hR�m��r^y��?rm<�J&��mY&����r�y�];�i������1�0�y��N��������ښ�b�p���y2�����;�&���(���z�!8N��Yc7��z�	���/��5�Ϛ���Y��N��/x%����&&����J_�N�*<�"1���v�Dv��
	�����M����X��o�xp�"���-J�/{��T��'��� �;H��A��O������<v�����8v���<�Ĥ-�aƷǐ���"���A6p��\���.7�E)6��ʠQ[x������d��o��;�����n7�|U����_�l�\���_o�\g���
4����T�t̲�ZP̄�ɨ���r
|I,/묙�]��M6�]"wp�튀� k�>�D���^�B�_�����]�`�C"+!��������A
�.��9��&��VE�FvA����i4����ׇ�hb��B`,ק�b��)G�������b娽h�nI��Y��w�SVW0����O�&�hJ�+n&�gJ}�H��Xv]�a�b��e"6�J��[c�Wv�O-Ë���h�*�k�Qʗzv�ʜw�w�x�۾V~0"2K���
"�D��0�C��|B��S��W�c�f���:��,pi ��6bD�7���c���fΕtu�o�`�}xT<=�EjAPt	5�;X�iL�Վ�qnȸ^��S�{D4\.d��Y���x�k�����-�#�tv��ǚ�"JV��(_��#ޞ��8�ZƏ����y9(���?w%��.Mv �ue�̽�&a||<�VN-�_j�#����Vk�T�n�zGEg�Sr%sa�pi$x�#������+�"�c֋˗�T>�%�Z��|+2��f�[a /��=2��a�@.%����'�L� Ȕ?��c�B��x�����i��
i� rR%؍q�Z����	�B:�u���:iKd�A���4�̉DEDD

���1���������lagw�f��XeJ]ݺV1�.V��Q�ِo�:���ሉ����	4�			�H��#jߑlHՀ�r��h�0p�9���KvE�������u7�:��Dٷ���M�1������9Lx�"TF�u�s���:�6*����ִ���А����`h)�@�T�Ƅ�p��/wM�g��q�������m���P����^8w	�;:<B�# Jq.�n�R钢�[cg�T <������1�a��^+�M�@ep3j���з��y�*݈q�[U�Z�?����#�^����ϐ��o�q���兣��-5*���l�&���jȔS���emp��l��L,�l�u��j��lؖ!�S�<e��z�t�G��˹�999�g��_2���3����^S
[��F��2P��~bI�pD.��ؼZ\}o�����HN�UZ�Z��Oq�M���1*O"�,����55����l����d!�*-��W�p�Լ��Z:��jO�=���G+.*}/�v�MS&W&8_�Ij�z:�	�����i�ID/�	c��	2Wn%���iJ6O�DH��~�#54��e'���A��,J�t
��"���:��ǘ`�����Vw��|T>B�lX�\�Q����4��c�5�WY�x�`�̴Gz��)��(�L�6�<^EF���ja� ��	ÏS����|��i�P��s1�G��c-�D�XV�U�&�ϫ��ϡ��I��γ���ڼ_��:_��Uu#G����3���ҧQ��$*c�f�s���l���C�P�')��l��ps׎f�v�&�uqq�Ҡi�t���v����B7���`�[E���j�Hz\s���ϐ'�x��ڕC�܂!���k���
�$��îk�:�%���[�Rش��'p���6R9�/��A�sM�/3� ?�3�A������i9<�:۫���vd��B%]B~��/1
f�fV����w��fT�^t�-�{;�z�|
�}��l��5���!w16)��x�}.��H�.$8zwBi6fB�;�rw6���V�4:���C^[��� 7�9)� 4��ϯ�N�>� W��^� v�����|�n��&����.7�p�uhѠ)��o`B�&�X�u����~����2 ��O-3_�s��Kp�1�Z�(�׎�mt���xF��F+i\����K�(k&��N�c�5`֙y��N#��_p������B:9#�`)������h���-�WyG�O��M�AI٘���[�8I	�cki����,� r�v�%��/��f��v��şHY�˩cQ�(��`^&4_��y���ca� ��H��*ĸ��)tVI�T�;�ڋ��1U+s-/x��_o�����/���7���X;��l��y��AGGG�9z�e>1?�B�JH���p�\=�G�lgMc+��@~��l�[�� ��́��]_�	?Z�h�be�0'��_��:�`_���EV �6�m�bl!"�5;]��Kr2�U�"k�g/C9~p�"�,�Zω�=�Z/��MXpl�J�P)0�������+��=O�\�a�c�tLS�k�*~JD��\d^H�gQf�z���Ak����4l������@-IΩ�����J2qЮg�	�ɶ�L��\��b0�~-x�}-�j§��N\p����f�Y5H�`����2���4�j�oB?��o�r�(P`��d�����@	�N� �UP�ɀÃ��
���U�H#V#$�Wi��ZJ��*��`��_�?�~�4�A$�]R������[XX�̗B1ZS�s���L�>��a��=F���4�,軡�zm������U���z��S�Y�Mw����W��{-�����]���O��P��u��[,�j�#�.4(�NE]_���>�EZ����ÿQ�g�v��[#�'|̔��Q�:糑A\��~K�p�'�r�>�\k����G�-:������o� ��k�.��W�xφ���x9צW|I�l_�Co�i6V���P,��G<�o��v���fP����z��Oϭ�pa�%�`氿x盺�&M��V
���<�z���F�Jd�X�	`��ç���uu�E�tBa��d�^�����jD鈫�GX�@KC���vn�g+���"PO6����=e϶3R��.
b��
S�y r�=s�?ep؍T��ܩU(˟Ȯ��n�C:ʗ₎\��ȹ�o|~O'<$	uD�\I���G��M/�����B�����fvdo?��P��}����\R��NZS����v�V��&;��%�!���iCdsHS&�#���G忝Q�B��z�\p��v�����T�����5���}AO�����
S=�#�E�����
Ӿ3#�����oq�YV�s��_��;I.�#>.�I|\ܦ�����ta�%�	�$#hȗ��As�:�0<|*���%a���|�,��$�1����Nf�y�Q�![�s���l+��M9ދ���u<@��$!�-	4ԭ�u��~�;U���F��iL�x���t���{�ck�=
ó������V~�e�pF�,2�	3��"�fY �C���4,����?5�l���49�֭KM{�p���Uۇs|�gzr��-t���+�ZB���MH�H�h&�e��p�n�	;�j�5�g;�7][R� T��[,{������?�	Z��{�<��F�Z��֠�J��Q�<�̒}��V��ԏ��<s��_��l����yyv�4�.���m�����ֆhW��rLK��"j�����bE����{7
����7��|)H�5��'���ΦWvLn@�.~*�E�m��I� �E��)� ����9uX.�u}ш]'߉�C	�p,()�{�5"�]�픽�,�uֈO?�WI{��%�Q�uu���k⭓��Ǖ�>���}{���ߧ��qt�f{��p�{��,��K��������#���Q�����6c�Mj�xoK�:��J��]���@J�6}iEs��5%��3���q�/9�HD��
���|s�����d���{��ī���g��a7�]��C�][���}����W?� �JP���=(
Lr^ �j��n�*��������Q�޿ŧ'�z2�
���nv���Զg7��ͯT�ݢ;��հ$�{S�J��Ű��_�X]�ךt�y�e�;����C������?sC���yQ�V4����#Q\}Ѧ��\[j0fb����z����F��7���g\�/y��<��@@ʚ+[VD
	�~��rkP�3+�=����9��ӕ{e#r��=��(�`T�w�WO�B���(��nsJQC���O��CL��O��oO�{�Az�W�q��'�΁�U��)c��h~��v�bJ@�y�<�!W�����ׁ�Cg���Y���]�+�G�+�q�3VY7�uI��j��'�":��Pz�A��(튿���mA���e�y��:������J�ǂ�~����G��_�~S��Ϗ��xx�q�@��LJ,OG�Jݺi���B�n�kF��z����XN�àrc�P������Z��l;�p��%��2"���u�p��9���t��Գu���a��D6��s^ˈ���nh�nM�r�f���u.���x���� tn#�Č�D�h�m��ߊ�`�hI,�ٛ}羆!��f'?�#��6��C��h�)k�O�O��K���'�+CH���B���0��q�Of�!�\ܕR�/
.}\]'�Q�뉫�
�uq�y�82���َ
��Rv(+o�bm;c�������a��Y[�D��*��p�jH���,Y�T���=�61qh�-~������h�.�.��@��`}�A��p �%j��L��%u�r?�=�����	ښ����w�����͵޴�/��c�0�	��@o�on��/�/.�u9�^%o ���l���⇷?Y�/�}au�BW_.�*`��V_z��=�Odw�Q�O�N��j���[ܷ�_�H���n�-񐏇�^����< bt6Z����SJ���6Dl�ۻ�w�H�AQ=`6�h�u?{�l��灙I��~ڜ�El�62)3"	EQ\�A�H������LLw�N٥���Y�����؎b�ʃ:n		!wC9�CD.���/��xZX�yݠ�o�tۯ�>χő��l#} ��Ip��.�DD�..����q�S�נz�� �:>7���$�����&[��b�QۙOf``]�F{���*��?_:mǪ.ۡfw�oĳ0�MK��;���穞a��o4�c���Å���jRa'
��K�� �����j Su&NT6N�:"���Y�3=�D)�}�Hv�:�	)���y�p�#FZ��q�m�4�HrZL^�s��m�,	h����a�ٚ\�ć�0�S�g)|��	�cS�uS�������墒B�kwL��d���[�/-�M�wM����8�_�en.E�/�����/���7Z2��R�/C��!��1艵���5~X�P<�~:��<�*�	GD����ap�=�ǊFP�M@�ܲ��A���e��}F�:�ܺ���ӻUΪ��K����i2Q4�|Dv%t��*@տ��`+Q�詂�|+[ѐD@Jf���*Kk�tD�Ѡc�˺TM�m�A�@�M�YZ��IK��kڮiU�p���I������;P����0o�kiT�V`S���پc���7��%�X:���L���m��� �c򲓁Z):o]��D�:�ʱ��襗1��]���9�;��L:��P���A�LX��UD��pG��f���]���Y�we����{�����>$�	�K��Fw�Xd&k��vb*�
��ųbS);i�N$�[�RY1^#�t�
�a'�r�6U�!�_p��:T_i���?��ތK���ߠ�/.���m�^��	ٸ���{��	׮�yV�g�M�ɵ�am���������߮6 }1�O�;�8K˫f2����C��@��@�h�涞����h�����`�����z!����p��z�3�<�*���,�Lo��	�� m����uKͬ|f�֠�̔��\XĒ�������wt�֧�r�},��Ѧ0_|B��� R/��P��Z}��4RGy'����ȣ_�;1@�7DuZP��m��F��'����$ƽz���>,��gE���遲;Q�Ocg���tY4��4j&��;��6ðt���@��u����l	���A�7�w@���CY\�z� !L?��7��� �˘X��b]~���X����?��p��FZx���otcdx��=�;��ܝ�������Н;w��,q�����/�����`�Q0�u{���l�cq�I�4������$��vqq��E���x�uA�UW�m�ؚV�9]@[�ÞD0f�"dʹ���l�*�ps�a����'����,P=��í�����=����b 8Rdi�71�M4uC ��oDӮ_����� v�Q$]�dⰓ�hP�T�G�8ց���X@���h���U˛ �~��_���Z9�o�,����y�!VF�~,ם<
-\ˤ�-G�ůB�bHS����˭`ܿO'<z��Io�>�5��X	f�gϞ=;G����o�;{v��ɉ�S�Nu�'zG���O?34337��3ώ�������o��k��б���⏧i�^]����)�eh�-�mZ�[f�L�7Z6ӉG�na6Ѵ+"�b����%=ִK��k&i3<��Jk�a��w~�y�!�򩃎ʳ��I
]�Xn�. ו�l��t����[?_�Y��@���zĔ���4ڮ�MBu�����1�b'+:����Ť�_��!P��!�5#���f��8�'��-T����[F��OH\cw=x3=���-���a|��
�~O���-�� l"�t��|%����e�[�q����V��{�G��o#�?B���=�䓷�r���'�|���nW[��o��o���_��ݼy���6߈�~�g�"��$f_c ezG?�r��53�n:V �����dR2�K@��y�Z�ܫ�Z�S]I�	f���AQ����'�XW8[3��^[׫<u����T��iˁ�e���#|��r��t��7T��l'ehK����y�Ӳ}��Y@�E�=����Z������Xh��\4*��!�
�y�����3S����}�:��Y� >hn6oڵ�y}����򎵀�'��<]'��I���r��P4o�k�=���I��>�bDVΊ��X&ebe�I��4?�w��F^C�J���U�������"����?����^��W�7ʳ�⽶�|���?��?���>���,��1��k,'�s�vN����$�0�h��) ��?�|ǋ��+&r}�DN'�����L���	Z�&�|�亶x���U����ѳ�xHH���@u'!�8�򄯯NZ��j�Z؆ޑIN���`�y���7�_t��>ͫ��c-�5x���'|��4���:�����M�w�;> ���8��De�C��UO_^�|�����
`���u�u�R�$�KؾI�L�)�(�\H0�E�N!\�[�C&�[~��-
?e��)|)�I������|o��G�xo�ӧ� �������n~�i���~p���׿kq|���A�)t�`�;@G5xk�p�wv����F$�p�'�K��m\�Ә-��mW��&�-IXw1�h�.p��WgiU�i�]����Y���<W��G^�1�d��+ԆP�6�>���X�d���Y#ukD��&C>����8]@-�ap�Z�[fh�H��{Y��G�L��}�xO��r���M�-]�:i:�O,�-³Ԑ�/֤ͫ����o⌧'����^���WC��+c������׾��������y꩗5%�L#<�N[m�z�?���?�3?�8����^q��h<��f���^���Yc���w���B6¾�wmM�֤�
G�v�3���3_��Y�XN�@���^��gR�P���� �m�!�5����ʍ�}��Д�Dxł�����#k�ӆ&2�.1����m�N��Z������!����)/}�>ڻu��I^=������=M[=A��5�� )��q�aM6��o.H�v������B}�Ֆ��K��׺ޡ	���'�4�pI��C��xY�F��2E>���Ƥ���j�F�SSS�?�����^<�t>yi�
��g~����_���'y���Fm�ԓ0KȺ�m�$!D(��`_۟,�k��մu�A��ĹB��X��&!����-�N��V#45��!S�Kc=�C����u�ׯ!0��< w��&*���"�%����E(�Ѵ'��}�hK��zJb��`.��& n��t��tB3��eWHN�&ҷ�� �}R����T�� yk��=�c�����O�����ݒ���>0�lM}�#�I@m2W�@�	�,�@7;���>�c��������^�_��+B�e��������ԧ>����*4R�Tg�ߪP���`�w2�h�dj�����{�Dʐ�<��WL<��:��S�;!sq�(�~O�-��e�JƵ-eY�"�|i�gYi5�}�� 6��H����C�������gI�,^=l9Yuթ���~������$!�����Yei�n�.f.����磍��Ǿ�j�!����҉2J�Td���[w�j7��&�Mޫ-Aւ1���I���;qq�a�*F�e�)��x�>�{��n�,b�bm�8T�1���Bx�jG2#�y\�����?���l�A�in�}�<�XL̈́R���1_; d��ߧ�+��"�>a�Ӥe��zy �%�EA3/�+c�z���ƬɀOx�\^
y�f�3��ؼc'y@⹼z6��I��o^��.�a�q�楗�t�4��,^��g��TtR�Q,�F�'��24X��ܔ���u:�;f�L��^��Y"|2(��E���=pJ{��矿��h�1y���������It�iI�q�0K��w��QM�
�`:Ill2��X��c_����ig� �တ}������A��qj!CW���`�ʏi�b������%�%�C����`,���Z8��5���x'OF4�<o��H��w�dS�O܇���Wkc�~����lsmXׇ��G���Xa�Lӱ*�x*�(2a�ty�&G���ɫ<Y$4�D<Ṇ�h����~�ÿ��7��e�p���}���D1{�ԩ)�T�]u�Ԧ�"멶��J�`����k��2���ɐ1������W-Oz�CZ��>\�6T�)��C�8�	�I>R����޵u�5��C �ib .H�|w��7[	>��O���Q��6���%	�_�:n � zL-�u�Y���;y���O�x?k��W~�] �{�w��w���3��YmM ���Gɦ�ꖮZ�Ċ���f�yp�Mc��oΥޱo���)��i��Z��+Wi~�q-ʑ�5#1��P":���Vd��o,k!��K�$���?�ׯx����+�v���zB�Y���l=��g�v�0�a���H7��
[��vY ��0�v�#�k07@�83p��r�g�D�'3��%d��vuPV�Y&=��l���K�,�ړ�jAT�6�ڡG�,P�*TC��[�u���xH�T���+\B�-K+�|�|��Gǘrrǆ�ٓ04c��ڙ[/r�'PO�{>:}�Wgͯz2��>i���]`p�������ɭK��]W���\;�9s[�#�xO��ϰ����R��ט<��XP�W�y���M�:K�]󸯝|_��&Y2�����bݔ<l?>��7ig\�U�W�$OD����Fx��iM{aa���i7��h�����4�����Z0��!��y
X״-���gA�6���e��7������.3V1?i�z}�� -�W��|�^���|��<��B&T���W��_���BZ����'��F'�� ���hdS��kHm��y�5����z���Wz�IZ�n��-��J�����B��E�ן�.�I��}є+��rм"Zx��ie����j"V.����#���X�|��u���I-���Q�rj'��J��<`=��'��~c��,It?{����Q����C?`.�a]!!�1!Th&���>��|�|��93�l&��T�853˻2�C���%"�q׵]����6՞fOhB��+&m^_߹�Kj�K��O��R��"�=9��E�-�1�6M�z����g�-4r��O_?��;n}ϵ���q�~>���@�SV�CyK۵�@'"#��Ӵr��/�,����e��6��yxB��.�_Z92K�{{��ܹ;S֣J��}���I���虫f��0w�j0�=��q���^��2*�Q3�fp��Y����2ڌ�暟\M��,����[����yf�����I������v��M|UZ#`�z�i�݈�ݴ��4+Z����Y�q^�|��,�wy^OB�dZ�&�,��}�-g/�cU� _9��)2�2������N��Қ�]�h�63�T�]7�)�������G��-@���@�ӌm�yn	m=��ɄY�\b.�ٚ0�.ם�f	ɻb���	�ED�	� �u�A�W/�>���j[��#��m�Y\m�W��v�0�:x���ah����;A��T)B��T)F�����@U���E���[�aV�"�Ўy�M㫛�Y���iK���ԚV.��CӅ��A�bx��N�=��h�|�]/�K�<�yBZ[[=�ۿ��}o���Ox:7�ݖ���_(������䱚uaC]��	e0��#)�t-��x�r�����M/��z�䀟�E�hc��8��ٽ�(2�8,h�L(܁|T��)mԖ�Z������p��j��f��ʍiK�nY}�'�Y�C�ܴ���qL9��	�/�V�É��*r)�NY4���R��%״j�o\�m"O�]�8���]��r�G>��%��u�e�����K�aM��Jow��mlv�7�UtJY�H$�V,��2�;8��50zؘ(�':�wC�� �	EY�L$L��&urtp���@uZ�d�h\F��5���K�<A�U_�c�-F+����������(M,�}MҠZ�ٍ�jWh��`_����w͏>:�W\�.�<E.i�<�aDEk�M<�]��KGL�Y��� D�Ў)���mԸ��׆Q���<��P�ċ/�H���m��j�@U3�y8�Y��K]u͸��݆�%�5C�tز����XPaj������B jo`���}�]��lY�x���'d����M��~��B��h����q��I#e����c���}7K;צa0�~�i7�y��Nh�����'!Z���㌀JyDp,�-��k�|y_@]�Hj)�
����O�CdTl�i�zG[9�fwwgptt��?�Q�?����y�k���ӣ��s`�!��#!Z�t�� ��-״�b� �9G�؝�B��u�gQ�+�u�:�B+�v�>��,�KG���l>��Ut ��������ZE��K+TC<܌:G�]=~��~7��<CZ�/��>0�4�3��O�t�IX4����N���fc�v-��g"�\�H��Τ6Uq��3$���X'��D@�;ޗ������l	��3Q8733C��c-��A�޽{' ڗ�S�5=0� W�a-l$���s�R��L�3遦����'�r}^-�rg��|��7��[(/wP�h\G�/���Ҵ�p*��E��Hڼz��q��(/�<89(��1��<�^#U�7���4l��S�_:]w��~����7�M|�*��>z�������1�<��"��9�2�%O-�ܱ.�/���&��D���������~�'�c_�u_�����6靖ml��:��{�	`3^>S3P�|t�1i�lO{��zi�v���˖�}|���2&���>S�X]��
�>0���Y�����)g���ج1RTC/:޲��ڇiG�zW���Ռ����<�iۍ�%��i�Ey�&ym͒y>:�v�vK���E�iٔ5��DVq��r]xBd[�OK��|����+����g?�Y�����~�Ҡ����~�G�"fb$b��)�p4P����;��)�3Xr_N�{��#�K@� �m&p�u!o""�cg�y��D ·����	���F��a��;�E��h���e	߇�9&Ir�:k4��;�����/R�;�|yf�w^�h�Ӽ"Z�aڜW��|� ��2�B���}2Gk�Y�"�[�e{�l��w	 kC`�r���v���l	�c�鰮���ۗA�!�-�,��0W���0�!��Æ*u������i��	��ԯJt4�T�r|kI�9�,S��|.��h�̐������,Z�S g���bNM�`�:!P��7t^'����"<Z��!�[�Q��le���ִݾv�2�N!@��X�����Zv��BP���ס�ו=�_>���!�O�[�%J	�R;����h:��)I���å��wAܜ�X��.�D"��O9J��}wg���y1�r[n�WKk��?����@ߥ�ݭan~�gh��u5�1��"/�`"a��cZ�f����$hF�e��rͿ>���۽�iˉ_���#$8�:g$_�u;kxX�yt��&�#��n�L����A%7��fn����ut�i���H�1��,���d���x��|}Ϸ���}þǕ�>h�]�Q�4�$��F�=w��֛�	��%.�rȥ]Hf�}��+J�q��6��Uץ�ަo*��x�F�6
�@e�cw���������>�Ǚ��A�֭[��b����ڭ=uK�"�kR\��#W�e�����m1��@�䡖*T�8�	��S4����2u���i{����^�� H�����"x�1H��By��?�>>��N�>o��y�4��Y���F���,��p��|���4�-�D�_H��:����wt��F��G[��.�[qw���H&��N��liОE����+�4�L:B�d|��TY�j�Ռ�um��B@���� �;Ȋ�iV�pyǝ(����`� x^��1o�5S�ΪK����Q=o�z��n�վ�Oc���d�����4�ٹ�����E�I��.W{�Si-����7�BI�i��_Q�6��]K�CV��r�B4���py�Q��P��F[��0ɜ�ix�&�-��Eՠ����zG�i �|5�ф�����B���)$��jm[��[����6��w��<��EA��j��U��4<���.-BC!��>m�a��*�� ��Y�����&�.���_�R%�o�ƌ;>Bu�7}�Wf��|}��Z�铽�<��G�;�b�Zc�˭���14	�}�&��׵����g˝�ݲ��w|�w������`����)E�;4\f������//�x�Y?Y�����(�=��iK]���]+��궭H�1i}���g���$�V�E"ӏ3)2A(��`5i��jWl9����.�#�/7]�嫁`{|Z`VVB�,mR?�I���~�i*���n"o���1$��s�0m�ϳV�t�ɹ��rf�<�����{��h[1�9�4-� V�z۞F��2;�2�f���Y֌V�_X/�6���/�Em��44�b&+Y���[�o=:�6���B�yϽ����5��('YU�|E��M��X>����1��Zml[|�"�5�!�x�}`3��C�7�W�$%A�B�/t�A�\�9e����no���}R�<�է��0�wa��t1���#]˂6�520P~Dp�'mi&���:�o����Ab���� c�1/	i*E�ן��|�u�W#�3��9�?4���#�M�Q <�:������A��s�Il�y���1���7�C /����\�$M2=�p���	-�n�����(�E^�w�B���e�{e���xgk���VJ-�;;��CãWA�^��Z`��灳f$$���̐�P�i�%�I]}��!@��i���|M4y� qA����BC4
�z�}�p	1z,�U�k	^'db�=�*����9	cۨ�5@�v��w�������Y �7��V-۩�1ok����O��o�ƪ�����>ỡe5��4�R������.]%ң�b�r���)�1t����n[u�|�Ժ4sǞ������Օ�+(�S��=�t-���[� �IY��1��]���|.�V3��9 �A�+C���-��0w��\��	#� m�-3�]���Mx��1K���Àn^�yϛ5�[N��Y�	�Y��غJ�Q/�����,@�t�W,c@YƮo\�ƃ�.]C�=�|�ܾ���-+cǍKW�/rP�Ew� ���&�~n�4�}�j�+O��L"�9���{�;��w����7n�3�H�Hײ���ȯ�]�nh�F����5��i�n�}e� ���;��-���z"�Z�>��umYЂC��}<j����ȖW�������.
E�׬�y��=o�m��Ӭ6�b>Y 킦̍���Y��:�F&1�h�';uh�&b.ݵ�uU�|�<��tzWѲ�7)�ڶ+�20���Uמ~�� O���9_��_����^Gz��]��,��y3D�^� -��0�+ t�w߀v�-HO"B��ݘ���Pd]a�7�����r��i��N��(ϋ��'>�x̽ i�v�;���'>`���,P@�ֽ�q-�dM��:*��;���M�B��'�?}��N�F�kQƒ絗^z���[&�iKjڈ�=����r�ĪsB��!��L3��v��N:\�<�����<`�sY&PUm�ۖ�I@hbh�f�Bޗ��	@H�8�d fbsm�jO�>y�a��)�&>��Y�B��㗣�v]���Ѡ��d�q�"�%��㶍i��Kyr�|��1��O&�r�-���VVV�q{�U�JK���������S��a�1.Z���k�	9R���48�ھt�����v`�C(�o������<�C� ��!���;����=�b�ߌ2�����f�3��kv�4;?7y"w\�4z͏���4���a�w_=c�_��eE#}��l���ƭ�#�3-��Ǝ(NL�����1��:o�]��XQ�N����F����s\�[��N�<q��˷^킪t�f<Ⱥکp|������D.��.���C��3=i��y-�1�W���A,��NHC
��ye���0��]W@VۉE2�ދCpx���x-k�]z(ckDYu�"�������Λ�e	��Ҵ�����W!މ����Yy�<Q�e�:�"vUd��?x�$��+�Y� �Di@��n}b��G��Lֲ֧ �|��ѝ��K�������W��h���l����_����4~��3���u�@اQ
�� +tO��R/�1�
��@ߓ6������/�� �(<d��A~�"z]Ӽ��%L�xZ��9纎z[b�e 8c��a8LӃ�L�I �����:q��7U�_��=o�e�㎱��te��/c�\f�j;���9�P� (��]�&rLdl苎=�׳ݶ�ȭX�����W�,=�>�{H7�	�g�5�h-q�����O}�a�rm8d��1��.`�,v �D�.n�>��0����c����#|By�j�m�uj����_�}��a�4�W.�C����-�-{o�:��������]�H6w6K###�Ҳ��^�W|'���fz��ha��ժ��[O�^�3ϐU#T��Q�<�O��P�*?�^�dG~�4�Ad롃O�������k�K#7���xú��g>�	g�r���/��� {�GH����/��>`+�ƭ�0�l��v����B���:�̜�0?����<�#���'�Wy��=/R�f~V�>���ه8��|��i���6�z�ͫ��q�ˡq�R���q߄6�N!���Ŗ���bhQ���/b��u�E��eF��NP"�9�w�]���,�9h�y�,�[����'�\^q��}Y&w)'ԇBGI�2�O!���-���h�8��ry�gh��I�*�:>--�>�t;�� 1��\���u� wm�}�Ww����8nd1]L�b�S3@6����1��U�����Ӂ�A��wJ�[�f��~�ft��ѱR��@��ٜ��`_[_�@�/������=&�&"Tc���䎷�>�KS����b���[Q~#� 4�|�"�{�ZvL�y4�M�d�<,����+�XWcI��{"+ݼC}�.C�
M��_*��\������$�ߎ��Q�k9���ڜ>G-DV�} ]�CL���	��dB�!�i��K﫟|]M��Ybڗ'�b��i�&!�6K5+��:�l�u[_[+��<Uz�;�Xzի_]7��'N�F��J-�����Q���CU�K��_��?����>���.L�'O��3�7R_w\�
�F�j�wB �W_�^ϹcB�i���}��ʅИ��մ}���;K{gm��Vɛ�yrI���%�u=|t�yU&-����w~��}�o���}��h-�����{�����>B�Uc ��\��7��bA2��&2[Θ��- Dc�H]���|�~~��e�3=��o$��+Dp��/���{���'�x����l��S��^P8�m�3�;11Q�r�1㴶��Uz���]��o������ϗ�տ�W���%�^�՟n[�]������N�^��dSL�C��-�i`�1�G�M�ӽ�|����ߌ���������a'A�L(B���ʙFǕ�'�Y��ןE��K�����ִa��5���ܞ���m18�8f5C�Fa�c��Z��C���k���5Ҿ�����d�ڴ-BS��o���Ah]?��o��;I��&o�$�.��Y�z�[^V^���B�`E��%���@��N�����0#�Ѱo߾]��_���3�<S�Ґ1����N�*=��㥯��?o>	ң�������,ݸq��]�Y0��+m�9�߱��ZX�8,�N��{0����f�!�ϙZJ��<�'''M�������|�,��=�Ib�����v�<��̙3�]�x0O҅υ�t_5���lL�f�.K�}�'�we�;����sh�[_CgUp�uY��=�o�~Y��e��
?��|rQ�7)3$�\�&x�{x���B��/_���>ǁ��A���|ݻwh�O�0C� �Y[�Sw��Ṁ�ߗwd����*S����rf�vR�	r�����u��b�4Z���뇘�}�3�֡w��y���Y��{O�����	x1��4����o7��g4�_�t�����+����ҧ>��� ��̃���t陧?]��_�����~�t��9����2���T�woo���w���u_�u��gϖ����d����iN��v�)�����f�]9�N&����菖��[��h���|���%+�j�?�ԇy����v�@��������ݿ3փM��vKy"�ܐ��~x��c�Е+yc$�ܽ�5�}c�'��{�<���]^�h�w����l����Y��$���v�����O,��J�U��A��ă�s���ZJӆ�1�U X�s\w�8!ƔNsgf�||����2U�>���l���_��wb�V� �^��Ϊo8���LY���y�c���h�ܢe��b
�Q���cX��� �Q�Ԅ�tf|6  �ű4<2�7�7״� ίzիJ�z׻J_��_bx��?5u
�Q������@֘�������)=��S�����(ak�1�������ܟ3<��/�����3����	����2@������<���/�������_(ݼy�m�t��eд��O��_��_h������ҷ}۷�>�����e4o��J�,��a�#��c��Ҵ�,pӹc:�.Y�;}�d�//}^=�B!u	��7�ƂS���h����@�6��|���	�!�3؞�2�C�b	k4��ᣣL�R���I��"c:H5ȅf�����E[\��o�yC��!�d�<�j�a�7��, np���D�=����;5ޯ���1���C
��%�������K�}�{K��_�x����{��=�3�K����`i��XS.�>��O���{������[�����6�YG�4��#)�����{��%�c��������}u�+���*�����!�{���K?�C�Z��������S��6������]�{���[{����������s�=���D����z�������:���w}����G~��S?��K���"��e�i)h������3$�x�Ԭ��^����{7$�b�h�!�M\\JO|��VbB��P����7Y��E��9~1�E|��J�4�;�z��@B�qt�q�q�o�4�<��jY�c�0�����
�{�c�z�
3�	b�����.�y7v�'���W��)��Ee�t��in������g��K�A 9�����f6v�£�$�m������%��-�$��������˿�˥�ӥh�\K��w�wM��O�)Sj��p	�تR���+����ŋ�~�S�7�7QƮ�̹�M�t������7 ��s/T��fff������&3f��y��zCV�e~~ޘ�?����.\�P���ͥ����*}��7i8y�/k���s�n#��Uv�x�����i�n�!���<@���AVOB4Mۭ�i̾���z/��!�����>o2ᓗ���2dL�,	��2���s������7���XO�Gt�h�A��?���|�0lf{pM,!@���2�hBn���w)W"YI>�m�f��-�~$��>�B*�+ B����(��(`7�.�O�AN��� \l�O�0�S//}���e���F����>��7L`���Y��_��ؿ���h{p�7 ���G3�>�1e�B�'/�Ϡ1���o0f�=LV ��6X���~��-��}�CЮȘ�'&N�!�|��M������3!)����� 2�$�=M��k�n&"�)�����Y���V����@{��s��{�vUˌ���s-���;�%��\�i��ayzM:f���������O֤"�]�,�'yZ��T�5E�"�q�q8�҃����m� ����׼njiq�}���*s/�L�fxx�t:��}����;�n\�=
q
A�>��@y�BP�scf�y �G�4#���z�B�g(}Vݳ�1?�c`��4Ž��K���� t0S3���~�qS#����ߔz�?����[����1`)�F���	��v����c#���u�+��S5bjʼhJ�q��
T��%�-�s��&@��Wi5`�d�϶c��4���k�v8Q�&ߋuz>�%�훤�6�ώ�y#������<��wߧ��j�2���P�hd�:TW�Q�-��<_^Y�u�m�g�G�,Q�j}����O�����?~�7~s�(y0/�Ѵ1�ǚ�0��?�\!�邟�7�r����A���P�n�5Xkr�?���]���el�����y�*�F�8����=[�{�	r�>��ۻ.]� M�z��p�e�#�4���p��V"du;��r���"� ��M}tD�JC99��pf�%.ɏ�n�3R[%"�y���*i�[ [����Wh%`.��Ǚ^�W��i�\�ֵ��d�O6j�v�]�D��+>��q���t�=��H������4�6	
G�SpB;%3=��%t?ݎ��<||X�#c��?-x">&��$�^��]�;L;[v��/k�4C�s����������opz�S!��ǹfݏO�{hV[�zB!�4S+~�g$�����.��4�m�O�Xuǒ�|`�����Z^��f��,�:$�b@�m�;�I��'����L�0��;?;;Gg4��􈮖ا��}�_�A^��p�q����礣{�e�P���\��ݙXh ���<�������=�~��B��������iOTF��|,al�TI�{��t�Bd���;wJ�?��Y_&H4�Ö-�S���A���	�L�Į�iV�u>�䏐<ɒQ�m��yV�$ol�0f�c�ueKH���;�ƭ�Of��=�t_��8���?����B�H"�Q��o��1�{�lj"ZKp;W����$�cDs�>�|�	��ǥ��0"y�f��6��<�E�F�!��f=?��ɤS�?7��h6�	_�qj٢�
�������;�C�L"B���F�'|z��:7��[)dZfe��� �=WV�4ż��u�����y|��"���P>1u�I��S��0~F0f_��O����aǕcb�� ml3� A^��H w��O4|��wϝ��C}'̬H�ڊ~�\��d̽��[�5
ʄJօ�D��,���t�j�|}��:޾	^�MsX^���cAF˹�6�7K.�����[ 4����䓧\e��M���1����g?K瓵Gŧ-aGP�\�jS!�x5�������:5Ox� �ov���Vw��{�z�e��b�����,�O^z	_+ڶ�4�d;�uZ���l���7���a�b"�6��!�4�<�ۢ�wJzW����q�Uק�tݛ�!���!�+�|��`�����Cad�Gv����Ќ�����S1���<ϛEj�^#��3k�L��|�<��1>�s��y���i�fƬ}h����g�˺�G�FC��*�m�#U�S�;�uȞn���*��&cY�Q�nY������5�P�>y49L^�}�K磅�Y��@(�^���}��	�I�e_Y�~�m�4�{�����OyJ��	2���C�������^��,	��^<���G�i�����AL�/ �F��zƧg>��R��y�&K�Ā���W^V��r���{�|���M�GH�M[�"㩈,i���Ա�+&���.�d+VΚ���a���.�Ķ��Q,e]�/��>�'�\��\Ǧ��pV==�uTh��;'���/���q��7���2eJ��p��(y��)Q���
�ˬ�֢c�h�ecȪ���i�aw*d�����j����}���Y�Bl�W!`ѯ��z�4+�#m�@41<<t*k����cfF!����{/db	�?��L�MC�λY��N�4�omw0�S��u�{�Џ�DWW6��Ez��6ǶC�gu�c��,��ͿH:���]��G�<�(@�!,%�
�H��;A�U/��S$����%4d�̘��s_'��1c�=�$\�Ŕ�7I<N*ZV�5�P����:6�n�ΝYZt�|�i� ��V�����-����2��!o���^&7��������ܞ�H"�=�5m�/\����y��mb(;gO��*��}�ڭK�< �Ѻ�.�%�X�Wfz�(�'��0�Y�Q�Ș
ѥH�H�,�:l{�� ��y�<��և���n��������!^E7��{��c�g��<,�}����?��3������y ��e�B)���5
���<�L2o�����4S0��G�Fם,��e6�L34Y�ic���/R����ړ̎}3t)C󊛾�A���y�f[~�|����,�x����ڟ��,���H��F�q�kh����b�X#u�i�Z���U�I�-s��J����7��L+	��(|�eK:S�P8_j�����?z�C֟���L�H5�~����O�J#u35�Duf�,f͒���,���:���6���N.��1y5S+k$�F�)"\�I3�����}�O�~��}��ڛ'x��'��y��~��A�]w7R��G� ͝|��To�wC���y274�����'��l�W���+\���Y^^��[��~��V��2�#մq��I��.�X}ZK�v.Y�iB�� �@{��K�<��{~�~h��Z�lz�N��Z I[u�廞6�Y<q\4�+���w�����,��O����kw:���tkV��󆸬��O�����ڏ��?������x�aCf�<��D(h��	��	A�p9,��9k�.[W���&�kV[}G��Io;�Mఞ���[��Y��A#[�t���XLÇ�d]F3�l3�C�G��&�!kF,M���yeŖ��3(��t^���?>��Ky�6��#������o��W���W\������o�O�v��:0Oc�����q�>�F�c���\�*Fxվ���wLyn�C��Esy'T� �a�6D�F�-krʯzf�O3��L��H;;&�Y�f���Q�a�qVdҥ���E4�҈2Jf�������L��v����@�S���B:�D��C����l.l彬<�:=�y��$��,܇�+��G-hd��5Yq�0ym:��Fhr�4a��N�K���v����z����E4��8Lmc�S�9���o⥗^�����y��ihc�2��� hIm\C �5k�c�Úّ�vJ�p:���˻�:���z���Q���8h�W�Xz�Į4hf?�N�[�GQ�"�Ь��lg��Ԋ�4Cޫ�?�і�<�v>2����>v��Te��j�;�d���!!��؎tM?1e�ibV�[g���N\�n{�z�2YH��X�f1�I>BO���$��æ+RＲ��W4��Ļ~�}�z#un�>1���>��y'KI��Y�q��~/��Y�J��[�ӓ�<>o���/���$�ۉS������~��v�k��7�]���h�� �	�kܭl#��;!��8;"��,�����J�4z����yzu]b�QԡS�<�p4ҶF��t�� f#�}'6]QZ�d����ȸ.�7Eڡ��2�B{�s&;z��M��D}������5,��>����y?L���£{{�f��� �=�{y3آ�S4}Fk4��E�T��<+?�L���h}�ŔW$M3�7�*R��~+�O^�Fh����\�h�}@��Ѣ�j�>���c����Q�OR�+k��Q�5�k"�C������(d��g�>Cд����ᶯc����я~t�x-ZZqB��h\�:��f\���mf/e�<�WHh�~y���q��:5D�������H9����'��I��o�N��ߕO��Ǉ�X��e^]b�����k��n���Z���@�}�֭���u��#�O|�C�r���G��y�UM�/�Y���.28��p���
����Z�af��P;��5M�h���!ĳ��UǢc���h��Hyn�5l���W�,��M�c�H��h�C�7W���M#|xT<��﷡],�=�B|&��������O��gQL�W	h�U~�}������! �F�U[�#�=�(
�2a��N&4�5��8�!��;�GU��]tB�H�}�(`�nt�E���Ҁ���0<p�	�qճH9��id��Hy�wb�>���T��^�d�u�d�߹s�:��������������ž�>� �hHA��!�B`��Y�y��^�n�갬Ɋf�"B)ȳ�)�4h����F��h;)�'8c�pY���~	N�"*�N:C�4��(�����mW���"TG��<��+G���z�v4B7-E�42��k�[��_;#X+I��b���nP2y�!�����������_z�;߱S�f�9vG��������ޫ���=x�e1o#����cEͣ�M��E�ڱ/�sȢ�7q��4���ô��:}ǭ�q�1�6�q�N<�Β^ƭ��WV��V�Ol�I��D���wpye��;w��3ڱk��=������[`/3�JV\����tT��j/�`ϫ�;@[u�6�^��/�΍>?�z����2c�c4�<:�M�Yw�\�Hc�/w�� 4����('�>���Czn�t+{�766n<��s��I�c�O~�S� �	���!F/z�8�xز��e���u��Q
����(��0e�ؚ�F�C�ЀSdb�h}B���_h���<4��a(�o����@?��4!I������"��"���E�:=��n#��P;=��>�?����s���]���=����N��}n+CkP��;6*>��fj�E��4�Ni���#�FS�O�7ㄮj�k6\�7$H��3 ݺ�@����F��Lz�&�z�9dM�!�=���9��a3iuTy�M�8��4����/�tu96�c�{��ePa����c�yT�؊���P�:�xL^GI�fs��;����3���Q���7�L�_����?�NV�y|�т��O��xXz�	j3��y�o�}4k$�ny�}����h��o�~4���ñ:����������0;1�-3_���8�E�V,��*�W'8�1B}��kv��w�7�=�������Z������b��qH�m��c��=���0m��qQ~�{���Vi��k?6��L'XR�3�~�z]{ff�����=�u�cմq'C��1�g#��<y3H��wBD��kÅ����
�'��ZÖv�=�F��K�@|^6^m,��\���jw��R�r���ڭ[��[׬>��O�D6�^�
C��z�4�`�2b;gM�Bv��nw�x�b�S^�ci,�V����7�b�t�ɀ�O�)�����2�·-��ڗW��C:PK�A�A(�����}���yy4����6���ïC8�dw3��j�<Bt�@�g�Е�u��~�N�O��b�nKJ[$=ёA�GL9�eƤk�����	`^����G��WtBX�� �-��Ky�,�<Kn�|b�'�\��Ӥ�3�>�e�r:����2�h��0���|�?V��ڣ������֧����T�ht`��u�m���4���
�G��,��H��G%̣�B��SV^�1y�9�2�E�5oM��	��Ֆ��ݼ�މ�/��}ezrB�G���u2S������v|.�|	h�A�>��?s��tg��<xp���o��2��@�;�0u�YZ��x��Mۗ����i�	F.�.�>�?�*_��B�d,�Ķ˵��� |\��0}�P�4��,M�t	�K��B}Q1���d�(�"��J��d+*�J"]�|��������ڱX96M����_��?�g^s����n��">��Quz��k��!����;fF��麂(4x]mC��lM���5��Hk١w�E4)W �ލ�"�ꯢ��M���F��KxԭK#4�kO uǈ�Ō��PxX.�Dˬ�+m���w>lŴ>�3�'-�33��U�cmDB���|�����8�h�5��1 t\�kV9y!kv��ȗ���,��1E�*�f�z��t �M��ȠԀ�ǱeƦ�M�b�r�t1�����+�b�I�ˢ Z�_���Â��ר<l�|Y�v�m�1to�4�ǂa�C����[玫����G4�5��д�lM���`�M��Z�l}���5"`���jaU�����gp�Ae-�]o�i֚����.o^�䜐� �bY� Y�"��Pp��F ���Zhd�X���#[+�i�R7�WBu�K�Nָ�ϲN'+إ��[��MY� ��C���w��'us=�C���ͨC���oG��1J��EZ�eM���������w���Ї>���7�i?���}~l����~v��0����a��O��! ��5��5�_hr���lV����K\c(��1u��>�C@��;Y��г"ڬ[� Ǥ�������4ҏ��i��������յ�߼y'W�V����_z�Z�hܧ��H��#G��N��(��U�֙�Yydi[!�g�Y@;h��!�����Gc����M(�a,��I�T�uz�gHs��ݼ]�)*�:�M<��0��Ex./O=.c&-E�~Ti�v�n���A�ٍ��~�X<ȏ������o����WMLL�� f�G�)�.7䲀�0ub�pgl8�,az�'��P��OLm�V��l�~!Pβ��y�ċy��ȇ);��X��W#�� G���˫{�s����O��"�r���G�Ci�&1zR�(_��;����qԧH�C|�eݨ� m9kr��G?��2���а��+�!n���jLY�>���g�!m,4%o��v�n��"c�M��	ڮ�o%~,��1��ژ�t���[4_zв�]�/5���UD���/n�Ɗ�&��& ��;��A۬�g���l�<�6e�]�<���O�G=�E�h�QO ��;�a಄�q4���j��l��o�o_?�c�@�*/f���7�~�$lV>��u�,����h�yBO@�P�Т"Pse��}�wPɳgM| �+˥OV��~�KY���>��>|�i�v���e.�bM�XN�:�~���FШ���}��X��F��:x��5Z���/伂���(��1 ����&r>��'�c��4�koщel~y�P��Qi�n��-kl���l��4i������4a߄�)��<u{�d��������H�b��]��&^>�CWL���M1Y�} e��<]^[_?�m_��8e�=NBi|6>�9c��%`��YB'4�����国�43߶2�f�X�1[� 6�|�i��;�>���z��������?�*�;��y��Ch� 4}y9&�脦�$�:E� K��M+9�Eq���+z�3�;1�Ǘ��Wy��n��Y��(V�Ǳ'�>�Bꋘ��s���\i��^���X���nom]�����o��o݉�i#���G~��;��]5��d��4��c}V�E�o�|����W�y�uڍjP�Ɣ� o��7��U?��Ϙ�
MZ��_���"u��n~Y�y R�-yy	��9K���˟>�˚e��u�ˉ� |�ͅ��f�Lw<���xg�T��ѓ�m����j��piyp���ʍ[�n���Av�����ף����8��X���,�R2�?'-��d_�E@/�� 6�A�d��=p��/r�ic@���+��*ߘ~�4Y�~l;:=]�u�}��i�%!kR�'
��/���fl�Wt����GC�Feu3��`�` �Z��ܹs��0===�B^�>�f]u�
�<�1d�(x���b�/���" ��X8�>!Z�ip�b�X�hVyE�i��5K�����.�4���&Ԟ�v��~Y`���}ߗ_^��B���@Jߛ sf�ǳ���7;���#}^Z^^>�m_G�/��sC쌼�`�����:�(�`X�����1�bA���<Aۦ�|��X3�*R�aӶk��n����>����'K���к=�ˁY4�ɍ�	q.x7�A���/��0�����1*ڑ^G���ݛ�6$�Y���\�Q���A ����<��cN�:�`1��'�ߍ);f�7s�*3�_�<��>-%v���a^]||�%Ě�_h܄�k�����;A�	�F�ua���,��hYo0}����+n!i�y ��^V���nޤ��Κv�5Aˏ"tk��b��A_8�w�#@{nn�\_��h��b�;�
�o�@��L�Iq/w�Ch"�ռ��Y�tn���fd`�ͼ~����� �l�֧��E�nv4���Sh��&���B��"�I~�q�n[C� �=q��!=9z(=�� sDQ�S�D�d������w����7�<��<<��P__�MfzAd�<�]\\�^��{E�?�"E��I����?ZYY}��ɠ�Վ�*j> ��,��*�e�f�m�y��t����~'�vnY��i�麸ߣ���5ҞF�	r#ye�⍘�����/fL�{ym�yo}�u��`�Gx�&���ͨC�΍���[��s?�sG�u���O~��8~�hLy߷_�Q��{.s�3(�-��|n}b����BF�˪W�bߏ����/���nD@4�N�e��g���h���i�Eʕ�yZq���k�[�F��{�m�k�m�:�h����8���&2ٻu���.'F�m�o[�������E�>�m_G
��?�� N����V��/� +6�X�
��ͬ��ֱ�<L=�x)f��"<�JE�jF}bˋ5���K+��H\�r'.�5���R��}��מ�r�.֯ ���99�_|tg�|��8���L��n�5/�؉a�;Yc��hPR/���G��G���۷O �/�!1f�"��iC V����x��o45-�~he�ɛ�� &��F��z'4c�q�tѾ>
���f��;��cq�z�4�`�M\Pѿ�mH��;TN�W�&Y�mDf��y���2��7q�=,��x-�1�����PNwg�{�k��I4b����WtL?����1�"1@��$���^�&����^B�bhތIA� F_��u�ʉ��f����m	iJ��,0ܾ�{��ɇ��Fh�H9B_�}�g�RG����1�7
����G��0�㶯)DE�6�#��L�����=�o~���E�iv���R$4P�����'hb��4Y �n!��������W^���kw�d�D1}�W^Q *ʇ��O#��W^�,�`޻y�c͖. �𱏧C�������������Y��u񍻇�����Ae\]�6혽+!W}�f���i�Q����U~9�**�t G�gfgg�9Guh��C����������Fa�Ce�~�&�,���X0Λ\HYY���A�+�Bv��_���)�|�{+��&!>ͪo䚽�*v��$�}�Zk�f�8}�i�`�U/�G!3ul����>y����zi����+ϲ�.mv�9�g��DC�X`}�L��.E�,1<�E�<9.���P?�	NL٬��@������1mj4͑�������?���C�T��#���'t��(YyeCH0��Ѕ��������+Ү�I��/������a�.����n�y<S�&v�w|�i$w|fim�v�Bߥ���<4e�B֤$Ds(��oR떓W'/�[Aa��u��^�=�2'�w�:�h�ۜ�y!_^E�F^��XD�q3q�����K?��?��W��_���y��#�g�yz[�.��^N��Ⱥ5�,Pbc�p��P:]�,�l��B�Ė�$�SVL����>:��D�ve1h������y�u���:�P��E-�Gt}���N�N�r|}�0�����[�Mt�d�cY �,����[~h�f2i�U���ۀ�*��^g4� �,��1���}�9F�9�J�����B�YpbT,8Ǧ+
�Y�教�\�%�B�&��c4�<��������;����%Db�+����
i����1�H��4�P>�u�y�<���P}�r�x3�6y@��-V����wxf���ݼ��Ӱ}t��O=�&41r���D�Ž�PT������++�7��G�+��Ao�"�3��1�Āc��	��	�a�'PC�4B��w���,����@�D&O����
����׆�<\!\�w�N� `H4_�4��6�&�|?�}Zw�Ϛ8�������'�B4���!p˫����ɕ|�x�vZW��*�i_9���7 �ːCW����A��sE����W��_|����zl����aL�R��\Ј��
�"�� t;$�� 9���z��E�מ,`ͣq^=\�,��3�y��L�wE4ʃ^�Z�Ƞo$�ڒGh<f����F�P4�Ƭw��Z�m,RNLcA3��1����^�^�ɗ��s`c��&&_�l&���E�9��1�Ms$������e�W�G�>`��N�ʚ� �4�����ʖM�,���w��Ȣ������41 ���Y@����oщ�0��==(���'�>88XZ__/��e�S���=�{$�wn0�D�!�0�[s`��L�`}t���~������:H��!uay����܇x7x��Ǆ�䳽�m�-�0�a�b9��a���v�4::b���민�4�����Jy,������|FZ�L�u[4O�t#o9��,�Ӷ�
6�6�@[�Ų�<MO���}ȑ=���?�#��ýߙ���U���������,Y�.���X �J+��DP��|c���e�\Pr�_��;h��6e�(k$��˒Sz�m��K!�2oR#r�e����D-}~$�ܾ}gz0��#Z���똘|e贾{|ތ��O̤(� ��ɚ,����������'�P���ǁ��|��F��[ �0������%�(�����6�eRpY���ja���{dd��O ��R� 
r�'A���>l��%�����m�n��4>>��l#Ͱ��v�s�!�Y_g~g�5H����������/���ғug�9��dC��vɤ%��a���0N�L}��u�$��m9R��c/~�/���J��5����۹�;k�1�I��Pz߸�K>�⃼��'��%�^�)'c��x�z?Vdԉ�7o>�G�F�������\'d�c�lh5���;Y�8��N'����!d���y4����� ����[m�
l
a\[� �h����F8oo�0+X`���0���Y;H��m֝���K%)��̲
r��,W��KS�`٦��Q�rj�8�א���dagg� +Ӱ�EK�����l�'�)`�5R8�'#�O�xE򓺱=��W���E� �}Z��35���C'�?i������[U�72ƶ{oo�t���ғO>i�}�S������O����c/O��76B�;v|Z���V��_!-��}��}ǭ�K�W�����u=�h��7�q�+,�r�omm������S����z�H>1i��776eC�G�7Hb*�&X�:��58�&������*�W��>`-�|�Ŕ�������}C��h�,1�S��C�t�ҥ�_�k��/��,!P��3�5�;���+/묽�v�w1 ����KSSS������0 ��y��͉&(�^� ��(�M�&����.���/7��	���P	!�K��GLY.\�wx\�A� �I���d�=�y�����Џ�_��_�����
����"]�oKKV�%��O>����O�Μ9S���?]��?�#C+ҍ�}@A�'`c����|ݟ�z�XS\S�1@[D�����"y�Ȧ��̛t�Xh�>Y��Q�����Hy�4���?k� V1ȜAX�n|�s��L���t��_�����yEY�Qt|��0���x1��^�|B�-i]0�y���C����&_��^(o]FtBtqi���(�E��;�[
�+W���_�@O�8Qz�;�Y�vń�w�ծ߹�����D�&���}����7��LΝ;W�5�t����w}�w�:��� �:�_�^�������������̟�3�K�@5�����+^����;������U��i�Y<,/�ׯ_7e~��.}��,}�C*���a�����o��o2�b��Nx��/��x�Lqla�կ~u�o��]�K�/M�u�uK�ܓ	�7�7���o|7&���j�vYD��=�s� Y����gi����o�^�h���w}���� �O�d��,$ǲdFH�dɏP�!�Ȣ<���J��2x�q��\M���i?x0M��� ؈��h	�1Zݎ�û�Y����m����cwV���c�+�$q�"/�^��׾����ۿ������5�}۷M�?���l@]@!�T���e8�v�Z�w~�wK���C�Ԯ	�Ԋ�~�h��0P���oP|�p3:�������-F��Z�)��MLL����8��������W��`�N�廸����=B�~��ݔ/�|�Ν�e���_��9o1�������߀�`�iE��ו��f�7�7����Ī� �g�wA�,O,0�,mm�4
��L@dIA��*�g.�����i�Ǖ�~��&��Y|t�Y&|�s��㇬�=˻�#��1Z���!Y��(���)J%!+N��Cw_���o�B�}�tІ ���u;3� �D��\l������ab��/ 65-]��A��=Č���&Z�ꝧ}�MjB���&���x&K�������������7�~�gά{~���-����|�o|c���`�6�s���Sԗ}ٗ���؏��mo{����S�o��opoh�<�~���&�0G�.��Z���[˴����'3ͽ{�Ʋ�r��{��
�$����|�7��N|�&�7n�����{F�4Nt��w�v@g��h�~���=��aO@���l�,_�^�֚҅e������k����u��q��y�s$��偝+O�~��� lHN��{_�!�ƒ~�E -4��M�b�yeq�KwO�~�0�bKl�^�v%q�:8��hgq�fl���X;&���'��0�nLX恋O��"��5`C��@��ն<Pt�j�W����I
>-)�}e�z�s�+ B���F�*���x�~����[�j4����߮���!gՑ}�r�F�P9�U�~i髿���$� KM�k��/�6ʵ_j��8��E�B����1=߽z�j��ݻ�tL�f~Y�z�z�����oh��lփui�ܰ#����O��O�ub�C��'?�Ic����O��OV�J�v;�����=)ؗ������3�����M��V:Y"���M�y�;����0Z���3�o�B���n[5ȹ�a�1��/)��6Cګ/�,y������`�&.�B���c_�!,�eW�7TQ��٤7�R��.�����]��Z�M��5Yq1���k:h���]� ��^���E*�̴y�������y�������' Y��X u���E@���Of_��:�ګ[L�\�I�e������:)ͼ��	������p,�mF��Ϯ�Ǽ5��pg�ӿ�w��q>#��������7�(������0�M �i��\-Nӈ�ؾO|�@�������͗г>�'ΝE'�,��G��7�k�_�U_eL���<��F&pв�7xMp�)JZ2�H{�����1y���h�&ܱ:�F;~����i���s/��f6�����[پg��1_Ҭ������B����=���z��1��8���}_��[W���x��i�uǦ��}��h������~ϝ��2��!����q�d���eL�o`b��`S�њ
����w��������Cm�i&�6�W,X�f�_ C��0�q� �m	�P;}�}��ڟ�NW���`C�����^����{�J�}�{��zt�ۂ���`�h����cn�鵶�jǀ5C�Y��,F�������~qm��n!>�}��Dֺe����Ϳ�7F ����і�>AW+7��,Nrؖ��~ڬ���l�b޲�#�r����/�w���ؽ�\��׽��p-��}Nx?h�����vV{�vVu*����>�ӧ� �c�6��|��Ѣ@S�w��)�}�k��v�i�n}}M7wr*+o2�GWS��Pi�.��M,b��ʱ��aZi������˰��P�Mg�T���g>��s'i��@,p&]������Ť���<sA<�C-�~V�B���w�<Np��h�)���~��+��+FHdO�<i@�Q�d}�y�sH��+�Z�D�	��E�`̓��Z���2�\Ĳ$�d�_&bʵ�Re�[-[6`�G��|jڜ��3�� ��	g�I�	���r�#��6V��5�avw�^v�&�5Y��=�l&��$��o����		B*W��ъ�2e��m�\��,Ex��>�yZ���]���$�'\��*?��$"4� �����K�%��*P��s��+����������r���[� h7݃������C�]�GBr�mֻ�ٙ�B3�< �G���3e��IFpc�RB�u�,�'Ѱl��M e?�6 �KӨh������L@Fʦ&J��ڜ���Í��.N��e���b�eH9\of��|E[2�E����w�Wk��wc�i�S�X$���6�³ ˥��_ߐ�t~�۳�\/��q>��:�D�S&N�[k9hyM�1	�̏~ 2����in!����_2Q
�~Ǖ->9�;�C�̲뭵�>����H=I��r��֗�k���=�����(67]HV�}#����S�0x�4��F�\1�IWSA�֭�SqB��&յ)�� cV�X���3�!���}߳� 9�6zP���B�H[]!)�ZG�-�i�D�t�M�ϴ�y�~rK~���!M�
x�b:���#d�O�)[��x��?�|&{�m���5'��N�$Bg�Q�X��%��L>��`Z��S@Y�E�M��8		[oV�yz�`wyN4e���Q&3�O"�e�g�<�9fi�:_��`%_~.���zG��Χ�}��E×�N�e��1�����_yc�ZG��L��=F�U��W��=__�r]hB�q�S?	Kc����E�7�g�f/��z"�ƐC�[ټ4L伤K���|��q�@*��y ��|�X�=�yB�c���1��`�G�a����uF�t�'�9��V+Oz�~]Q�S1��#s@����=��jцm��\x������%��|�~;;<���ǦCۦ�������:V���0/��2_�i'�)	���7#���z��gn�#����˰ö���
$~x�o�&B�t��4���Y��w,�ZDl�+�;3[/]�>8���حaY`S�3{h�].�}e�R�^?��0���S��� �(4��tF�W�h��D���IG�8Qp�Us��УF�}ڪ�F!-��������Y���˝�ԏM�ړ*�*�Tm��tM�e�X:���t2�UF�d�[H�o-���o�O���M��i�~�"�����w�VW^E���a�tv�8�����S����c��{�<�.���'�	�@�n�~�m[�୯�x���C[�*b�|�O�S�V��jm��nESs�ǝ�h���[��/��F�l-�������aڸ��:�Nβ %��?<.d?t��v�����>�<z=���R��J;t:�� �L�jtx�>��'뎇��ö�ퟘ��kw}�J��K���Q�n���h��<R�[�o�ǉ+;\^����ɡ��B��'��d�~�����xκ���oC���iv��iO?x�u�ҫ��dl�>�iv��bL7�F����BH�貘U�'iB氬Ɂ��d!��yB���8u:�[�G�}WɌ�a�v�7X��k��=�2*�j��'3k?����%��'3y���_y��C��k$v՚�X����?T��_���Ր\��i��o|Z�;1�ѡ��fҠ��������ͭ�U�4�ʷjqU�"���X�٣e�CZ��N}r+�kZ�r�GW����]�7K�RV��Lޘ.:.�����B`�hm��!ihc��0f�7�}��^xܵ�C��Я� I3�f�0��.Y���&潬6d_�)7L}����>ڡIP^9EA;�<zޑ��<�UY� .?�1�qp�6�I���`�UÞ���N�a�LVi.ח����j�h|�[���~���1�n��[mڽB�A�'Wܶ��V����;�����/�ǲ��&T����p�*i����ON�z����7Ii�N.��^hc?�Y/c�(i=І��*y�j�0R�7J���5�Ny ��>����}�R|��;n}}��W׺��L��yכM� ΢�<��
	���k��y�am�$��1�_�Zna�rY?�)9?�i�a��#xS]'�^�l��Y}9���.x�	��:h�<�����+>�vi�A*�!���8�+@)e	����P��������KG��)�}�,i���i?v�֭�n�j���>�? Ӹھ�;���(��"������d���E�vq�jS���kg-�m����&��C��h� !o2��<�	Q��"���q�����ei�n:�/|�p�����ϢMx40շ���Єx�Hz�g����`�,��[x��,Kj��C���1�$�7EqE�#�_MG�8�	]66gY��e�+����{%l�DjT�����EA�(>:d����Y�^��
Gw��h��,���,�Ԟ՜�Bu(�!�d呥��m��rw>��,�ޚ�&>�	I��h����O�ɒ>�+7\�����M |��>v����@���6�/=Aq���G�]wR�e���4�偓�{����͝$��%�>>����,9|��s�<��tL�2�j/vG��価��d�o
h���q���&Nq+�K�,℄]���1 �2�;`��G͜���i��+G
�`�^ž��h.H���}�w���K��o�G�,��_�C<�Wow��d���v�sߤ$v�f�f.�d�����1@�C�ʘӓ-�.�Z�I��\��M|c�v�:���*�{����n�r'܉`��U{ݼ��b�Z�s�]��']�x���q�ȥ�<����:OO��r��7	1�e:�k=�4���0�k����pB/�9�2_��y����G���8�qV���"���	���CB7P\A��1 8B���w����ڤ���Cee���8b���^��Ŷ�'�&{K�[�o�~W�P�m�	�-t�pC \���±�����������\<���gQ�ǭ<ƱC�[�8���`7���v��uE�2�ˮ������ؽ������gmr�M�o4��ͦ� ���)?�jq��xW��I�*��#;L��������lS�}5����h�9�A c��x��vR�`��! ��\���?�C�:�Nz`�6������My���^��/n�|�}ejZ�h���߾�!:�����б��'9�'$��I�.;,���{(�����&���ҺX_	2�+7O;s5/��.�;��z>�`/:���߭�![E-u- �(]���U�]9�¥Q#<��g>�����W؆���'b&1ulF�\���}�yIMm��O"��,��fV:O(��
���j!��*!��,��.X�LS>�����c6����-:�/�m�X���ut�#m�A��eP��d��g�=>�۷����M,����;����s����+2�B��T�.�t?��6��	��x���D��Wlu=��W~t}yg�����u�i�Z����u'�/���׭���C�5��<U?I�{˻}&c/D�P��������k��.�mmV:��l����?���o��o�jF�Mm�?��F��T5�6�z�������Zh��|@/i�^Oty�-���
[)[b<K�|��j����~0YЖ{!��w�^.X�	M�,@��/MW�?��}�|��f�PR��>䫗��q�?��&���ٵ���ͥ��&/����t�B����a�'�v%�~l=9Ѐ(��n�Ln]}bn9���)�r�M�����Ld�{8���N��,ri��D-75�
��zf�+/|� w����S��!��g�
<�s�5@�����z��?��1x����_nZx��[+������f!Pu���[��+��P����-�7yp���rA8����t�T�[=�Ȣ�5��~���H�UM Y(���6���$���}���Hh됛N��W�,�v�Ō��4�=t偰h�Y@&��@2�n.��Q����{ǥ;��z��]`�m�y�;�-®B�+�7Y�t�B�	�jZ�&}���{��ג�n��S�	M8�;���]�b?�A8��U�� 
W�К������ex���@�5Bfx�98���Īl�|��V#����S9xoPֵ<�v#2Q��U~׃Q�����L㚒}tO���u9!S�~_�ŝA�m^h���>�_�&6p�ka�7��ж4��}�Oڙ��\�mM|������K+j�`����*/:N�5R�n�l��ښb�m�i����'H]�Û.�������i���� �;k@c�Y�������'���ߺߤ�G�˛���@�=-#D~h��$F��)^�|�L�P��ȥ�𖌛Z��]�	�	χ'Ϻ֎�{�k�Uew�n�z���*e��2	`�Q�����4Rc�O"%t�ڭ�򓿴�W�� >L�B����I#�;�&��������~���s�����s�]FH���ꜽ�z�5�s͵��8�[�r[��2�#W���}�<^0�������:��}yIm��v��MRl�O.���?Y�q<�K������eyl��.����x��tt�����#cc.ߘ��iv��}gΜ�n��x٤m��a ��Y���|�!^%��U[���Ej���ZR���%E��c���	)��X����^��f���;{^��>�70�u�dF&�#e�n�-�n���p�,x�බ��p����e����_�N�d\�7�J�d�������ѕ����s:w�u�����y��ۂF����㢫[��_�-�ЧP�2�2��+�#iq�m�j�W��漉r�C�8��,@69�b�2�B,Ruo�����0U����N�C2���Ő��)_�,s2���Zk���)�����%�}vv��*k����%���{`b��-h^�;�����O�g��p�����(N�1����'m�۱���3�iK)ᢰ�����#�y���Xɔ��}��x\�XwS�a5��P�P�ʈ�O�Cl\9���?7�u1%�����
[�h���Y�u���C��_QK_��C���_�(�r�V��V�ݨ�NEseL�F2A��� |���!άo�B��F�	b^�F;�\G��Oo���oۿىn�A��b)^��qg�g��~�=J+�>���9�:[Q�y2r���Т�-�z����Uf#B����K�t���/�l�~@�ҠH��m^����0)��v)�H;F�[?s� A�#��
���GmR�T��oJ_�:�%H��nQ�b}V��;����J�Hly3�,r	S&�n���c<E�L	7]3�W�C�P�1`�Ԩ��[Ks���z��!�����j�<�l3�-E ��/YF`z*6aKfԗ.޵��������alv�q6�тhC���n�!.�W�D�[9�hJ�Dn��%EU�/�u ǲ��V�8��
"ӯ�ŝLT�����Tg�6:�5Z0[��QI��W�����]�,��1n����ׂ�_�bcQ���\�����c�3m���
�$�#Y��,��}������n�(��nY�Q�΅}���Y
���u�z!w���W%�	��Q�1m� ��5j�_a	Mq����}�֓��H����a�F�Qkq�����h+oR,��l���673�H����u�[�;�!@����k�/|V��8oppq�<��bD���k()����E�̽��a8I�9�k�d|�rw�a�����v#�9���3�L`���FX�����y��M�K�p��5�M+]Rh-�~^a�r�� 	y�6�s mWO�P�Q)>���~yBvyW"� �vx=9R��QP��:(��~P"ˮ�;ϥ��,�����#=���e�2�u�=�pd�R��}�>0S��1�K#k
��^ږ?~k$m��'��u���]�L�hTv�q�JƮ��e��|j��CX�:�2��Tw�fz��ނͧ�p:0*e�0ru��v'�C`�b�/�m2K�l�)Nc�~��-�NO�WXCLH���C�/�M
�&�2��S߹�Q����R��L����6�� $X�z�֨`@(��-�W�V8D�m��.�Vjş�&�^F�"c������*�0��*���ʗ�C�.vwq��\�Ņ;�4�6iLNe����dVS9�Y��q�owͥ���hǷvƞ*�]4� �t��P��uF�Q?�`�n<���d�V&�1"+wA!B�h_T{�O������+:�Ӡ��Ƃ�F��A=ƈ�˜1��oT'bt�
c�YU���k�(ZB�]N�{��#��z2F�ֱ���@è#�n�~��=��X�''"�rĮD��>��T]bЗ�hk�99yx�`U���;B��4g�C�i�m2{%%x�1y��a!�D�i�/Rd?�%�>��{��G&#�R���r��~��i�g݌�U����0���zȠ���B7:��6�j��(���r�p�W��K$O^V��V�a���`�a��F�	�?ނ��;1�S���ӗ��%����y{xA����N����0��<�5����H{�^�6���IF������3{⾯���U�%�+B�]�w��ym�j�	�j(��4��

+;.���+��!@�vm��6P�a�� +���8������>�������9y(�k�P�a`�N��b�(�;�̾?F�;��AGM��шZ�񔘔Q/Ʋf���u\&ed�1��`yV������H�>����6��;�_�h�b»���(%�	`�;(kD��s�K4�VJ�	�g����[(���� �*�k8(3��-��d�I#̛I|��r�V�j��H�u���:�E�{N���y��S���Ü	`2�q�!J�Z��1�FB<���/��๻'Κ(��:�j*,�5o}����{��==0�j�+�!ڸ`߸J��Q�=_�uމ]��U�R�\��P_|�_nv
�6.B7��_������kp�~y�4Xv����FZT��r2����W�� ����h�2l[G��ѱ���H�>�%Ƣu|h�3o�z�w���c������c� ����W\O�{Mm-�3D�beޟЌ~H���3�ZZ��mB�i�����|�"ش���V�t������%�{��r�ζ�{-؇j���q��?�L��9sd�?.�r�}K�Js'��aI3�ϟ(t[�s��a[���w�b�������F���`�o]��}�o�u���I(㰊i6)�o�܅b���3��k��؇�n�\M4;��3
sìU0�I��s?�H�kfЇ
3�+��e�c��@ZX*-�Y<t��2z�'�h3k��Z�19

����J�É+Nϐ�b���Q��m�}(%t���8�mc�;$�s_C�E��K��N�Ņգ�3�ӶV��5˾���PE=Y_�W%�FmBF��hDݧ���ͮ͗K�Y�nY��)���
���R�5w�a	��i�O�y2�f��V��f�P�'����2[:y�W�gn]^����.+�|�/c�Q��U��^�B�94�_�R�����k��ȹ�<�O#=tԇ�:N�H_v��(��5�(�w��78���r ���\ZŤ�w8��bf�����8{�AJf ƒ<���8�!��|�Q۾5�U���!�'!�H0ڌ ��v~j��ӈԟ�)���޻ɨ��:��d���w͂�~������<Y=�'Z��%W��9E���@�6�->#�����X��"3����@���S�i�� J��/�L�!F�`J)�MJģ�M�B�}h���@^��$�L����׬[��^na��uzl�W�����?�6Ja.ņyp�,W+�O��k�_�X̡��4�0WR�������_�~mX�LR4�P�i(d$l_�
�^��+g~��oҔn��ʌqr�v^��Wwe�G�Mz�5D|sʿ�j�Nj�^e������A�se\7̈́7�cWOk��V��*0���=pV��2[�}���,ڌ��M�9,B~2���=��Z&�@3�}:% 4�!Ȥ�o���0�Vl�����z'H����w��-����C��<�bT�����r"��F�X#���q.9�q����%���mxr�s�|���]���W;��$��<=.�6b�'����^��?���v����p2� ��V�$�H���P�}���y�#ӣi�����a_�6>����ae��B+2���,4zr�$���m�lI�$L0B\��/��ٍ�-id�8�����tCa�ha{���֚6���3I]y�_,)�_���-�R,l�s�3�����f^�ծ�Ň���N�������K��n]���Fx�����r�UAu`9I[#4�@<���h7<�J9�'R��ÐFMgk+�|�re����P�����hjS�9ŽY3'k�.6��'�U�j�|�yN6.��A���g�D5ϥNM�J�A������cz�9�o
i��-L�ofX�v���y���N�F�	��ax�}i	&n��?51=�xkp��h?L�5*�/�l2|N�w�=9sOi4�[��Wi )Or�M���=�-\|��睄�٢�nXһ�*ԇ��B#y���95� ���ч��T ��m�р�l�|��?�zol�6=.��,lY_e�\��)"&U���N��t���j�u��*5���E�
��>K ��֔�!��j��<�����0��O��['v�4!zN�'^�݂9�.����Y���dT �z�6�2.-}\�`�ڨ�wx�f�bH��\҂�FH�5=pB��b�X[�+����+C̶v��8��������?h����[��7�i+S�BX�wS"]���g(IYi��R�]��1�.4���\�;�ӱ�^����r��?|�#y�i�@�hO�����iBW�>fL�1n*}�A=I����e�}K:��pw8���l�+A5�<:r��P{�.�� #$��k[�\-²�_S^�ĂedD_���b�؜�Nh�:U0=����]}�ǙL�ϓ�*�x(��me,�x2f�eP�u}��	\Nǟ��}ؙ�ʪl����:�诂��f�&3����@���p��{Q�n�TF��+)�u�Z��X����_w�u���R	�[n��]�n���9�֮�����bj�+UQ+\�>$��g2�S�����3F	�<^~�9<Y���-a6���O�0P1�h���B��/6*!V	�9")a��6��GN$���^��:��B4�C ���F	?$M��A��s�hz|�P``��_��G��z������oT0���1��Mq�у<We�R�W'Q����t<K-�$�[T㨒�����k������I�}u>��	�I���H�M�=Yw5�Kh�b6^��>�I�͙�T���Y-l<��Ä�u/I�mڻB
�g�UhY4N����R���L�S�4V��Pa �#<���w�¬���ʚU�-:��l:#���q�`f�3��ן��y�~fR����v&��#�=�+�+c�>����ϝ��r��)��g��$7x���oJEh���]���Q�	a���Ђ�z���mT���f�'���|��i�ڑ+�p�|jMs:Hw��Z���"�g�>~�����W��$i���g�*�)�x��H�IK�x/p��V}���x�V@���]�!ϸ�s�����{S֚�ܺy�މ9K�!R|O��*���J�;��$��D�:��U���-��=�Q:��v1o�{i\;RL���_�vK+��i��`��#��mIpq��ƐG~+��/]�g�Ґ���ۃb��& � ��y���1�� ��_�&4�EE,G�\�i|�26����hwç)�Ӳߛ�Q�f������]�3��n��+�|��P?��Sb�I�bNjȃ# �����dʓ�|�����"�8�A�� �g;q���&�p0���]g/^b�*��N��&�>���)k� �3�@eȏ{�GfJ��ZN���^f[#�}�I��;OV�,w�oGfK�G����BB5[����䁟�fҎ�G�Y\�?��ꮬ��M���p��3cF�֫�+˘a �~�pK��;��p�6�PP��2 L�peb��ǛuB;�h�����MB���Iԁ
¡M���f�& �kPz�O0M�������G6�ɻlM�`��ŷ�VðIkf��
���f�Z�.�x��WYrf�b\�2_;��[�f���s,����q�3�6vY��e��K4���	3��^N8���։�N��QwK1j p�$Mp�T:�8�M�/��c��_W�����ϼM��]i�z:�� �<��F�a��RI�b��"VԂ&.�`T �)r�I��>u�×~9i�kb']v\\v�a�
���(��88���Z]�\���?�#',��(���U/��ң0��b���m+�0 �7�Q��$P>d����t�y��\��GI���i[ f�jʇ��F��8��8�c�}��i��O�!��&�we�h�6�dA.3��\�tx���g2�tOD(av�1��O�
�e/^=E��gw<y�Ģb�����}&(��*�.��B�%i�-Hi�e���=M�Hm�dQ�	��]q�1E�,>㿡�_���ۨ�Q	M���f1��U`!���W�P�'$ '��c9�"�?^��'TL�<���5���7S����wBM�ߥ{���?Huq��1�{s�~����,F�l��H�58F���+W����1|����eP�W8J���zq�|Z[!�95�eT:Cs���1��L�������ɾ�_"O��<ۭ�Ô�/��os��v��a��0F��Dףr'-n,l��]�&�rңiE\(�ת�82+�ͧ��E�5(�g�.�1��[���
�,3�N2r���_w�7��P9`�	��8�'Y1!�Ej�}3�`瞒�6�U
�(\��&3�z?��߳ͅ�Nv��o����׿o?���1��b<�1���]9�1Wx��}���W�k]7)��3�Ux�q�	Z����'���B��V��\���'���d�?SO�9H��'���=�^ig8�?O��e٭O��̇$����x������<o=�z�ONG���8��q��P�81�{�E�?i������r�8� N
����_M�K��P@�u���
�^э��T�:r��DS��9���^�0�$ʶ�ھ�n��w��c�Pa�d��DTܘ� !]t�pv;���η��#U�c�N�����~kn���V��.Qf,q>�Nf�[3�iF�Ǽu�����x��
������sVgb���� 2�P.n��_���`;k����K!^�O�]�g�d/�T��>�����!� ��������2��\�w��L'�W\�ݲR~͌�ʸ���H��hu���]f�6;i��g���kz�3��簮��Og%��{�!�sٖ���>���z�Q{�v%<Y��V�
s�Ǒ�ʩy���O;��8���<]Z"���q�!���9�$����8395>�q�����yF�"~UA�w�tQ+�<]�
�Y�K����ZH�ŉ�q��%���S秎ӂVb� e���^�F��9�鏏T���$���E���=eH��be�6���t_Y��Ðwn6Jۤ�+�Cg��Ոi��8�f���Řh�-�&v�1Շ'�o���f�({P�K[��J��'�B��3�{� ����S�z��Cucm�*Q,���������3�o�T�da�6�W-kI�����S�.k��: �y�{�iE?�Ff_��BA#��i9	�!����	��?�^?FF8Ai)e=0}6*g|O��ң�z���>Cu���qw&�)]�D<]�E����Oֈh�+��M��N��oK+�|���P)����n`�"*̏թ}��B��)�����o�93w{�@���B&���%�'�T��v��I��
���Qu��4䰘�	����3ћ����Kѧ1;a�?��:nо�w�~R��i��Knz6��J+����	<����a�Tt�s���G�E�/-0�hA���3�	Q�������,C^>P(��iu��J�ǧ~�r�Y��8oVMC�79�_+��e�������Sׯ=���� }'ѧ������g�wy��	��]/O���9�;�'(I��I^��z��dt�>y.���/:�<�3�_��år�K�U�~f��Q�Yw�[w{�M8誧R���2�{^���d�B,�/��'ɥQ����x��p�����W�I3d:��r��m.|R���יE�,&<�h_^�z'o�ۙ'ڄ��G�%��rS�J�]6 ��[�B�L��+s��|"�� ��S.�*���־�૲A��7ur�h�ŧ7V9tl�3��2��	�S�v�6�*73�ԟq�]�X��r�����P�ɡ��P�[���T��B7�5�}��|�n-�qrT/��Go\p�<��^��q��kb<�֊�3*V��8~e��ۋ���2����h�7�;ա�����M��R�\�r���ke-��;hs\��I @9���=6%^8i��P��Bs��챂n	n����'Z{�L�\#-*���G>s�g�`��4h�������>�A����0��̂��V��帠T*�v�M�՗��~�99�1�fX]t���Ӫ�x���H�E���b}ܟ�Z<�>�'��{;�_���������
p���?޶v�:	��^}�Iö�0 ��azB&�]\�N�]��A���f{��d�L
M���_�ҧ�ɂ�yă"��1��3ֹ=vT����ʛ�=}�k�/6l�-L����&�ͥqd�OW~�E�~W�$$,�W��2᮪�Oʚ�p�-}����`-���MF����Xg;cLhst���4-�*S4+1{�+܀@���{_ݜm�6��C�1U"|r��������d��XZ�*�A���J��0��w�.A�zs�-����˟|S������`\�,R.��v�y�Q|��H�.
�8���8���%>xz��p
N��CĨ��F{�5/� ��>�x��2����~�*��X��Ogm��8�S㥽 V���f�GLo�%L��?��K�z�}���T�mU����["��ܵkղ���!H�"�&��&���ݕ��5ޫl迖��8��G���P���*��zG'�)=��ҥ�O��>Im�W5텼��]�⍔#��,��H��-ս�������*��_F�M��R=��{��y܁��y��a,���O� ���n
�yi`J��0֠�NL+�.@�~.��y�-��Ē�{K&[y~Ӂ�fܕ`�"ρy֊�Y�,.:��DԘhSs��"�L,���o&��G�����d�B��SI��S��b>|�Uh����I�I����16��t+��6ls�yЌ�4}��L���_����w:uS9�%�;����8��p6�[����Yr-N���'P����S�~/��+�No���'eP������4��-��&�2&���E4��ޖ��x�������8$��q꽡"$!8r6g��ck@]J��W����"��������,Ks�r��T���;�$��8oh��ud�$�^��
qn�O���*�_�2�ޥ����@�n���Q0��1o?w\��n�ɵƞ��l[����p����eSa3j���i*��Ѣ�[�}��z�Ao�Z��� |Ҧ��e��G&��c�5�1��'���'�Zό�B���1~zE��ft`�Æ��ڞ��;z��Ӛ2�ۂ��Lab�-����Ô�:x"�WEK�AF=FG�cF4�B�s���m��]���gc©.�������vV�fY�iK���ֲ��{�l,>]�O���]6n"z����� ���F#��2�s���҈�0O���p��aڊr��wn�ja8*���8h�菾(�}8���CJF���~����{x�|#Y/Yza�4;�
�4�Wot!)�X��4)|�}e����l�}u�Q�Ug�!-�L�3��J�� I��&3s�, �]��I��{��W�u�O6��֕r��&Lt~Vc���3�7y��}�}XG��O(�jt�H`n]>V���W�W#���nZ(�� !�8*_��]��y�H{$�&N0��Ӂѫ����F�/?��͡��Y��I߷�6�\�G�x�Y���q��{��T�ajK8���9P4f���:�-j��Ί>�g�.�	Q���4���8�B��2�}��1To��W4Ne�"�\�����!1?T�@�N�� �7w-�!�G�����&����o'�I�nwa�0�{@�p� �Y�^��K����j��͇�`���w&4���^����KY�Քl�|��=S�k�AT	3��W�j	�﨓+e{�ʒ�?��2��0ץN3W~��@N<&C�Wt��7��'����/kϳo4��n���#vd�L[<������w)ߐ��fr��l�ɘVvԡ`�{�1�96�]��}��M�A��;U���gU0��MyL}D?%r(����WaZ���ߺ��\*i��i}c3��ҹ�m�4�1с�'äe$�Z2Ґ�HX;2wG�|�+F�);��ώ��us���|��-Ljm�
y�!��R��]�b#r��j��!:E�Q����䊬�9|1����~�p�vjYѬ�W�Q�u�0[�d����l�D�s@��[g\9������12#*W��?h6*�f`9� �-'�j�c=�rc�]M��g�k�X�K�*�L��i�g����EQMV�_�q+L�5p�4h5��{���(U�t���?�y��Ф.T/�T��h3U�>�]RlW�N}�w�a�`�2b�Й	�����a����S{ޭ�^��\�N.F�UtF�o�0j�k�lW��p��b�"GGY��a�k�Aߵ k�z\aCT-,�����x�1/�=�e�F-T*�\���#
`P��Ů7h��ց"�U�����2F�nZ��I� �;��-���u$���^�����	n�����+�g�B��SQ@,�%�^�1)�J��23�D�jg!��HY'�[₰�d1Q��5"�j�f]QC���t�D��K���*L�:�PGh೩E����G���'��v�1�]4-n�m3.T�j3�qY�<�*$��zD�e47����G�~�fq����T�;n[F��Y ;���j�=���}1U����\�W1�w�7�,��-B:������6�N�2)��EJױTP��V�c�>�m��ug����{a6P�eJ5Ϊ\�F�Z!	pa	L��8����"�۬�-�+ ���C��(�����T�#L��6�F�Ԅ�#Grԯi�J��}z�E<�`	�<���]��c�8���s.#a�w�ty�gs�@@~�tNy���`�������2?�j�A���z	;}�G�,���O�� a��|ϰ:Z�g��������H�D���^��gA+��!��Z��*�xO�t֖i����)���yԾ��x�4���tu)��A����s`7�X�2
��_�W�51�G�u]��3{nM["�~��Ą���*_���:aa%��M��4wIw`3�<"���C/4q��c��ƌ{��I`:	�(h@�e��2��(B��Ņ����pOF�W��� �$��;(Z�w ]��>�]amϑ�,H}͛�%��%7��y�0���˱�yk�%������9��[\��q���f6�4�G��Vh`�.�t�yIqk�_AjՏ��(a�:¿�����j)����k�LA���W�$1�����wUzZ�S�9v���Xv�?o��q�QZg���Wan~�э�M3v*_(�ҰM�߆����17�n![g%�$�8(Z�H1�#8�湪�ad*�+�P�+��k��}��!:-x�lxmN��@_�Z��`GV_��p���⪀���iȩ��@��vP<2�a<}��yI��j�s�Z�,��7zaW���btmO�v��r�T���>M��p:#`{�ϭ��J�ڹ3�X4R���ѵ��M������ev�亢=;��74a�
z�PO^=�i������N����L�k��g�ۆ�|{_k|�C>=�$�k�_�Hҩ��������Gw����7��H��S�S���6�PK   �cW~�޴� �# /   images/51dc5037-8d6b-4f3e-a32e-636e17d8257a.png�eS���5<�[ ���5@���:���;,�������������ߪ�7��5_�z��^�z}�5���(�x�   ERBT ��z��þ}34�  �����K�������,�  ���d8y%u�S�}H�	�6I D^�$��gt)x�l}C[�Y�0x�0�0�Fl��0��oU$3(�!ԇ��_}>7>���^fq:�o���K��Kl�D ,Z9R��"�a�}�:���\��5 ��;:�A/80 Zp������{mUr�����&�2@�R���b�>��  ȷ`��op5�I'�"�.������C1#`1b�	�k|�_p��Ul��՜]�����z��]��"���|t�-\�᩿C6)�\�0�n?}�p��:�y�˘�����e���K9��PrY���Vv+�3�)"Mߋ��+�oU�g���R��.�ƖY�Z�1K�İM���"�{��ľ����{XLIHV�\���_{�J l��n���j�o/¶>�W�/am&��:�,�T��U�+/�,�<�N����c��*�u��s�R
I4�;�I(���%��%�-a�Q�=Z&j�08C?C	� `;`>y+O�N���p�y^"!�'˪����
�Ϲ�����R.���H6�0%q^�`K�d[g֧�}>E��Y�N�~%1��'@�Bj���|��w�@	�C%�B� ��A&����VC	�������G��Zc�BL�CcC�r�S���nM�O�(B=��e"��Ġ�Cu�Z�\�к<A�BD_�!xF(_�±�A�Nv�����r�[��=�+\�?�)�����(�~�6�L>���\h���mP<��F�g�Z*	���a��W
*��a���zr����~ (�����oP��B?��/�I5����A'�ɭ�?K܃ڣt�}�h��x	�ѭeI�ĉ��.�Kߋ�7�R����Ғ�5�N�=ԙ��U�;�eI��D�DU�Ꮊx��f�%�A��	�\����x�(�XӨ��$·P�����y���N����$�CL!���)L�UHMjNhNܔb��
S,�VT�K\��O�Rt���q�Pqtf����T�1Q1��n�Y�ņH��|Y�dT�TYd�T��ԔX@)>���LE�&!W��ߢJ�*�	*4�4�4ˊn���*�tL?�J��"�!R�i��?�)����ܢy~	+U)!(ȫ��o��+g�g��;V�L��Kl��ղ�zֆ�z�$YK�N(��_u_�>T���j�.|����4����Zc����$��1z�s`��V����p������= �/ϙ]�������N3�auӑi�ҺfƐ�oq�p)آ�.�(���L�+%�Z��TB�j�v��1�"������'��_��23%��+�m8����R�z���k�k��+�kqi�_Ȉ�x(D�Pԃ$�4���#�"��8�9�t���q?�N�_t��?T���o5��~�]�����*�=���0�4n�|*��\7��W0���P�P��~R{���ϣ�Wc��OW�q�v�x�x6M�P_Kw��y���r�8^&x�S�j�aѳ��Ǳ����ʜ���q��)�<��
w-W�S�ωݑ�/�'�é�������5�=������m�p0�A���SO�Cc������<C���E�����QVEFP%+�n� :x)~?u�iQ�$�������j����H7�Fi>x����3O��C�f���k�C�����U����%����|���������oz���qi�$9����?[k!k�k���?O��̟eϧ�����rc؉p���!>:2:Y�-7�vw%;���b#�p!��l�|����@_̠����u�i5���k��Q؜�����$��VO�|���ף�i:_:�}��(���4R�ϮH���~������ ��~&���+j��WO �#�Uq�a����P �$����h<'Z�K~B!r(�/��éΩ�)4�����	�	|�3\\���/���;qÌ��y��vCi��(I3�"�H՚v{ZƔ�_g�S5mm�6��H
I��c^U�/��2:46t7��tȤ����ޓ�86�7ѪY�c��(Z�`eZ#��5���t�o���0������|R���o�Wꇪ����_�'.&���_o�z��g��mV*-Ȝr]n)+d�^>p��,�6�����k�8�W��-Q.RV���[�zn�0%�$:�x�9��R�����i���;/<�>>�Ǭ,,��+�`r���<��u|~h*W)���9�:���=�:vdtt��C��|ht��C��:wk��_�;SL�`�F�i��	�ÁE`�)±t�����ʔJ*-� _�{�f�"�1�<�+բƲ�ܓ����Ca�l	h�&ȥ�lxn���l�|7L�uj�9us&|�{l������1�:���7?D�,�e�bwA{h~ɾk!3*Ϻ�o��A2�?�k����K�*4w��+������-͹��'#T�W|Y^���Kp�h��zD�|�޿��v�/W���m�m�Yb|�s}����7�:HY
��h{(S��^�c�g;�L:R�Q���.v�T�+�^��g����_f'f�3m�-��͖���X�S��h/�����T3�Q�,Ypb8�<���_�5��p>d&p�#f�@PQ@�� ��$���B*�'���,���Lt�M&	+��<P���Uw�<�z�5�e�Q�j��ۋ�S�m|vK=������K!�������a���-  ����E��N��#�,[
l�-j���/K�z�!���F�HLw������+˙�xK�CL�\��\Ց��e��9���)�į[m8\�+���*���"Kȃ,�x��y�}�i{ɞ�?��������o��0A��P,�A'-���&��x�	��F��ϭ�����}�&�~�|���W;A��'~��*��������Q 2ꏶ}�-�N�l-L���#��Ţ�����������A��)1����M��#�ޜ�V��K�zN֌D2��������*��-��6��F>$.�>޲=gH�ScCssZ6�{/�r�o�1��&�1�d������q���	�{�r��X���Y�Q�(�*rZD�	�Ǝm��.%�������~���eOVzF�&hD�"�u�?y�*��Y�5�����]Z�!��.>�v6&�6n�N�����|��.H�1���������o=T&���`�����ae���p-w/�D�|B��Tf���w��$�\���8�=�*��-"���_ΰxnhcll^�*.)~e�����v>�_{3�e��<��u�;��^xy�d��<A΍�	�ֽ7r��v.X�j���C��!'R,\u~���ߧY��i�u��S8�}l��0�����γ��-�K�<H\H?��m��]�u���E�yh{�	�}��b�1^V�VvBi�O�F���|n?\]]���rfJK#Χl���N5�(m�[��F瀷vr�81l�]��@�)?�U<�.�?(�!� �u֩ή���4L��)�Fq|����-�={�%���;.x�g�qqO�{#���-ߛt0KZ�l�)���^��-�D�&�O�/�sMz|����q�4��j��!���]K��ƕ!d��S��$GG�d�0�Ƨ�����J���k�INf��fMԧ&�
��������eu4�'D��BE11�"'��-ih�:��EMͼ�I�|mmϞ��"�%�Vև��S]|�L޿�a����>�p؟Ф*,�N޷n^����H��KZD+8[�.�[XZ�n��	8K�Kցw�N�{T��ng���_�����V�.��5���8��he��:��9�����b�M�l�Κ������DCS���Α��ӌ�����۽9zX���d��D�_������V>ih�->48$�w�*�ljBuG�����̳߼*.f��Uj|�Ɣim�2먫���ۻ��	x=v''�ܳQ�����#�'����*25o�����3MY�E����(v�1k �W�g>;n�iM~�]PX8ۣ���pol)��?՗Ҿ!��\����!,@�;��������QJg{֟��=T��[(��%�X~�fO�l��>�����j���>����kvik�I��6.�<�>px~���b�����M~�lQtx�پ�{q�>�|��>^ϙ&Ά�aR�;��Tw}ę�ߥ��dedP�4�in��̷��6��-��E����!Q��+�',���,�ٿul���xѽQ�E�E�|�k���~5�'DX��dV��5�T񍛅 w|��@��������i�w�����7���TZ�n��޺��b�d�r籴�vg�Pg��%��L�#5N?.̹�{!<?�K���+O���8��/�l;���it�^�ml!(��l:��a}��]]�!�A�����u�]�j���!hr���5H�PWt�?X���"Y�M%I�`3෴�؃kޒ�F�:�֠gj&m��?EN�qG �׽>uSz�W�do-4D�A���>���{v|=��;�&��6���赡x�-s_�i)�Gl(�O���{����B�hb~7YjvwS'FwS�=�^J��ʾ��S�~�����g@�`E��@��Ԝ����fJ�G����䘖3�(���p��5O3�筧'��l~>��,�s5� ]q��X��X������"ZaA���>���(|��#�U�������]ռ$���zw6���j9�_�+�v�ϯBX8�u�O���[%�}nK/{n9>I�>>���񝌰e!�կi�i�������̿	�4�ۑP��dd�����[�`+��&��=���hze7$����[�%O�22��9��2 Pzz�{�������1Z���ab�Ɂ��=���6��B��L�gwce���#�A�������V���u�ʳ���LtBFG"�{��0x2j3��5���9.~��7�/nx���E[Aa߆�(1�7����(1~Q�7����r�чhЭ��tdw��n4e���O���&���0зt黺ʛt�Hr^�G ��E&�I�3�Ή!���W�A�g�u@i�j~� g�7"�Mں��U�߁�g{A��ԨcL�שt���r��Zٜ<��F����{��o�K��鋻�_|j��h��)0�$�t8=3�|ɲ��E��Y�U�������&W�Elp��#�,J��Ʀ��i������8��v&���k�Խr���������	q��6V,g¥eN?٘�Ug����t�� op�(W�T�0KJK�@ ��s�\��s�f^`F�t�W��-����	:�,�f��d{pw���KM ��5�B����rK�Zh®in��D JE��K ���gƻQ�<w9xz����O60���ބ�ʸ7+! k@���f�h݆<%�/>>9���d��1 ��o�cm���ѩ�����o=0SS����U�/��d�?k�z��# 2�2�98TX�ٛ������u�Й�Ҵ���_����{�]|�꒸�#'�\t �Fr�ps
60�[�I�1��r��t4��u���ױd`���p1X��3�rr��`���3���aò���uz=����UZff����M�qv�=f�,�j�i#�������٘����^�f�r����"�����]k 2�U�(46����^������Z��7V�S�	_м�Adsǚ��XVV:R�w���׹�)�(��ݵɵ�l?w?�)��_����"�>|N˅%��{�[Y騕���4v��������J�� !���Z������L�8�3�r*�ظx�8�Q��ƃ�q��})0�H���\
?}�]Sn�(�?2�&�Lz����F�Zg�G˽]e"?��-Ώ۲~B&�r�:[?::�,--�im��i��Z%̯�į������R+��e����vt2ڻ���t��ʁ���7SG�!��{7+aMM����������n�
ʾj�Ct��-x�� ��.0�����:" τA9<�%��郿�qy�a��}h���ɽ&x�u�����i��M���c���I<y����
[c��������ӛ���^#�'8]�Q8�y���0�6��ڇ}�hb���O�g���V�w�E�=\����E{ﮭ�����T���R/�_�&?�,+�+Br��p��� n��>��{W�OԀ�G�~v�ø��eH2//�׿��5Ij��S���M�Y���_�8 �݊�f��[[[�I���I	�Y��Zy�{��VnZ��+��އY������##��H�v�����O�Ճ�����b�Ɗ&�5��FFz����}��=Mmδ���`E{]c�q�9$�����-��_�����ߕ��&��\��-��<,~~N{D�y#>�cx����<s��]��Ci�*>x�݇�-�*fq�q!��h@��)�����d�q�G�|W��J���_��Q�~Y�r�^����?$�o-�Ƭ"�گoܟn��'�ϋ�u��ǫ�~��W�S���ӗ�T&A�ڣ�B��C~�g�(��I
!m9��fs�t�2Ӆl�� �:�Ň/��L��ou3[}8sh�������%@M\� cXEa��Ї���Х&����׋�:׹`���nb��g)��M������E��?9������٥�vK\#j����:��ǂ|�~����=��(+����T����.���ݯQ��V--dd"��de�QPQ����<y���[Pm�׆�M�} �Bey=�c��Мyө�&�'h�i����#<��[����i$�-���:���"{��>���J�iO��H�����Ǭ���|���௭�����"����A���<-G�}B��c�(D$X�п���	%��k�����+�"�2XX)00P	x�m�z�������mu׊���m���E���E�99��u�~\�r_ �T�󐘓	%9�NI�\��NtT�*�[�	��
Mh��6����(��J�O����n�ߗ~�f�$QkNlKh�u��q�$'G�"��&e�w�@�����@[x!^ң ����N����{�lSm��b;��k��xu�H̅��)�ɧF&��Ó|1K[�Lc�H�kx�O�u�k�����s^[e~��P���.m6�͐�.���!��&���b����*��zV�Qc��Xa�����V�#�͝䵮�럓6<<���h<OOO��SWؙ�X��<�v���y
��gH��\#�
1��9��5W_t�Β
,�V��yB,-�Z��I�ј-Q*���hS7=Բ���r�E{!�@�&�U�^�&�ı��n��y<ʚ6M/�x�:jtz��KQN*P:#
��ܞ_B� �ا騩����!ly0�nc(b� ��	?��:H��)e��3���#������շ���˅�����];E��O����\O�ʕ/�$bd�HkM��L~�j��:�a��LT���~6޹�b�����r���9����8O���6��ϼ�y�j%���(i�hh�:�c��ݫ�.�G��fu����$�@9OM�Eq���,H!�P���[s+z(]6���b Q8Xʡ�Lw��8����ь��>T�5d�^�6o�Bq�?C��p: �6O������5m��7�j��<RRQq;84�w�mn�	�ܝ<��@�s�O�p�O,�L'ZC���	�$�.
 ��W���0C�'�+���ӋJ��dB�4�N&���[��:�RQ�d��N��V��o�������o���}.bYؤ�r�%�j��i��D�aD���w�<SDg�(J̠�7�,
e��$1��Y`�@�oE��ǟ��{�����QEw: ;[q1��Vr!T>�a]�y��E�IX�V���=�Vm	!��(Y��>���e�وn�V@u����1&�0���p
��DFE��d}8�J�<�,�cd�1�8lMK�˛��U;R���l�����x6l�k;A����I�������ՉG�}���X8��H1ξ �p|���l���#U�%P�I1R��A���8R�����#��z�pD��M&��`����۽{r�GX���[��V���|S�.A+�w�upС�aL��_�~㜥�������z@��9b�Eے_�}z���"�uv��
��a$?R&R��C�B2op	>MB9@�����KW�+��$Y���
.а��3��J^)I"�"t_`D"����k��N�~k�O9��l��}�0/�ڦF�8�fK��o ;0�0�s�v��� v��)ֻ�b�b�V��r�@�%�M�ȹ�0U�f��@&��Ҙ�;җ�N��̻�G�RS��M�{ch�s�n"(�J.�G�A�҅��������â�Z�ڌ��]�6u���3_ � ��@,*��
���Ê�%گk�w�t��6K_��Q�'9B+�8P�F&(q���d�o��h����m�^�=t�K&`�م�����+�G���nv�ܭ^jwk� v��.F�5��J&��y�"U����g��Q����4�b{�=�&]��/��K�xD�(��n�x>���3g+4O˴Z�ee?:��
�=�s	_�@����3��p� �- H�A����U��\°	$w��/�:�C�Ob{*�Q~\�R�&N���N3���JO����w�|�}�-��������W�Q=9=���H:����_�%�g_R�fZ����Q�����]�8Z�Po�{Ʊ���-�X�*�������~z?+)F���������֮��zl?\�N��a}0��ry\uބ��x8{<�ӥ�`���		8e��e@�m��K�}�F������F�Є���|:�^�����P(�`�KC%��v|\�������T|�S1Ć��-�Ǐ�+Q�������cy5$���{�>���示H���J��h�!�����-%i�TG����4#-*���'.n+s�"���e4�� J  �ē��u]x�z='y:�>X?�X*�@Bt����o����	�Q�ΞdGx�	'���0��`�n�M<33剟G4fY�y�}iA�m8����89.��C�O�>�=��u6}�m�h�^�K��ao̞waa�Z���7��Xc���`Z�ae�'-�mB\�$���VB�/d
�5���B�����EN71� �$r���ϟr���F��3�dǈq�����GW١$$�Y�(U-�c���?"ΐ�>�5@�,����H15�����L�靡�����8P+b�*��D��V% �i��I۔B��,�t/p����D'�@ۀ�Xf��|D`��@u�U��@�U���[b9���=aB�9��O����v؍a�j,>��G�����<�l�؈^X�X�4����A���b֓LU�:/+�W���II����m�d����ѧ�z�@˦���Y]qT���|�,�6$����������Q�n����x);JqI�	���E��~\ǂ�<R)9�Ήz�DK�q��ʠ6��Ci��|+�F]m�˧og���G!7�s�-ee�.	�ʴ�&�ZE2DQuLu�!К���:N�cNaO�o����x}��?7E���.Ѷ8_��{l�}�G)��^Ha[E�u"FDp�;��L�@v�)���� "4�˻#���~��T�����D}\\u�X�G�l�cFM�y]g�Cfަ��)�s�J��m�j�hBR�3i�wi�Uc�xɵߺ-���@)�󹤃����{Ζ���vf��
����辷���إƱ��\N]�̮ �����D��J�n��3��ښ��I"6땲����Y8 ]�����!8��ekW=�S��`����d�X�ymC�۳'T��	�ϱ%;{�D�Ʝ���V&����x��o�<N+�\d�\��N����E�՟p%!feq]�L?|�p���`ܝf�}d^ه)u6*T]��^�Z�L@􁚚��Ƕ񅖈`�NFT�(\���D0:�G��Y��ĨIƄ�vU�	y���-��o�+��6�� Pߪ��ߠ�]�'6�-�)F�_������CPs׍m��G���u~����?Y�T�Iq��ho���`�8^�5Wn*v�������� Fnǃ-b��@���$R� �`���ff���6I�IXXض�v"Ć<ȩ�3�<(tD��r9i(���%�����,�����TdJD��ښ�-��T�GO���I�����Z�W Y C���C�����b5L�y��
xLM��u͉c$�調@���M�N�Q����D�䐃k���o��]�GX�}dR@$BpPs�
6��ڀ�"O�>�}�R�9������3tj:�Gf�/	��ТK�[�.�F�ܳޗ�Ć�0h��u��J�J���x�D��qqq�ؽ�$��uurڮlM�q0������W��L44/'��WyO����V�eYM��T	��?�=A�Pp�w0�uO���؍�BP��R�['�����2�rW3_|�&-D��?��f(��M-df��5��I�L�4�L�*��+p�+��ϩZOM�Q��� 05�=�w��a}V�g��}U�-��a��[�ۨ?�i�����U"�ͧ����w�r�|B�˭`��Ҵ�̟sb�BB����34�� �X�m=���:�Í�2�.|�[tB�����!.I.�}"���%H��C�z�νOw�D��,V21��7��3M�V�;8G�C\�1�CZqa�i��+ၞ ڍ�y
�����J��"���R9�.�r�������	�����������Hh�"��E��DVV�>�Xv�x��&{G��=V�����Ǒ�Ǳ�,�4P�^m����d����F �E��с�� �|/���C)��W��������硡�JJ�:����MSiQ��8�~n>�eӉʚ�Vː��#�е�#�㒈˴�ΐy`I����hh�����,�H�Z����r���\�S\�� ��L�� ��e�P�����>o�\P����2�}Oa'�-���ү��N�7����&a5B �3�w2Bl�Q�f%f-�?Gy�~sZ�Sq�]D]a����Z��|�j��������"��ع��磈������������Z�5l�>ӗ��燠kq�����F��לh��W���U�OL�(7P���@�k�"�",J��U�sE��u8oX�:_�qp
<��T��6�NN��K�T<9�����!�kLu��<��.���_�U(s��vŅ4�	��Χʀt917��MO[�q�5ddl��D�We�RC3v�E�H��� +��G�C(y;��d\�Că����>p�7!��؀�rt3`&;
�n��l�����	R��)�2���\]1��M�X�g�����)���a��<���}���-\e�[�U�9���tT5��:k\��҃�����8[�8��[�� ��&k��3ցHWAa�_�{VUI�8������M����۶}؄��8://�������j�3�w�nh?Otd����B1bf��7<u^��TRn;�����,f7�h_EsgH�"c�Rh�F���5��F�$.�%I�|P��$'U��CQ��q݁l�(��j�g�V�*2���X��6?xMH#����{���#}|�V�����!�ZY~��8�Aa��ԭ�]K&�`D��E>�N�F�Q�_ʴ�E:»X�BX�钭Z�o�SNW�qȱB]hϹ��{�N�~�����~�,A��c�+_��h��|hU�Va�c��p�(��%%�������	]�e��Ğ��ǔw1���≮ɮ�$lw~����>��)�Ƒ��~Sѩ�3�w5�#?��`��^�ku�q���2�};+��"Ac������7��q���C�o�и{9�DA����\X�夭śV�W�wԁQ�:��	`B�hq��7�v��#����$T�1�U�K)]��䉤__�@������A��I㥖n��J���	8�f���qҴk���ns�G�ץ! 1ȇ�^a<�
���0��O
��V?�;�7�~L�2}�wj�B0�Nv�8f�R�0.�5�ͤ��|-a��B�n�}+窬�1��V�*��\"�sc��0�u5���H�fQ�P��m+��5/�b�r��c���i`��e;T���x[��=��rpO,6�Y2ɀa�����^4X����kYd�^l�:^;�y۹m�Ƭ�҈Z2(���ߔ�� �;w�B�Q���fϷU����a"�3�5f|�vg4��D�A��i�q:�~����	ǋ�ڮ�3[�2�
.(D�3�*,,D����ղ��b�2�2���.�C�r�w�B��w�8����t5��h�f�e�v5<���+!1�
f�Q��r�gX�_K���I�V���������b�`�#�T��8��"�6�wB%�!8P�Z��)ֿ���̺�f�|T�.�_�2��8�����!�(�C�Z��}�4�`}�<YW�q;�-!�N��:d�*<�/�� �NF��5����ã�P��$nhw_i��g���ׁ�� ���g�of�q�x�Lڠ�1+�D͵�]zh�x!*�%��ǳ����:��|��ݷ ���:>*��8�M�?ky�d�z>��:8�k+��"nz�1��B�\C�tmd>MM�Y�	%JA��ZIڴIpM����BY�K]��X�����J��ݜ,~� ���xJҊ�loo7�q�s��5�ԨTd��:���Ԅ��X��k$�4QlDPB�c�[r�8T'Q�U�re�2ߦ%�AT��%a�^�H����-=W�E��<���o9�5������ �Ū��u����4S���~���IA�N:���۩��_؅�����*�%�6a1���sDod��cbE�������e�1�M�};W��Pu�9YرXi���܌�l�Q)�)��M����%&~p��e��|�A�a|ڹr�3��<%����}D�ui�u��l�_�Uc�p�q8���92�r��,�S~�n��l������� +��~W��Ta���B��4���Ԟ
\>u%+%5�#��.�k�pHL�EA�#I��S	�v]YY���;�j����}���1�Ƽ ��j��J`a����,���sp� *��}a��� �.�+yP}K(A�_�Z�(z!&d�B#h��������^l�c�Y7�o梏�2KQ��&��ɚ�Qpl�A��z~�I��ҏ��|N���+���ņ?B��s1�S�������&!%����MgԨmV��%���C�(k�1�X\�_�3'�����J��],΋�bT�Ā=��Id�{�a�,}x�o8��kg���y4*�^��/mu~��s�h:�<�y�X[�W辸%x��q� {դ�E��5k��i+����A��ݴ��
^:��g7��S����&�<��R�IHAv�>K���ZgWHN�T��aEئ��G!n���3��}h)�>>*^M��"�tcJ�o��]a�n!-B�/�ܚ�*B�������RY_Q<�ؐ�=*���
8 *edB�ӒL�A�C!�<7������+��mf�Q�ۢ\b�G�&<ڵG�)H�ݷ���_��S��@tf��q�_����IҮ�-,.	td9������)�& ��Ba�$zB����]\�C�'>f->{ӕ�&&��ܫ5�q!��@���cmU���p�������[3�L�mW����SRT�����c��q��㬛��}�2�9�MN�
�@�=F�/����(����r��B�8T'j <���8�P���޲�� VQ�IY��TH��8}�#���#By{h���#M����v��2��A��Ǒ������~Ɋ^���T��Gÿ�6m��	���{̶�30<����LJ��$"m��8(̚1�o�sT-z �'���Čhr��9eH��~N��@�R|v���a�E8�-�d��E/���}Ȧ�m;����@��
�4U��ܬ:{L�͆�B-qA3�O�A�m��q��3�ل\��7�k�o�V��G+$C������L�Z�������h��Rʘ��ѫ�~���� W0�t2��P��bj`�$k�m�X01Ys��x��6_x�2���?�}Y3^��-��-)�je+�u�K��h�� O�hl�E�\���R�W�/������f
�I�y|���
�.�3h,ȣ=�ʗD]�������^�6ŕ*��&�K���Kd�'��I�t�!M��քH�����F�E([S�۱����jy�2<�Ie�ؖ��i��Y�A�����U��~��F��	�$oN�%�/G�O�^0�Io�%�G��adR���Iic��4ԮuS+-3ᐽ?irA)#NG���N*|^w�5����D�M|��ޡu堣=��v-m09`�R�Ŧ+0�*X�y�.�4=�\�I�US\\LC�tS=��Tr'���ey������i2g������"3}��8.�D?�!�?���C�F"��m��@R�TE�TVJt�#��E� |dU���"�'�����J�3�5��d��0�2�T���X�d�s1p���DbD�1FY<:�z�IU%�DK�>U��4��j}:�`��J�Z��g��r�HY�9��������/�~8!� ��Qo�?Kq����l�����E�q'g��!��=���&}I�4��P��h;����I����vC+2��fV)��1z�3�> CN�$	fͅ�O,��5�Q���cOm�j�����2��%6���Mn�o�#W�+�֓�0*o��d��q���؊I&/?�%�(#g�\cq~�~8g۝��L(G�; 1j�����Z�=�"N�����|\�
�Ak�����G����:A��K�ko~�e& b$��x���d�ѹ8X\|���l���)�.} �ՇR4L���ab,�ՈW�����~Ukz\o]vmYP����������}:�?B%v��'3��Lw�m��_��4�F�e���I��Ӑ�FM�yl�M�+t.���ߛ7��m��ʏ�;\UCϔ�>pˬ�Wmv<W���Y:_OIkg)c �~��]��	�����g�`�ɯ������4���2�:��j>�va�M]���A��jȾ�4�l�oL &��@�f/�=��,�tp7z?j��x�(��$`98;OOK���&a�a�����/ǝ�c ���{yn�v�dt�V��G=W���ݑ̛ P�&1~�Q0�Q_l�䐔5�E�*�D�|�L�P��Dj� J��ɯ��Hi�ak����iD�TwI����q�!@�O�X� ��+T� =y#�K�9����](�0�|���aB��&�X:b���;��Eڷ�y�*z�2G��6B�tZ���U:F��P�A����hA�hA��8����c��e,�H2m�c���ބT�>�A�`T4a)�L��"D���ŵ
�eH�Cg�)����ց|ْ�^}uJ�#AT^\r�IG9�h�aiU=tԴ�Vs�VK���S����۪����l���(�ɽl�������0��{�pO#��Z<.�>t��^�v؞���K,��o�5�����,�S�P�Ů'������,�������Ia	#4!l�k&yl������:?V�:�u����4 c�'��E�?��v
*�wNќĽ����&�P|��>]�����E9���m��9ۢ%3*�N�����.��hvb�]|4�8[A�	n�U�b���W��.ؓR����X����=��̐��F(��.�%�`��/��b0\����e����7�Qa�wd>�$��0i�}g_�*l��UK+�2睫������ƫ%�;F�=����H����:��6JC���7N�ǥ�������Wk��W)L4��vK~���i*���:�i>6�8:=]	O�,�F�[� f��w���l!��p@�J���* �;�L��8�H5���HQ����uyf�	e0�vT��>����>/5*�d��HF+��E����|�bf�@U1@����b��b��n������D�vd��&���''�2PC'�*���Ő
*����_�w�{4$��q��lp���w���cIU5��p+�sJu�*�Aό�-v�G�����Лɛڰ��[Ԧ�]���jb��=�p-�	U�?%u����ǃb�*�{�Ou�m|^┴54���:��Χ�����F�m���nU��]�kZ�ʨ٨:<����KN�\Ap���ZZ�O���P?�C���0�/t�I���6�q���Cl
8F*>,�ҭ��8 ��8��?��B3�h�h�fի}mC�6/h�*���A�4�Gh��Ô4.3�p�����ќua>&fJ�J�}m��]{X�7(
R�p������XTE(@��Iord|�o�=M���n�.�1FZ �El��M��&#����H�:�å�	�Ҷ�8�r�r�3�J��-��3�A�ߤ��}���r?�z�~�ݍPSL �_/�kY?4 �x��E�� @�'�2Qk�`wwO&x
5<6| 7+�q[��pg�W���W�0j�ֶ��}L��gO��`Ss�G�l������5-��Ԍ�K��9�[7T�)�s�e�`յ�:�+jz�.55 ߋ���<�HYPJc���R C kI��$2�3��9�Y��Q����ۊ���� �r���+��E��D�2��$0�3*�"@O	�%5j-Kt�ڹ�0'�i���c�/���1nA֠���K�[ LK��}3@͢���Li+���v3��/�����܄D���o~����@@��
H�h��+,xd%X����>�� �lI#a����$!̂g��NN0�_���A��:��U���U���s�U�����_����`S�֙�k�O�}��y���@f�1����O�*9�=��^f�?���-b��c{�>�=Ͻ��x��Pjy��l�n���ܞ��/<}������s���%��V���x�S���	��},������[��(|P��N:c�F�C��.�	�%ǉ���++��5�M ct���%��EDd�5k%���kHo$���^�	�@_�~����G%]mIqt�����6�n���x������QvH��=I&��}fk��T9��r�A���&B�O�����b,Og������1a=]#v�9lCp'���@F�ROM�|A�d��
)P��H=.��8,]d��`�|d�ʝ�5Z��y(��1��E	�n�N���}�����M���Dy���bԭ���/���˸*J+j��o�s߃��?�\��/T���ҲSvL��~�s��]��u��;��;Z[�5v�\�o�����i9�ek���'�S�ǎzc��  "�X���l���dR�� y��,m��2�!��$@�AQ�X�J�ׂl�"7h� ��=��|�N�@R�L�%:r����%�o�eg�3�İ��39�_ Q�D�Z�,{�ڮe�	��- T	ʖ�f/�n���	�T�#Q��sx�ܜm�ӿ3�V�찊�H6@��j�K]N�ǝ�ͤ��`pg�}:}�K�K��Q�$J$L���v'�>���O���O� ���q�({�罬l� G�g�]K
:����
�a����"iK�=q�0�=�6@lg��b@����������{88,����p94�՝Lx�oh�c����h����]�X���w������{5~����9f�+���KJ���JC��^vv�7��*=��0��AԗD���z,u$�)r�'AQDX(#
���{��"f���'�<��;��+ �l��H�(����Ok�=�S#h˞�o����rE@��p
�H�5w��L�K
� �~vD�6���RWF����zF��"gtn�_,N�I�j��I�ö�|HV�Q;�5����<[�_��/�8J�"UΟt����>Q��$/D�Q�f!�#}�p���2+�l�&~���� ���
'cW��c���P7�����ܱO>��r_��|}n�����Aȃc LǹX��`6CF{�������{�D�&�p�'��z���x�J�� �>YY�3L�t���Y�q��b�iKo�ױ7�#W�WЇ��}��eb��u�޼yC�=��/�~�Xg_߇&�f6���-, ���mp����͇����n�r�� �j�K�T,����lIQ�73:�����1odh�K�{�Ш���g�H��+�XN:��R�LY���gT`]�N���q��;��v'�2$����I�W����E��	�&e/�)�x��#zZI2�S���%@���H��D4J���$��������w�����U�I��E�6����5�b����õ$�'�5��S3�0�af5�Fg#d���(^ڈd7:'���	ؔ���5a�{D� v�&#lS�Ł�l 6��md�s�"FU���a⡗���z=ǩʱ� ә`4�Y��� �_������w����2;��Ţ��	���?;Pe(M��FRpo������J���	�3���c9p�
�y(�"���+y2�}����4O�-��/�K'�kgN&.���d|�����.�r&�&0�p
����N��z���+�\n;�h���--��^�t����p����LYY�u3����}��������n��Ց��;�{��R2r��|H�-$}����+��ǿr����n�\��=�梾}��U�q�˨�ү��%^�(eCe�n�����0@�-�V�G�tHƲ]���LA�JB]W�V9c~7�� -�
��b@Y_T���^a��Е�LsU��m���Փ 5�.ur�:N(։f���kM�$@�Q�FꚊ�C���J�1�ۤ�N����#���ߖ	t�
�LQ�g�z���:M�[
=x	B��,�q�z��,�O�؎i۔4G�X�䣾¿�G�(~���h���T��n� /��p>(�C5@���bGW�f�S��N����ߓ�%���L�����S�����'��c13���4��ŋ�:�.~���n�v�~
��lea,o��'���V����8' ?S��R}��!8NA�w�>�FQ	Q��%|��;AJN* ŋ;���s�(����4��Q\����\��ǎ��I��V�mq"'��k_M<�*��������:y��џ��|>�{�S�����"ړ�����I�عm'�������;�z�zbh|��L�"�R�͍��HͿ������6ZW��w5O�r����d!���h����@���S���H����Q/��+
^�F���������!d.F�v�� 8~���ۖ)��0az^A�.^99��=
�C>L{�-s~2��Z��	b� 9��e{�V��LS�A L��t\`*� k�2k\��J��/�SZ�p��`�_"�"��?N@c4-�NCct��)$����F��
�UI�#b����a.ҀV)3����Ѭ4A��#� <֞s�TxJ~r����#��[a���8���O�>�p�u�Î���z���)@�W�S:�^
ѐ7����Tiy�� `���t>�҅���֯��U�&&F�w:2$(1�NOMU;vx�x�������p}g����� <_��%��#@t6s�y�-�S�R�^U���,ĥ�BKF��i���|2��g� ��O^��<���)����$ |���#� s ?���g�x<XNk�"��
���po���K7������ݳ�kӅEm�9�gsrr������a(�9����C;N�i�����;�S2
S��N�)�|X�¡��ʼ��w���[���ʾ����#G��4�����RQ���ӓ^2�dz���l�"�ch�	NB�WZR���ze��^
 <��~�W\K޾�ςQ= Z������̈�����5��$3�I!�i#q4��رc؏1 R�Xږ�'k�5F�������7����M�������57�66mo%`�0E�DZߒ�tD����=�ެ�ϵ!�zNN5֙�C���͟��1��-e�I��[�v�
h}�N� �Q����D,��(1M"��?'���!unWX���жA��%ˀ0��s��8^������A.�rPg"�9�2��s4���>�3 B1��c`  �������5����؛�9 w2�2�G�rq�ԁ��y&2��a�
6-�Ӕ ΄�S	���5.Y��ՋR�����'�8�hM4W�^�����,�&�S��!�{����Qq����
�2�2�
��:��{QZiJ	��G��yzH��g䚆�7��+�˯�[�������z�zoD�O���X9�����ɢ��s�֎�"+**n/((ԑT+������|���������|��pF�?�Y�41"�[��ݾ��/n�Qr�6;gb�����ɉ���{��s�?����8�h�@=6	�Wa��G����6����F�yEE���_��{%�3=�q��{z{����9{F ���\wF���E�Q �;�ܱ����)��N��öN]ji�P��5)I	33 0'��������a_'b-m-�~���d1�h$�{�؉�-��[x���H�.����͛���'`rV�D��j����N}t�H�l�L}���U?��~굋2���-�@u��5i�� ��t2��ROQ�� CC���O�t9e������,GP�vh�L8nR�'	�$@8"!�:K)����L1$��u��A���\���C�9���02	߬oh����ݯ�B]�����ONd���"����M���p�I������F���&6#�%M.�+�S�D�U��Jt��'�G��GDgIֆ�N���	���K�^�5Ӥ�
�(fĎ��Z� �cT�^���I�5Ӈ����x$/?����Q�t��a���K�ill�?22�a([�/4~<� .��ܼ�***G��RWװ"[R��?��ȣO�<r����������3s$M��,=_U���75|��-���oe����#�C� ���n7��  �A,�Q���yortT�oE� �2/i�zD�Y�8�X�h�:q����SO�����Ԋm��i�=Y"���%���Q)S�칦����;'i�'NȿU@�5b֏�D$zV �A�h8�����6�I]Ѷ���5�`ndb�\*�HS��k/t;0�>Id��ה���N'����uq��[�z*����Q�ֹ��,��vF��7u��E��0���>}���9anF�bI������7��:[���<��)X�*���rBZ�fMR��'�Aec�D�(]��2����v:d`R�>�eٻ���h���}�1}����֭۸b"utxd���挏����� ���F�)�q]��<��D��@rI���M��������&LD�T���e I�V��:��k�E�IV��E@�K�&2\�D@��
-c��#sp��3U�-�)���;L}M,����}�.�����ٕ��w��Lڅ��5X�����jj:W���r3�x�X*��s`�)Y��Y�Y'jkk�UVԬ8���z������T[_�'��ܭ! L8=[Ҍ�!o�$;���?�skÉ�����p�V�[[Z/�?���;8��_�ǜ��T+#i���j�r�XD��A������8e |ˑv/**��񳴪֋"�cT��w�}�I}���N�mB���.�[1���(D��a(b�t�	0gϞ��5P��T��t�>m$��<�3�#�\gWW�,�����B�G.�4S,�M q�mT��,�/Y�e�3QS�:�ͤ4����IU\A�7�%F��c��f��7� J;a����HdS"�e�' �D�6/�D�L�k�8K!l`ǹAwZ��qa�k��E��/�w��X��;����t�8q��� �
N��h5t�OF�(ى�Gd�}�!8��rǬ
�^�(�|������s9�,SJ�0?s��OL�݆kk'��Z8Z�&�.@�4Ε�A�\����פ5R����!�s�-����.� Kd���H�F��f�� ��i�R"�f[��;�D�Q���,�0�"�dyL怵u:a&c$e9��("Hu�DM��iõ�;;;����¦����v������K�OljbLd*ؒ�}�}�5_l~n��6m�g��m+.�E}6끧������::5�����p8=��
gy�X\�BI�ꪊ�q[�wvn�j��'�����`_`���wc��ߢ]��Jd��$,�#��ƚ,{�29��z��F����Kō����{�E^e�:/#;�8 ��{��%U���`��"�蔀M�q�`���D����T:8,n�聿pᢤq��m�V���P������u���]
���5(��D�7�LE*��-�*U��6�ھ�����+�+�|)	I���?�mh���W�Ի�LG�>�7�.�!�#���� �)Uh�izF�n.ζ�.���BE~E�Lt�"�o�9IKX�(��"ö5)ÚUF�QLx���</̦Й
%�E�Z�F�ҲgJ,'��)�>����A�� �W�������ښڿZ�i�X7FG�Bcc�9(?�C���w���kp�Kq�J\B,c=Zġ\�P�A:n?^����VJ�{ ��	;(H��!	�!2%~��l�H�o�mZz���-In��@m����#�����]H��h�^�����/��Vj��!��}�).�K8��fge}�������¥��¾, �����{��s������ĳ������PIIي�ֿy�35�<��7�{�~2.�

��xYX�RS�Ѽ������m77,��^q��j���k9���Ɂ"�E
utI�K�MC�d���h-����w��!/>3饧$�N^��Vz9�^u��<��#�白޳���

�¢B#�
�I�S� �!�c�-�IQ:j�L�JmP[�.\h�S�'hp�a���
���;n��[��e-���M����g�����Ow"��j�r|U&b�6 ״?�������Ӳ��Դ4J7{K����k�Z�Ykב��b�C�h�� f��`K�F��?��֨����K��)qM��[�5Lx�S�"`Q����oP0I��ܳm�5�Y z̤�^'����iKTN��d4��wD�8/ap!x<���l��d�s�6�p쾽f͚�\�q��6J�oxh8%�r8~����	�l-�\	N^.R�D���t43.����*A4��__��,�a#�@ƃ�N=�{о�:������׍l�ו�y�r���'�@zW+�*'�~� x�cA�@mw�5��d^�ƥ���ЕI���ܒ�a2G��\�H�n��vII�7�m�t��`ڪ��Ui[{����gO��-��k�}}����ᦦ���]�<Si�v�?��oo9p���?����c�Z~1��->��FBQjfzhڗv��������nn{�Ɔ��S��ә�g�����}'�Ce��iCR�l.^J�Б8�E)3+�+)��:Zϣ�9�!����%a����J�1,ꕕU`��U3M/2��Q��g�§����gZ�Dl��Y��AS"Z�,?W"�<�{��t�7m���:d�|��}��y���;��Rk�ŋn�F�ߎ��V,d �zY$#��u�+]##F�"�cꕲ�.�Rɫ�Ql][�;�#�c����yl�����$b��Ř�&.z���vn���!��Z�6W'�3Aq��L��ѫJz[�I����uyS_��@Q�\|̋�a���	N	��$�I�G�_H�r� 0���Ӎr��!ȱ��a�8�����i�ܙSP�&���ёd���=r�.����:w!Hd�S�ZΝ���R ���O:~�����e.��Q^A6S�^�l듬m�R#������c�B�7�x�74��Y"�]X���wn����:܆��u�x���i:$,O�F�t�m�N@���@�Bv-���[#�:v4���.��ck<>[���~�����rUu�3e啮��
Ҳ�З�go_g��s����H��8|���zoEE�ث��r}�k�޵~ד��������Yk�RmpH�Ps2�=�ũ��yC�?߶c���z��_��=sӱ�G�@�."#2/|V"8F��n@�|T�v�=��t�(�͒���Gy��è��x��y^yu5R��^]�F���uvxO=���	x��e{E�P�)vI��q���[�S~?#q�ƺF���'q#���=3,|� ���{��������V��
O�:U���y���Ȼ��g�`���"�a[�D>vI��F�Z/VH8\�-қ��=/�h�(�Ѿ��O�y`�ƍ�%�bU�3�u��i?M]�����)N�l�%�t��6�L�f*�����0r��s��DWO���Y��+ jv���0F�-j�i���Fn�zg9@R�,�$�t�%uu�ޥ�]@@k�T���!�����_]�v��lڼ���������韇h���[p�߉�yB�r��)"ݜ/uh�$B�A�%$_R��p�&ц,Q���S�����zy�����aKKVdiD�; �8mfT-I��h���%c�,�ɇ=��3���e[���:���;�]^W���A��>��|��w�~,b�s Lk�vUخ�pH�4�&�d�F�L@�[�:;Zqm<�{��յ�s������<]��Y��N�v�:u���J���^[�n���4lh[igg߱3�?xh�m�O�������|��0��C�a,R�^I~�ٍY�k����sFW��uu���~���������D��h��rޖ%�%��3M�E�Q���l/~Aǅ&��a1���xYY���[��Vy啕�0HXGN�{�	Y���ʕ�Lf7�qL��'��%O���� 茆UI��[݄��m~�'/7�>��O<z%�Ů�������-h��),�[� c�B��;B.�1e@~�z򆛴�Y�$AMa�p���l��Huud	�\p.9�K6�#e���Y��9����m{3�x.�|��* ���;��|竧�W��ph��Y����-�X�~a���I�+��e!:���sKG��vq���&�<A]3�!8-_\�~�7o����՞���/ԁˑ�k.���)������Čok��7�?P:48t��6\�k`�
|_���H�2�f���@�J�T���$�I{_��Y�(Η�K�	AS�e ����a9p��c �*��̶�9R%@�j�̏S�I�,e̮�,qm&H�	���N�bM]�K��	漇�<��QA����$?:��A�ޑx�뇎��+*�˿�m�w��9�kZ�W�ᅹ�	d�-�/��h���x=�+��p+й�#c�����By��0��0�D�۹�W��r;_�Σ5O�9���>�W�9��iY^vF�|}u�=o�q�7v��,b���f�sOm;r��בJ�j�޼�E�<����|Yx(LB���'��4��ӽ�Ĩw��oth@���ؾVQ�e�xE��B�j�l�|�QD~=^z���rQ�[�5_�5�2�e,�X����JdX��d�����թ�f >�,̍h����?��k��}߿���g�������;c��͈��m:����?;aMA]���y��R���a}XF���#�@0�b�:_cߛ�2L[Po]":�����X͒h�pBEδ���~�X�Z=��)���joF�P��S��S��>'��P���F�[k��ʷ�j�PGM�(� )�uiq��I���4<��~XQQ����p�S�?
���b��>v��7���>��]_Wvooo����L�{J�PD��gr倔\f�p�����l��p��zV:�Q t��D����
F)��dA�ɍr|8&���ĚHW#u%�`U�WIvm+�3[`]K_�g�j��O��|�~���ן�����%�ю��	���IB���T�g����	��=��t�i�0K'.)x�UH�T �Y��_��������YQ�no���7��w|ztt�֙Ht����[�ly-+N��Ƀǳ�o��/v}2��ş����5?+i��(塷l���l�>��H����Myz�ӟnkm��h4�:�D�2Ǜ�[�JKJQo�t(R��J�0��*��B\Ow���xFze� ����*�4����1�4��?z��ݘ��ߋ=�k�堐�����.%�q
`���b��Lo��e�'>�]�~�/����\52�3{v��;Z��tv���n��T�bѠ8��2����t�X��.z�bUa�xɃ@�蟎��z��p����FH�@H�md޹)?�����T)L��OR��t���ʲ����2`���
0������nY�-8X>]R��m͎V����!�JxVU�@`SD�edlTj6��_'&f�%1�M�?�=:��C{`��C�~�����w^Xj��~���kc�����f7�Y�ž��N�빑�����p4S��>���($K��sE�t6��h�9��&�~fO����wCH3�Y�8���p- N����+�9�)��nl��$�#bX��9�k_V�ő�*k[��n�a��s��d��	䋨~gЙ�CZ�L��#�Y��B`׹��B@Ot2$J?��n�~-��v��7� ��V�eI��QZ�f���������r{k[�ϡ6��`�n8��;k֬k]N��q��Nh�7vt}����~��S�795�Ήٱ��l��\D�??9}��oh�s��c�4�f-k�9 b>n�w�3mˌ�����I�1� Sl�Q�E��Z;���J� -~ č�C0��l��r_��>=�����T��mR b[�8�H�0��YЁ+�ra����4�@�5eFSR'$鋋bR�Xؤ�\���︓�g&��[�|���cG��/\�8��߉�XPHS6�lW�N&�1���g�9ї�'^��o~��Gܒ�&��r�~�`Qe}�Ѡ��a��h��V9Ni3\�D*���BLɂ�"$��<w�ǨZR�����i�	#ekB�
~$rᜉ�/�~D?�2��`��&�����D'��x�5��ܹ�p&�(���#`@�T��Cu�s���~��O�܉�ھ}{���x)�5Ǐ� &��%�Z8K���� (Zk�RKH" �׹t��������b(���g��s��P.��(]�?�KV�Wy��t�_( *��bۣ�1��/RN��5b��6+�$������moR�z�ض���E"��M����{K�/�u��5���E��bP�df!��i�8��({��yKA@\ ��,$Is�=� �%��IB���R�>����'O���-�W����x�˫G���Ç^8z��/�9s�N0 b�#�6n|���j�BYWQF�������?��س�M�c�+�Q��cQJ�}v����;u����k�{_�b/�W��-�¹N����SM�߹�3����0�Q`�ep	� o�WӰ��W⽓��H� ��A0���[��n��==�G�) �9�ʱ�Hʒ��9,
 � @���vǗ�1�����2�KR�*�1�dTD��*Up,��x������T-���|�o�
��g?�)^ۣ���w�8�u�	%�|�يH3C���V���+>�>���M�.vYXY{�zQ��".p�f8���g��'��	t!������(A,��XD%�;��v7����q��D�p�d�
��ט�et̴x�t�*����n�9@(S�6������ՑsC�>��G0��J��=fY[e��aϓ�E���f ����NB ҵ���b����P$���'���d����>��Nݍ����y̺aC����2wжa/p^f�.����0�T�m�q�(���N��� �c�r��6`�� x8��B�3�-6ལ܉*�I��J����T�P8�X,�x/���� �W�m��¦�'�M���k�X��:�6�O�'���y5h�PgG	�q �H;�I�*�<U���)���{���d��>��z1x����n޶�q�V�o��ί, ZO�p������e�
��֍�6~�����=^1�}�N������?����q_�M�`.t�sA��2��j���q{���֕�)JO�*��z�599��g��O�?��9�7 vV9�pa�b�f��^z5"lF,\�Yoe$�	gd����G���b�7�oa������G�e��; ��/.��F�z��0�/�[�PJ-�F��ʔ`�3U��0-K�%5��FX�?��EcsQ �sp*N��X��q6�, &�%�l�(jycH�S�0��FPG�A���D�F������N` �k�&�{���^�>w�컰_��~#������)��������6ϥ�xiE��g��`tN"i��t:CR?��w�T��H���*�]�5EoHY���I��E �^92.�����2�7I�:��!U�P�������vl�rV('�fT�FIa<��  �A�IyҚǆ ���}NKܴq�,�S�X[!�Kb�Q#P:�A��;�N&=�r
n��� ӏ�=ך	�l[���<�0��u1$>K��Iuj�����=d�ׂ�·ـI�'�l�X�/��ۿ+�/~^���<^�B�'���s<_��R��%u���ҷǦ��c� �S�'���Y �Q"hd;-(>�6�cP39x����+*�x��/Zu���"#����:V^��ѱ�g;;:n����U� ��ld�ޱ���Y��#+�t�vۖ�S�m����{��;x�w&'��5�K�FR�f�_����G��R���ڢ�+�F���,Hފ���Ň���Yk�u.	�T���Q.nqL`��8>!�`d'"���o��D��C���HB$�t1@��mۼ]�,k��9��!�&�ٍȑ?� ���a�M�ӑPU�P���v!���s����wtuuݎ
+�(���}��9���E+`����b-���4���{��H�gt �;���/����u������5��Q��C?�a:p�w۞}��=mm���< �$�d���1.֤~-I-�����aI�����2UX�>��&-��IX�l�S�N�z��s���6�Y��S�7��j	���P�N, ͖3:	�I��4ȉb�(�U�2e��2,������5�
jB&�O���Y͖'I�(O*S��az���y� q��e��P,&!����Ms��<n��D�"�Kp'�墬\O5L[�1��K(0�'����w�� �5� m ��N��� ������:�VS�2� �ε��6�>XO�u }���6s����P�m���p)w-)oɼ �o{�-�D�B|�eB ��s��H�W�$�m�"'/��"0D�m��i�~���:;gO�<�'��l�j��7c����\�n2;+�u�ZZ�����(ش�F꡶������_���"�W;9��x?���<������]C��LUL�3<���#yw�D/�������jr��hƏ�� ���m�b�m1�t� �l���K�k&"u�����Ij��0T���?���<7����L�A�'y �&�Fѧ��5����.�y'O�2u5�+���.0�Ɲ�t ද�)PFkq���(�Qڲ��/�))�cqĔ�����r�!
�p��Q�5�'I�����V��X� v����ٱ��ܳ e����������U������i^���ׯ����=�X[{��� \+Ѷ�#+��%��D��0�fS��H0��OI�� 3��)��HP&����'h�&�1�(iN5�i[�d�3u.$9���wZ���x<�X��\h�I��~���\�Ц���!�(��0�c,���Ǒ�T;�����$DͶÁ�c��",l�K!�)s�
��q@��.N�M�K*[#�Y89�1�Qz�� �vV��f][�ߧB-
T�ii��/ɏʕ'H�]�cuQ�4�/��@n�4�����ˆ�ׂ��17��p��1q*L�FK t:�Ķ%w��f�KV��G�ݰ�N��j��S���=���{H[$��8z|<gY�DFNe�#�=#ȳ�R��+d,$�ÛC9d�4\0l�h��>s�3�6nyM�?n�[��n ���������ۭ-m���Z�lm�شcǎ/���E;��@�ߗ��SW۾�'>�݇�h<}���`u� a�8��~~f�Pb�}�؅��u{��>g7[&@:��
�`�E�Lb�6)f
�� Ę�L� U�����P�"�O/������i���3N&|$#��(������r�u6q�Z��\	&XP��a5ι�0M
�3�J�IT,.��re�@���I-�� ��rt��H�,c��d�&�x6�y���X�[��Lgg�(��L��ܜ�C_�ڗ��WV4�T�t4ԯ{���q
�<��/�S���/�����ca�ǘ)�I�`��`����+�a�s��pW/m�ph��0%Zg4:6<S�-y�dTj�ܐ('�:D� 8�NfCݓ�W*�a�f�H��L�#��1�O���v�m�D����1�+5b ��`�I
W2*�v�������sҖ'%??_�#�4���#�?d��82ԏ��<.fxl�V�|� �Ds� ��D��cfp�?c���\�� 6�]��$�Y�Wl&Bq�(IQ>�L�V(7cy��4����Ly�1�%��v)/�.5�f�c�o2�G��D�暰�Ь���AL&�v�n:ɈZ�a˚fhԉѧ��Xr�Ҷ9�=��$�':IO�����o�c�T����2�S�̐D���_P6��_8�d�}������������������%>��s����O������q�C��Rii�����f����(NRS3��L��;�?|d�M/>�{�3�wͧd��P3�F�mI~�lY^��7U|nˆ����o����y��Ç�2K9��ɂ����pD�7�z=l����yQq�WUU-)K��*Qi�=ӲX@�F'�ދ@h�b�Mzٳ��
���BI�:����#��>&��,�P��nذ��im�ı�%��� h�sښ0�U����>��� �V1�����Jy&�?��J]��`/�b��O'A��H�����Q�d��.>���U5���V�����TWս�5�/�����`��g�r=���D^��Q��I�Z�z�ۅ�?|��T+�Ը���퐑�ܴ�O�$���j]�!IN�X��!�ٚD�k��	�E�����(Zں D��T\�C�(�����rL&��������X"����T>�XEv�Yi�={�f������vJ^�YЃP�dy�[�'��,�����֘5���bNV�dL�N��l�قg�0�+#ߪ�Eٿ�����I_2���)���2�@f��t�Y��d�=>���w�I"DK4���RH0y
�ukG�M���6�n�_����"?髷���l�b�nX����V��f��]�>F�G�a1�fȒ�=Dx9F�J��A����X�h��m�-(,Z�����Эaz����u�m�-?��pYE鉝7���Ԕ��O>�6\%�����seeU�oԘW������������uN��;��,JdA����i^q��hCM��޲c�c[j���~�ڶ�~������u���l�t2��`��-J������mE!�ABzP�n����%� ��Ⱥ��6>؏tn�˄�wQi�Lc+,���R/25�=����ӧ0�3 ��n�O������akV
��hǫ�剃LX[VBլ�����=rFC"|�S�eԚ$#t��N<������<u�8r�x4�5�ר�-<a�CP����4/��}XV�rs����W�ݸaÙ��rۋ��z���?�����}�j��6E��g�_-uU_�jl��	(�yл��C��~�I�7����d1^��.Y�IҙF��Gr��1��J���+�aH��x�1\t$��cT���u�F��pf���eee�� 4�a��(����'��ŋ����3����0�(�����@�c���O�;D��r�<���I��&�()iC<d)�� ���`�wU�K��ǥ�����2l~�1b���c%�<I$�ÞS^���OmH�t5���L�84�G���h��U
mzA��C�nN@G�D� �'¹2׏��f[Y�ڇ��k�u�e*��ה��xϘL�#q�i�<-c(���t>�Q�ݤ��펾�}�E%����z��X��w^��N��g#�����s���z���;�B���ر�U����+���[�u۶�`�.[�����+���O|��c�g�y����z�Y)^q����"|��-��z��5׼mc�#|��ψ���$����vI�;A��N�Q���{���@��,�`jM�5�y��F����AH���",�E�e�%�u^�H-�ڼ>��7��{1'�qʚ��f��%jD��j��LD)c<���YH[��ŢȔ3�l�֖�1��,��fb�Ҵ�,PZ��ق� 9�AD�:Ȃ��4�3��\pI��T�3��0�绰���dg߻vݺc7n�jX�>�a��/|>���}��]w��t��;d�\Q/���H/Z�}&x��KDh�z����8l��+@��-f��y�F�#b1L�Aة�F�����9���X�� ʂz__���.	���bo�ڵ����5�� V*U�ʰ�g0�=�p&���S�(���@��玠^XX`T9
�LW�rBS�P[�՚�� @�䩥�b"ZuM�k����MŐ��!�>�׍�Ĕ]�@G&��%.Z�f��j<�P�bT,��{P�c��)���E'������0"y��t��7f	�Ki�1[NS����޻�o�ѱ)��lѨ���8l��i��?�/��҆8/v���탻��20lq�m0§#J�L�з���Qú�˶�7q0o�U��F���>�T�۷�=�������)��nܰ�kw�y羭[���A�^���9w>��?|���O������;���9�#�@���<�cm��n�Ts��4��޵���n:���H�eZ���
���}VSdr�G�ΛPj�X��x9H��&��2�)V��s�HƢ�����z�|�^1X�Ř��	���z i�;~���ЮGm��ʖg�:aL�ZM��L�R�]�Ɛ
���F6�q�N�ŰZ�-��P:�mhM��D�3n#INJ�U\��K����� <_�!Fr�d��8���41��5���!p�DKԓ�u�{w������)����߬=x����@�_J<��)w%,Y�7�a7���ԱJ��ӹ�7�V�] wL2,,�0B�yR~NR��Z��t�dA�hT�%��Y�t���KG�ۚFą{��";�
������3��+���J:��2��%�r��qU&��2q�� y�����l\��+@��>�)��y�lZZS�Z/V�A���Y¼'�Ko��a�\�>)�H�[j��a!׆؝�R�%l��>�"#[������ ��׬D�t�8v_��	\��N��i�c��W�4S��>jj^���w�s�f1���s_$#C�F�s!J'���Kw ��$��tf��4K e�P~N�I:�tT�%:`ċ����=�Yٿ�i��+(*^�%�Ă�:��Hq?�IIa^��i���=�|���w���$�xih����Chy�����������kXv5ׯa��������=�̡�xotr�t8�&g�S&"9�E��F{��t�T�o����:����1�d1<��d�x�� �}�A�
� ŉ����hE)	`�V8u�	 \�DLBꅺ�@<BzO��O���x#�(���Qa�����[��mpd3ӟP!:�y�K"a�(!0c�Һ�i�O�O�2
������������F���kY�K]�4"��0FTT�
�rAӨ|N�L��y�$�i-���Ȍ)U��4$r���c�l�-'N�<�x��w���|��7��a�������^����_>��#͐��4����J�c��ѫ>��fIG�}��%F�J�N��a:�+��&���%��PO��R���.��Tږ��(A�\#jf]�%��3����dkf�82�S�L���m��2���ԣY���"1�ȍ�a?�=�Lc�X�O ����qf��%���[�[���"2�L�_)-)���"A^o��Zr�b�.nG�p
���a%!�Ν���2?K'�:)�@��Agί)��6�G#`��&`n~'��a�;�����W{,�/#?�{�8|6�$?�r�/�\j�%~R��������!�%���֐�.S�pΤc��(�-�\�8Vmk����y���3����q��Qv���ZS�S1ڏ�5���m��yU�=7�䦐�y���OU,��_`m�5��?��ӻ�766������v��y���zl���_���?�������.���������Z��#�k#SI�;qz��9��[75���M���q�,iIc���T���u�<�4'nX#<�5yg�g!J����:,jY�֛��^�&�k��G�y͈qtlD�$����{�%��6�I��>$�NR�Q�[�P#]���=�P�JD)&��+Թ�E��Xa��׋	b��ERU"2�T�I��үuQ�P�XwdC���\M:����#���$.�`Ć^yI_Ki �r�f�毹�|��m}�k_z�����W�?^�_��_���cG���w�ߙ��lF2�2e ��E�o��u<�:m�@7Y�P]��	1r�4<�*KL�̂nդDa�Pk�!v�rι ���"l�����!���
^LQ[�ɂ'�,O�vn��pQ��Z���غ%m�.@�OpU��&��]Z�,��A3�22�T�"Q������=�lB�L�%Pm|fG���N����X�)H��aF�mn�19w����
�A�G��
�' #`�}�OU���3ִ�+��˔��SC��)o��M	ǖ lF˞C��JG�-�{�$�)��h���*��LE���`A �j�Bƌ�u&*�<N:O���Q���s*N�f<H�DYU�b;��؁���@Q���+*�Y��Z�ƪ�򲪩��^��'�x���Ç	�(7MMM��QF ����Zp�S���仛7on/-)_V»o�q������{�������������䴁�dop&-o(���h��������ѷl,�^�Uy �6�ō��f��k��7�Ө&Cz6�,��,�yyϽ�}�����{����,a.6|�d%#Sܬ�u��"����
���#uZ m���^/����䆽[o��G��E���y�h��Ȳ�'/~�Д��
�&ߨ�xa!b���A���ފ�w2AvJ���o��&�K���Ga���m�Т�D���#����W��PN � 0�ĵ��Hx���߿�a�>��_h������������>�i�.}?��\�%�I�ڇq:���MF �#�v.���YI1U=���ET ��a륖u��� ��J9i���j�S���P�R,�G,��!�ak�
b
f��ߙِM���m�� ��gS
���x�V�S���vLJG��� mg�
J�Zt�l���s AΎ�5W�8	����B)^�5���d���e��.�qt���ŉ�:��(S4i-��c�'m�cڜ��^ /�V�m��#�&j�j��ЅH�n�]��}���N�f\$�d����y!G�5��сe	��8fc�=�k��#^��a�B�)v�����B:e�N��S�td�#X��y�~��kU:O�Λ�:�?|x��'���}ǹs��ߎ4f�errs�e�x��iMWw�;�;~?t�ܲyK[~~�U�v_�嵶��w��o��D��G��l��y_�������J,<3�7N�F��M��=�>�u]���������^0��K�M1m=�HX,
��)H,�$	2�P!�<�<Sp-��J�KJ�w�x㗞ݷ�����K�R�h��$ƳO��,t3���)n���p�u�yU��^Ei�w����;�v�!iScJ�1L
�) ]���X8�Է�,�~�(Y�i8�lǎ	dz'1���9.0ڧ�dKL$VMu���f��m�i-)	�:��E�~���45H�4�ԅ�H�}1U�}��� �E��LE�?G��>�����[����~�܃�����#H�}��/�Zs�R�e����m��o`�g6R�<�~?2�,u.�6�*cr�<�t�$3�f��c�f��&�`�јJ�2
�=���^#A�A �\�6"���X�A b�9�@GG�?�e��L�9Ү�ط��d�(l�`���/�t7݀v��iX�N�~�e����2��N#@y���p�9@��c�
�OD���8��<F2�"�d��LKs���vC���da&2���yBV�#���%�1S`%ZU�uQS�G�kԶ���(T�f��܇���DZ���v�-	q��ȵ��:�/����N-���t/FDy�o4:2$Òi�#���B�%,N�s�^O��A��������y!�.��U�gbk���>��f(�.���Y_/�=/�K.�����ZZ���=�\�5?q�B�{qo�����e�=�H���>��a�n�喧6l�Й�W�����;x�����]??3��P^���e:Ƌ�A>�X_����l�������9<�x�Z���x�[�6��9�HR��2-MO�\&�Ģ0�8[�����[��[��y��'���������:��|���+��W�<e������8��X��R�QC��YY�`ΗyE��1�gN7z��Ͱ��Y�`fk4"Ma�kJYǬ*��.Č<��'�Kf7����?���}Ӈ�.\�(mQ�ʕ,����˭M�[:	��-��R5�M�S�j�^i�"�Nҵt����;�G��5�#�����$lw(;+��vl�~�����������;�7)Պ�8�pp�dT$�P�;���ۆ�"5�b�2��q8�e2[B$��$6�1��}&K���s���*��`�1��C����uY���D;]�ĦÀ�6��t�)�ݎ��DFn���)x~wII��̱�.�دm[�bP�D�|o��ΖK�2�Y���1�y%2�b�	~���Cb�u�-��E6I��~�F�x��L��(�~�0����N�'���`A��*΋�Q�_��$3�ƎڝO!$څ����m�ԯ$�ϲ�MRM��F�<[ҰY7�W�q�<Q����0È��-�u�+m	��z��0�$G_T�8�/!���)�K�"� �&��Y�L
9؎��x�"�d�d�4	�`~�xii����ַ�����r�֪�З����,��=~���ڻw��<�ː�}��T������dᢹ���[/]��1��z��'v�_�����|Y �m;o`������>�{��_��z�B(�b|!�&��d��^������|�ؗo�ڰ�� }�J\�XL&��6��p���eq��2*���S��m_r(9*�eX<S16t���O>����x����"��4H3CiFJ\H��{�s@a��(eG����1�ks ���7}�{b�^��<��&
�� %��f$�2L`~���^XH�Ȏ��<�p��Buǝw�Ĩ�M�¬����d$e/M�M�RS�:uNS�`iSq�uF2�uXB#�ĖM��-�E5�pYܱ`ҞH,~� �;�E��駞�HEE�#۶n;	@����σ"[��h���2s@�@Ϝ�݂Q C�� Xj�>�hs28�S:�!`�F�ƅ�D.F�X�	ܥe�`�W��P D;:K�h�$�!�|�D��?��d?�]��om�V<�����Y�f��x�ȵg@�@�l�8�����1�s̄p�D�����^fT�:Jɢ���/Β
w�6x�cAM|�g$k��<)Q�q���f�h C�e�I���������Œ��gJ���3�`;	�xYBۿ���%��E�י�
h���8۾t-� n�u��=Z�X$��.�x�(��@� ��e�WFĝ)��~�h��tp9O@3X�g&��k��謰��L���>��m���y8t2|���eR88Xf.�7~����BqqU�����_�t>��3�hm�9t��/�m�����"�3EũI���L�{<����Ȧ͛ټiskUU݋?��+屧�����=?y�R�ǣ�Է��٩��\�8s����(7x��4��+����dFZ��\/�@�'��v=����:�����@Z#�	�li���dp�I�А�8֒���C��{��>�?kimY���߁'_�CꙒ�Ԏ�[qam���H}z5h޴Hႍ��'he���r���Q|��'�"b�B��lZ�\�Ù�*�����M��ma�L�c�`Y��<pa�O�����6YԄe�EV�hF�S��D������Z6FP���j�[P�t���¥��(��H�iZfE �x���: ����%�:u���v�(�2������K���]S���*��)cj��{��6?q*���D ���C8��f�X��ږa%T���ņ�>D�y�5�˛62+Y�D(]�����f<خ�t��8=<L�f :��H0ق-�CH���{��Kb�LL�����T���:���	�l��9���0�%|�<�>z����F02�}��VD{ `�sX�k��s@�d9B�n
!��%��Ì�L�(`U6R�Ot�4��D�ǔ�D7��������8�[ɪ�m���K���N��2 j
�HJ��ejzB�%�7E�]�	2UO�%�TR���	`F�d#21~�1�Ψ���\�p�X��ۋN�qФTF��Yǰ��07��7ly�%�/ci}Moq��#���s���޳�i�_܉ˤ@�k� � Y�1	��u�6�<w����������tR��?��{6>���_x�,��f{sP����T��������-5�_�is���U%����O>��'O���^F�Y����(KF�Gf*S�L?�]�7��zd�C�}7_n� R�� <~�X	�	���	2�`4�c��w,�����8d��L��΄��]���8����޳���h��29�Z3��p���h]D��B*5A�'��5�N����S�t.Z���;:$r� ��b�jThD�ZY%f4ugy?J��������VnU#CU��hD�`EL�*gL�cq��0���О�wQ��挈	�&���J�U��tεD<�\��Ϝ�s��s�M���$J��Ju��/�]�l�̰̄�2���\�-C]���Hu{�wPP���h���ۃS("��`aqec;�zUҩ�cTE;���r�E��P^ �  hI��5m�k�:�$��&��83-���2g/=u8*��s�{ҹ$�S�8� �'g���P Z��8^�J��~�O��m�BA�8<�*�?�']Eq��ۼk���t	P�^:miK���-f-�<�]��$t����XǦ���V�����A]R��?K����K�8�JLeF| 93('!�W�G:�t�y�� �	�W��!�D�kt���m۶��Դ,%�^'�q"�|�Ѳ�{���X�/@��-�֨��*֩x�P�����=VSS��-[��B�UVV���{(�<���>59�e*#+��=�+����?zCC�7���:Q\��������ٷ�o,���S�|0xL:M�*����`�)$����%\��*�2P�8[�NL����M �$�~�w<PZ��;�t��}� �tx���3� �yS���{^�I�F���hӲs8�h�
�鬯�T��׹�g�)�d)�b-�[ J�X{��%��Ŗ�:)$�
 � ��`a���%�?й�*J�&�R�!ёxg�r���b�z�z�(�'�S"v:�$�a�eZ��j:4��E�6�2�h�@�Z�#�Ŕ�8��Z/V�����m�$#�L3ak2� � ��3p|��1�Y��M:\j�TUa��x+8�(�~��m��[�4�D�Y/t�ې!9s�D�R�� :<�>I�|�ý�m޸I@��a��ےs�t6�[�j�a8�7�9 ��c�w0=��0�}68I�8���⌀#�j������^$*WCW�Dil�vXꑲk�r�z}X�X�>8�/��^|���ŚDu�M�iQ���x�h��RP�P���p<� ��E�li������r\CL�3joo��Z�Z���6Q�d�#�q���n!J��-����w�>G9�'��w��\S�5S���.��Y%:hp�N�������.=֕����p���x�<����lچ���FaMۍ0@�-SR���7bl�x�@��u���W�V�v�eo���f�����މ�������2@V��U��Pv�PCU�׶m-zp熊�<v�ҥ�=��g�B��3ӑ ����I�R}��l�G�Z�Q�t������^�d�|��5�hr~�j����D @9I"4,�q����E9J�pB���F�2�S�4|n�i�� �?ᙱ�	f��T�T�*7�A#��	����;"`8ri������M3J"�Xa(�a�GF�Zq)�����ށott� �D>�b�%Y�r9)�� o��M�j9p)��i}�S#v�bF��O6#��H��oؿ~�Aɀ-mS��WZX:	�� Id��_�����Z����[����m:X���F�������[��嵂	t��NP��	���f�&ii���n��ۺy���հ�Z��&�?R��視=���Y͔��/%pL�3 ���܀�AR�Y���>�"����^���Ad{/!��,��Ӵh�j�κ�xb_���q%؉�#�T�x�2����N��I�����Q�G¤��e{.�9�}����m'P�Ɍ3&<&[Cb�J��x�-y�MMPl(-�!��m�����A@��*1T��a�:�%8K�pZ��Є(�K&�UOn~Wiy��m޺��I�;@�ȣ�W=��3�|�����p��q��ԜN�B�s^�x�֮[��͛�4oX��;?��M���{�����̭';~qb>�./���OΔa�9�H�6\����ƚ�{6��>����5{����}���925Y��E���V����~FDa�E�7�(��Q�Z�酐ue���WT��w��,�`M�8��+��v��S�ߛ��땂�NP�D�O}w8^�Q��mo��g��>l�]#G*�.z�U�]#^I�rF��Q0Z'�3�	T2p�0+#Q	�H�E`+��i�_����x ��������<:>��P�Te��'�L�"��_"x�0��Zf�um��r���j�M�p��Ie����5v����։<�ӹ�K�k9v$��ED�^t+K։y�md�n���="�#�q��miK�a�`�miԹH�j���q�f '��;s�;��,�1{�	�lfU��2�����r��B��K7��X6��Cb�Oi	co8�l�3@瓬~j��!���Χ$qYY)�Dq�CE�;����&�.�si3#��1��[j�f��T'�t���1����M�k"#[UC^�P+��~$BW[+�jAܖ����0sH�������i �~N:&����� ����q�ȏ��]N��k�����f�ao=��y�
`F%0ɘ�� s:Y�B��`��P�O:f�K%P:c���Z�l�>�ـ]� 3��k֬�Æ�;_,��8@����f8����soC��CX��6WNQB^̖��Hn�k'�FhQ?�u��'��ֱfͺ�7��o�_��j}��'��&���m�#���gos�W���f&�+�Oݽ����ז��T]tY���T<������)*�DGT�زD `�p-kqIO"R��Lš-�288����5�ftKF�,�l����E�5igC͎YTF(��XxX����||'IrY�f�ј$�QH$�H����{j��Rk�D�a���HP3�M"^��jz�파z���HXG����i����Γ:�k�K��y��q��/�/<�o<ߴ���3���\z������H�ڶg���MQ' ��/ux������؈]3G v,���͈��[�BJ��0�):Q��xr�5 ��ܞ,� Q~��^'r)0���w��?��se��u17���AALeMm���2�ֶtZ�.��$á��BB�в�ȏ��1�Yuw�	�� ��}���6z�$��1.`�'p�FNG��#U�C���!8��Y ���zyx |���$�î������3M![���B��ԁQ�f'��Q@�m,AMsC	�Ŋ&����{-�KĪ�C@�s�\���t���T=�Ex �t!΂�����?�k�*��m�>H��kD2Z&��.b=�!,����O��)���ÌK]d�㞃S-�Sr
%s^:z�Y��g�����9��EPW'�$O��(�a��}��������]�.��p�~�N�|����C���~$���[�Mg��4\���A�j���ۿf����o�~q횵]E�|�ۡ#G�}���Ϝ��3#���}�k�\/_F&f��,dg�^��?��*��-��'6���(�������CC�(<��sz��Ĺ�3]Kmn�|:��9 t���4#�OGԃtx���f{G�,���� j}��Ց�JX�݋T<�e!:�
��f���^�u"tD������@T���缳gu�`�)u����:5M�E� GJ��$sۅD�h�GR����s����� �,�b�	@�,���v&++���iD�E��OM����6��/T<�Q�={^ZߴS�3�`{��_P.�ֱ�p���i�H� �֨
�M�Z�%�Y�����7c��� �B�q�.-\<9jSR�\HM��2��=�Y�M�d"�(�qCxcZ[���z갧�Zq�\�pAH�� �(2?t�X"Q���d�����|�Ll�}� ��ˬ�OGg9T1���VH:<<�N1cQ�H�e�{����mEZdN�p�lI����jyb�0�@����b�Dڦ�!�n)���S�_�2�7|	aa$@W}��`� �u��1��K�q��O�n���ҩ�ׇ=GV(G$��CA%����ַ�XJ�����EKj�dA�A.��CWG�9� e
d�][��#�4���~gʞ��Zµ��x��H�I��ҡ���ڸi�H��g����}��~v��,���2��w`�X�E���A^���*k:�����X�]�a=#�֭[�����]���?\���v�u��ѹ�-��K� ��è}gB�)3��g�Η�e>_[���5��wnxuF��G��x��ѯ�n$1,����J���"R�*r��=*�I��>����/�`��LZʤv��Z��΄Qkҩ�v��PO��ଡ଼o]PX�h�Pz>�xbǼ.(�?u��ǼѡI�i�ʃ�*d��e��utQ�0�����nm�����/���c��x!2��4:�� ��X,Z����C���`�1{�ԱU�Lu�,+����Ч9���S!M��B2�t7��̊��M�\Fp0�!@���o6�s��f�	Y�%=nA����B�<��K��txF"��8�O��&��f7=�&E�s;L��� e�r!O ��	(�MW�8zpn�l݂�Q�q�Ց�!�O�d6�pE-�f�3��	���I�������7�M��־)h��«f)�,r-H[�a�'T)3,���x��AH
�uj�*��^>�����Q���Ȝ��Y �˓����z*Ϳ�D�32���gڌ�� �0���'!E2�֕l�!�_j��+�6ro�4.��(@�e2n���!v42K`�ML`�=����I�@�8V���O!���^����؈���?��{탫+���[�Jm�mg�N�:8r�H9T�6b���FGG�"*X���В�H$�O��&p��^|����!��Ϣ����~�ص����ok��?����Gc�;bl�AZ�L�DuY���RC�9i�gʳ���+�US�{��8�Eم�g��>������F�����(�Q	�m�(,,��/e[Y�b��Qk�d��aA��,��%���:4kh��^�D\����-a�<D� �!G�,�[em��K�S�mg#]
��7�tjәF��C�%k�M��d�!l�@��)k.B�]�t�����ں�"'��`;:!<��7Iê��!�Tң����?x\<nQ�"x���T,�V��%�I�?/�o�'.���f���K���6�h��E-�\�V��FwV��F���$j7љ��m���t��O����͙b$�E��tM��4��P��4���>�0�b�#�388�ȼ�;q�ԳYGf�q-��(��	��:B�=�#KZ���#Ã���cF ��BD�E�N�c�:�Md���ۢ�g�X�6;��ǋ��	�C��:td�n_J��ui�V����u9�*�+DH�<eR�a��o$ˉ+ُ��f�,'!�2_��X�A�(&ʶ�`R�gT/
�p���m�����%q��:J.d{tm�c��i�r=J[�a��a
��r
2�^/�j�p�E-���K��bF+^zܑ$�?i�G7#�ґgH3p���-�CWү��ǯ�{%��E�WҚ��-wIG�^t��ٷ���|���X�Jp+��qQ�����y�l���Q������ׯiFkMWMM�5�<t�)���Gk�����;�����crV*��2qc�F�@�9/3М�xdmu�w
3.ݴ��ǚ��������859^A	F?dq!`�J�Pvf���2'}��:��ź�$z�TۂR�D�eDn��K���қ�dU�EcD%�^,��+��F&�<5��Kӑ-0�o>E��ݎ棈�XPĂN�&e��)vY1lmK@3�9F�"���X��/��t'�d�Z�[|��N���U�̲��>MY3e��qK ゜h=�@�QҊ6� 7uDFv��f�vj�N&�K��u��&�Ut�M�[p:}���h��ly��o��أ,�_b����G�_�����LD�}��r�X���AnX��N���#��&��ܒ�A�a�3+��XS�b�U��M؉�^��R�Җy���HxTA:t� �F��F���ux�!2�4،�^�F5�\��aYL��s(�:lY� 6ԈZ�b�ŜKL�4`������K�$>��DXǋΓ����~�r�2��� �C]su���=�
��:3�����>p�D['���0��B�kg:)��!��u0������t�] �v��A����CD|Gkf���Ug��]�g!�,�;5ġ���u�$&}w����f͆���s���~��k�+����WJ�=�u��Bun����1z`4��."���75%�"R�׭]� ��jk�ݾ$ve��[{��c���;�������9��� �BHŧPa��0+GN[afΩ��������/v�l>y��?NNm���{s��0�-��0�Ù^6R��L�Sa3����Gc�l�Q�{�ϐ�"�HY}seq3�̅V�Nٿ�� �%�G��>X H'#�"S^��"�6Ɉ��H��(�d��ǎ��p������T�_(�|��!c�4�%�-ѫ�Ie�Ґ�:�X��R��uS_�����(@�a�,���k�Җde��ĥ�*�#(��HbZ�m��n �2��~�F�K|M��`��Z6�8Y���:A��W���w����cI�9���R%�I_8���`��I��t�$ڴ4��z�^B���%5Z�(h��^>E6�<it!U1���7#�̧�e�.���=��C�Ip�,�>��\(��&��-'P�G�Q��^g�stВ����r>��wWV8I��B'�/�7�?L�(s��΋"t�[c{����;^q��3�����E���:��4�����y��B>4��D�#1�:m��!a���ck�1���� �|R[(��g)35c&N�T�F�!�5� l�F�0�!0m 6�uߏ�᏷l������g���Wy���Z�
�oף���9}��ԩ3�Z�P;ވ�d)�,Ә��C$eJ���m���;0�2�3�����?�*�?����g�?��LS���N��k�I�T}aOs2X(� <3=e2-u�LFj����������H�lt��@6=��׈{Y �L,��Y$�
�hr(@��C훑�tDS��`)�9ą�]0*T��i���p��ysJ���Q%h� r>,�>l��
O��{��G��@g*� O����!)>��a(HzeB�c�AJ�o.�[�K���Ѩ��`=Yd�%�!I-S����u�Wr�l���Y�@#��4�+M��n��n�����\ti�׵uJ�Y���:���ɫ�H�L������#fFu<���8*�k��6��þe>��8oooC�Z�����U�&'����M9P�`�&5k��n��FQ���ђ@Z��a%}-��j��ܐ�t ]���oqj��Ҿo�3R^Yt�x��o!2�0CHt�;@�զ{��*Z�Vg�<���`��3"�O|����Cs%�w��ԩ\�\�X�%�bH��˶^�������4�@&@���!��tF� �T��l�y�9�aكC�$���9!\JFL�Ct^�>f��>�2���cj�Sڨ I}q��y��)/�PǨf�!������a=��d�������O���/9�e�O����sϿ�<����;�G����^��
7o
q�u� z�Y��=�(����X�vWVVR��?�0�b�j��gN>��ȺC'�}��o���-I�P6�]lw�KFK���x�<R�9$�mQT���R�d���T�������8%�2pl \�!A	�`�(�1��X�D��iw�X��s�53�698�Q^c29���Q@�<:|��'Ǽt,�uNb�+F������3u�*,�N0l�Pk���ѕV&���TZ���-Q� �h�%�t�ׅQ�Q��+GI\�%Ch��,�M�Ť"��u,��)��b��=�ӳt�l�I��@j�l#p���t*��-��o���Tp[�V(����d0#/�Վ��T�`�~N��x�c:�ud'R����p���*���I`%PDl�5�;�ӫ(/�(�ʭ�P�|<H�̄�8S��p*�j�:�S���߉ӭ�i]��wH?:�U�&Z�X��":�]�w�ȓ��`N�a���oy]��U���@�ɿS��Y \c$�����$9=Z%H�F�mk�0�e�u溳}��q�e;�Ij��I�$4S��q5+��H��M�N�	�k��{L[�Li�%:F�W���C!���z����7� ��mki�T!g�e� �����끙�\���'����Iҙ0�}���͛���vͲ��a�����X��g��g�N�:��ȑj�>��͸qk�pL�wJo\���`��nx�0�k?���������6ԯ�*�~��������>�����''�c��Ԛ�$�2n�#�$���%��˘�9��~F�`�c!�ca�����{�d.8 ̰u)B����"���B���`2Q��Ms�g�����4�pa���QŒԯ��XȰ�Σ�
���8�f$Z"��]���H��03���,�XĦ���lnC]�WYY,)>-O�U2qͼ8
2H��W��R�l��,��f��;ˍ�$���Z�>�?H��,m-R�� *Q��.M�mA�)jq.u�ԥ;b�Q��2/ەz*^��gQ�4���(	r����� \��*�+p-�vC����u���'�9; h�DfhK��F��a3
�p����6h[��?p��^)"t�6�-W0����f�
A�����:�iu�,�Вפ�LgSj˚MbiM�x�ΪsB��8�8R���*�PLm���7��f��?���Wu����(���k�n�N�RW��:aJ\Sқd?�k�8�j�?��v�����v5���~�/�$t�mffb��CF:e��$+P�=gk�f5Dz�L)eq�󒥁�Hs�o�N�l`��#�����)�y:�VU��*U�T��	K���2��m�wܟ����:X∖�/З��H��#�>:}�tIcc�ږ�ֻ0�d#.�uH!��M(i��7��>��E�����s)';�paQ�AD�-U�UCe�e��5�cW�P�{�9���4�;���ց���x��2�?�'e{�D`HMS��d���BXD}x-�d:��ĉ�=�
-fq/�_`ZQ}Rԝ�DH����La�T)j%�)���H��DH�8A@�n�2v�S���\$[%#�@V���'/ .J��c�Y��� � ����R�F���7x�eh����@bCT�a����X�F$R��5�����dBY�l�ύ�[׼(�����gي�ȟ�*���ח��ٌِ]�%���}�i�/օp�C�m�=�غ��M-����5hn��Lr�s:�d
�I
Q��Cn2��2vC0R��<k��C�_Fr���v��Κ2AK��Q��������~�'�����.��K�@�җ���0׍��!+�*���
�G� 4���=��:#$5F�*�Z�>W &�@����̆�H�˔=v�>h/��`D�t�t&<���r�:	�r���Y�6-w��%:W�K����,����t3�US�d�+YT ��I���U�=��B���2�����q�/�_tV�ʼ���y#����aŒ��a��AI"��H�}�E่B��5����<�L�3��.ڊ��4hl���w�iX�k6m�t��Ϋ�=�W˲Wp��=�H����'N��`���q3�z�o�q���&WQ���r3��Ci��~�ut��y��G��ǳ���������z��>������h+�����T4u���B�|r8��]��\>(�����jX8�m@��]"a� @鿅9�o�9�uNT��li���-A6"v� ���D�Cd͊�4� :��gx�$�h�8��d�o~Z�\�%"�����D�r���������DO�75x�{��2o}M���e
�1d/���d�艷�u.�S�D�%��Hh�M��_|K+�_��E��h|1ŭ�������c��:�Ck�6b��mY[<f[�&PI{�2�U��@W���(�� b��J����>*�%�K=���ّ
��0t|^�NI���c�<�B�������A���~P����� ��Z�ukii@��FV�����Ԕ' �V�N�NU�SgJϷ���k���iR��yM΢�BSf�&�'���%Z疩vqTنe}L��Q��V��r0�pHg�:ez�mJR�.�%�Hx�"8��:g"9L&>>�$����dD����6;��خ)�P�`�l�l>�G���Ѵ��0{a�q�:�}���<�����'��7��ɎmF�2�Vd�!A��3�b��9��Ŷ:t�as8/7��o�馯f��]s��;��s�~��Z�|��O�:Y�Y֛�fz�5���q�T`���%ڃ��j֪ �q0N�ѫم��	ĺg�+ʛk��P{,))��P6~�<�\ታ�O7^�|���桱�M�xh�?��7� 0a�%����/`%] �&�'SkZ���/cAu�%W
���3B'�Z���h�L�H��d�L6!,$]Q�2B#˕��HQ��=Ű@����i�Gp��.zѱFﭛJ��5�q�<7.&5jy���Y#$:�p�kK� :&K������$.���f���&�؀����f\�m
����۴�I��[�Z=�/Δ��I]������ܤ	D��3�D���v	�Qr�֣a�a�Yz�U�3AQ�aH��O��1)�!0�'���Z��ˀ�|]�~�������YL[# ڱ�tx��3���k.�����}^ ]�L-��Q�5�i�qjd�"m#����>���ٚ��kc)q�=窒�&nG���:���J��A/l��HU�`�b�=���
�LG�Z�>�Qq�����ө�}m)[
�z����ҕ���y�z��;�O��_&�$�-�	p*XfђJH{�Knƙ�bާ��S�C�w�F�"$A��p�G�}"%��k�θ*��ޮ]�Hm]z�Q3�%�
�AL�M�80J��ZD r�x�H�(3�0�=����7�O|�2���2>9?n���[����:��X��@�|'n�z|�B����X2M�������R��=�4W;R�����2zo��ڗ��?�!W$�?z�R����u�>���/v~���*��\;�Áe1<Yw���Ƣ@�f�N���b�VR���:Am,��EAA��[��Q��V������g���bj�U,vE2��:�B-ܦȅ�� ����"���77x��d"��(�ͺ�����`yN���맦Ry ��Y�V0]�/�.j����r@7mEt �&�!�2/I�ۚwb����g��,���9R�V<K��.��7j�����㕔-~֊yM�\�fL�e'�4R��e��1z!�S�rFm}���W�gX�a���e��dh|�a��w��Ii9d4,��c�1��[��᳑r�{���Q��eC� ��HX�?ڞ g���k��]`������8�SД�ƭ�L��<a�3�t����,�B��(�1:&�Q��S*�d"Z�����k�'@G�9&,i	�{���7Ѹ-���\r��L�Ԭ����%�N���n%��1���'�-�ѕ2�C���/8�3g;^��aȒ�7[:��x,\������w�W� �D[#��v�<��2o����<L��g2���;�x|�B�k8���4�;�&с���@n���6o�rAq)Zu�����{_�޽�?�3?K�>{1��j��Ξ�Ĵ�;'&�7A+��U�;��*�<1�zq |&"�����zߋt�0R�� 
5��>wϷ�y���������_��o�P˻���ܵwMunQKG��wv�!e�f����f��~M����Ȃ�5 �O����h7=��%�d�A�V�k[�YA����y���A�]#o��1�U�`�+�I�3��=��
�	���9�;�@e�F:�'�`v{w�W���)E�Ǎ�q;�=�t+�*@h[�'�����F�Ky�q�#�o�/i:�t$Q�2�e�ڬG�u��'%�[HfBvM��dA�Z�}=.>��O"Y�:��Q������ �x�=�a&Z��jk$
����J�E�G�dp��+�6V���m�0ȩv�\�)����h��:fz�D �Q4�K�E �D|�	pR��L���sNA���1ɵ�z5�i�H /  n�S����ɯ�{�������g*yDKfT�Ő�8�4%��18��M�6A�����P�������#d:��%#!>��y�%� �_�����v�X�I"�3].��G����!;��������E� �}Ih=�|�+��܈��.\7xQ�3�F��ɬ?�vUq�f ћ���|P�=2Ko��k � �ȘU8`�8EEd|�̰f�rF�'>
��c8���w�V�s�~�,}���w��hBu���G�?�x�1���Y�P7�tw�Fc�pT��yXdR5��~V��u#�� ��Q��	������"���g���%%%mxv�U�b5�u�y��8�������m.+�Fz0:ٌ��e!�D��4�Y�t� 2� �<b��<Q��G�p�d�t�f}�BE���U���L�����D� �aa�SS����69Iyra�7@`���lWg_k@���gƼ5��R�e�����*��4�^t�����g !�	�a3?*B�miD)uX2җ<��&I���	�*�N�I��X	�\��Zj��)��hXr� �|���"��'�֦}&���4:#O*�ȦAt�"��i�ʆJ�����	V,��
�� ���AF�\l�c��d�Z�ٙ��� 9�]������Ť�F�v�,	l�����۶:��,�OF�L�RzWR�&
�a+�@��ul!ڑ���Ȥ6�9i�q؂$?��!�P��F�l�b��2��N3H n�o�cZ���m�)f�[�%����c�*����M�9t��\L����vT���Ėx��S��	��\H-�zz}�5`����R��i�q���mo�K��y�����O�#� ���[��Nj��
-x�U��w��=��;�
d�<	���XN�~�x�$/J���sb^O�`p=���c�����+V�|����^u����,?}�����>/>���=����P>[���C#k�V*�\�ū7g�i1z�|�I�Lea��������# ����5�E������eR�PL@�}Ӧ�s����\q�6͗�����Ɖ�኉�(��fƍ:9�z���{�X8� �$U��e��VF�I���w޴6�ՖI��d]��3�.�q�hg�([^��s1 ��ْ�t�F1-H�>=ڴ(#�r�mO��~.��9� x3ϴy�F"x�H����]���'n��Ņ�k��@���.���1�c�D�F�K��D�]"-;���bM]?�iI]XmT��%f�l�D�M�z.�3}*zi�Z"x�f�x��#:�S��2m�g�Igm�v�~��8�W8d�WW"���[)�GI`bO�f3�G��f'�v��+�
�sB�^8��~�@E� �U�#�҂�����c�4�jE�����0�/���@n��e{Rs7up:�}#th���	���S�������M�m8�FС`��\F�"]��>u˩�د�8Z��E�E{ڭ�',w:&�e�s14�/t��ڣ!8�<��X�n�j�e+�d{��y����S���pr��Uo��O��0ے�k��{��O��HRD�:0��(�� 'r���,�!��С�H��:A��C���^^�Qd�R��[�֭]��A*���p-�4@?:[�Ol�������\��۴C�����r������+��$��%��������Q�N�<�ts��lL-��0�}}��F,B帷���3zO����)���b�a)(�bS�Eg=��(��t)�1�� �a�d��އ�~��jW-s8����;ں����724	��",:`%�&%hh�Zm��J�#�G�˔�M�6����*3��Y��D �<� S�����<"�$�|�F/�ơ����5�7w{�˱�Ndf�G�k�S��2w�}̜�F@'`��G�tQ���e�˲����ES�mAބȆقӬ������V����u�6u�]Z�DQ�@1U�L�D�̚�X#CF/���HX[�&'�F��4�r�%�M4�ah8\����z�xV�W�\'�f �� ��֫�s�P�*�f��caj˪\�Ѣ�-�S���ؖqO.���_̃��:���綘���tn� ��%�@ �d+4C�6�585=*R�:xB@���Ibl͂󐟧�2)��>nr[x��F��
����h<�����>�{	<|��Tؙ���є�( /�(�Wf��Y�p�׿f���nKK(��J��{Ѿ׶��s��ed�(�p��^:[*C�N�E���d.���l*� rn��Jfw�a��f��i�����rf6�`o:���L�c�8��7������ߦ���ׅ�!�<U�$���n�a�;c���u8D苗���Ͷ��-;lݝ�T�������N�<Q��ѱshhh#<�r�|��v��g�bA_�m`�DT�9::R�E�-h�=\1d՛����4�%��(���\`Y_����!����4W� c�K��b#�)����-����/" ����h�D7�ǅ0?�>BB2��|#?�DMʡ�a �J�#۝)L	eﴅ'i!ݛ@k��{����Q����>��e�n�3��օ�⦍v,�[^��_|��Ihi�ֺ�_��XDҦ
�V4D����n[�q*
�}�
Bf"��H�Jݘ�'F�/#+��Ա
�hY�p�\��p�,�WZR����{e`�����J�4���e��gWC���)�!{,�5'e�k�u��1.��ړ���c��������Z"!���4�)NQ�<+`h��:���T�'.��V�x�S	L�N�uI�"!K��X�9ݙ�JO�ayv�h������3��$˾K��\�G!��}�z�p~�&@�A'��1}��8�w� �l�:R�zYt#u�z{mi�D4L�_�_�,��N��)�v�yg�O8�~c9N9WF;m������b��z�� T&��6G�>Y�sIr����-�:KG����ף�"�DY�H9�v�mR��I�Y�i� p�<�S8�2�ۢ&6��O��##������G�U�z�]����"��g���S7���q��/6=�V�L���Ϝ=S�y��0c�f�d��n@�
���})�茋��]#�lD����K(���͔*�Đ��MHfL��rDfz�.�	�h%��(�8� G�.��#�	��adg.?X�J(gD���Pś;і�H�5z�Ktb�SHPx!�'���)n�d�
� <��EJғK"p�Srl��� �ҟK߫`���m�����iJT�u��k�mH/�u.Ό�y.�*&��`�c��Ia�FBR��Ȍ֏���Ա�F��*���g ����Ĳb��� �`)#:O���EY�<�<ߦ��rls��:��L�D�h~��hY�z(�H4��~.�Fȁ��	`~a�3���	*j?5��t�v=��UC^g��ϝ�
� ��q� ��\eSsH�[dU�z;{�CP���>e�y=
��#]K%r��![zm�6K��A�{�u�4[�c��ot��u��7��7h\Q���
A�����xI�mm$�א��s{b�EgQ�	�[�-q��qёI8�̂�e<H��$������� �����ɸ�T:aP�c6�DV�,�/haー�4ؙ�fƏ�#�C+D�k���m۶a��~q��݋����6�>�9�?S�b�^xRjb�+)�����+��҂�^[^��[��ݐy���g�=�������/�C�|mOo�x��X �F�ƢW ����&7 \DNLc�b#J��+�1B����W��%�_�ZT�@�FDv���ϭ�Ӗ���-J��~u���?Xzu��d:ls��;m
A�"4�A2i`@Cd<�y`T�Eҵ� E0���3�c4b ����T�>_��(yʿd�\����0�@kĠњ���(A��$���R`������?I$��#T+�T�p���~��p���,nL
��Zd`?hW�a�/��5"�Q\T$���*0j���mǁ8>�
������"�n�u:R
0@o�Y6�U��M=[�W�5@�w�~	~X�yޙe��n��I�#W��!�B{���̕���~9h{7�.��H�C�$2�y�����r�ԂU?��5".VAϡ�1%�-gl�h�7�X�
�ؙ�*�d'�i������w���6'O�|�=����~��:�	�O�1�ʾ�S�2�ͅi�=7�4��a�kD�>q#(�VT��\�*��� Y���0&��r�)��!z��db?��$�U�tl&�wN�ﹶ𳨩ϡ�e��MayPޔ��SĠ� �1c��DgQjD	 ���ej�r�쌙���X��u��E���d,�]y�m��~�y	σǏ�A�`���3���;���^78п#F�`��(b�Z��iX�3 �a���Q�c#��f�.�x��₯ �;]#��d�c�ϛ�.�:o���m�
��i*�2����H�]Ӌ�� � 3=�ҝ��E�^�s�D-�)���,I�ʀ|�2�ul&�� %����T\�$������{�i�G�\Aɨqљ�sd�\��Ff�^�D��4��9�zF&A�EU"T�2 GIM��mIUV�$1�T�H�\X��Q&�Ir� *�T%��tth7�L�3O;�D~Fzr��11�T��.r3vԐ��8�wA�Y�`af��E9����=�6�e4
���K�O�<0�K�Lcv ӿ�N	+6��Z�� i�a��4 Hj:�nD߬��N�v��D�t��ͦ-PD��`���\<�"�`��D�����_W��j5�-{\�<��E߷���x`f�}P���`׸r��䭴N
�s���37��8!�|��B���N��y��"�+[Ť�#��85���6I�q� N�,s��H���>#hhk�0[�^�������õ+���7��a��	b�q�y����{X?ߺu�nii�N�^3Ft�	�A�����:��F!����.,(Y��q����~\��m��T����/�}lxp(�����FJ+��t�B뺺zn���}+^�4�|@m���������h@�v\���e�ʔ��M���+�##U��2J�!fa"ti��+��H�̅��;�+�.A��I��EFi��n�H���>;(D5.
�(X2���y|<�������D�iVYO�� �"�)�\]�.ER�y�m��� �I�s�"zBb�N�%jь���%	�=��7>��q��5�G66����� �Z!mC����8?��eDj���p	ύ�iΕ�$:T W�p��.g%A247o�|��0Q�� 	i}a��vRMn�=ǲp��ʝ�E�)X�V9ՏC_&@�#���d
;-3�+ �MR�@�����A�8����Ŵ7� ��&ã6����s3�̀�8g�vv���?L�K��B�cw�dh3�/P{2��N�������w��K��%�#�A��ID���'��l��������ZI'[ByM��G�w�e��r��!�q���:�b��1kO�\�ԙ`G	����*(k��vN�~$��N8`�l�a1��Ȧ�I4�c��$��u@GǇ�R:Ar_蘒����#� �G	�$-r����KC��}|l4_7��Y��/З��X����~���<��gϞ�}��'?x�쩿D���-����I[�0D+�p\��ۚ�ݘi���("1?n|aS>oN�R��sf�iqFKd#�&�2Z�y�X�DV�=ҌƐRE�>R}cXD�T&޾Jz�C��SD?\4�����p2��2�Zה�>��,i���~u�L}���V3\�5t򘭧J?8o��f?Zֻ�mi[[TuKD\LI�^ ���Ĭ%Y�2,Q�]"b�qĩU_]]�tz� 8�#��!��[}p[�ly@5�Y�X��`ZX��I�Oql���YF����������&��H��o��8���IĨ:�1?H�����|tvuz����2�#:1�'Q8�����/������w��@:�FWH�<?*c�M��`f����
�h9GƵR5�3X����������a[ ��IID��lI���lX� �H�j�5��q.Lbӣ�3��F���&�z�NA�8���b>\��t�d=0*�#���`�I��<\�Y;\3�_�謔I	�8̠)��.{F��:�"$�*�5���TX,Q|WO��x�=��X���$GK��-iǜ<*cR5r�|h��㽌qӐ�m���{���<��>���a�'k͆��P���q��R�������[��.���0�%01��H�����A!'��ś���#i[
�H���Y�ID"ن�=DB8�����kE�5ة(�k]�iY��E��x�ǜ�5�?�d��G�ǈ!�E .R����;(H����[">iOb���%�d��|�(�+��3K@S�
�`�`����?�c�8cZA]��:$��P]\�y|h	���lG���$[��H���5�"��~9��m��Ɠ�)k�tV�t�v�HR�[B2MJT�����G���� z]g�?~��>�)��*�Ul�r�;qHO�$,,�.���[`��[إ-,XH�� �BH`	!Ŏ{�%[�z����g�i���y�ygl��I��_��[�=��{��)��������"�G�����~�����;�1)�O�E{@�09�����s0���U|��_�k�}����8׆t��^(q9oN��8�� ^�(0��c�� h��x���6JP'�ֶM�3U/���p�X	���B�Wl�*��w8�V�!7;��G����AyYۿ�!�	d[��zu{�KKFKJ�&��a\d�)]�S���PKsMs"�[�r�0�q���MNO�Kz�P�~��(����B�7�8�A�X�Ql�!�� ?�AL�bo��+�9���w w�m4F�K�P��2�
�m�ֶ��/^�`BE��c>lF��C���� &�s:��u5v��g�V����/�J֩�B�0��9����RK�s�"6��@N�/��{�Sp�~��̀ ú0����L7i�@���HERY=�K/ٍ[e�ԄZ��o:A��"�N�0D��̠�nr�F�2�	���C��&$<a�:p��ax�N$Z��PߪՑ!�d�VU�|,7���m���vD�� 1JXb�Wc�R��k5���J�Z�cFJ��+z`@����z�d��+>Ya�61R�K@���vu &��կ�u5:�vcj�p#s\�c�. 3�\��
Yp���ܸ��ي�ڢ��]'"�X <��y��B9�2�z�DY�y���`c��Ș3Ϋ�"(c�V>�`�Q��?��k,��+�H���JЦ�Z�"(BN܄]T6�A�`�e�\����h�<`m�pfݽ���F�Љ�[� 0� ����ar=!,"K¤d���������d�����7==yE:'�9�k�tiE�����~��G�<h�-o~��/~c,-��_��>�׾���~��̹3ս]]�dd=���A�"7ꚩ�^$�����)#��y3��r5��T�b��"Xb�����\�p~��׹(�@�əS	��tL�3�Z�'�\�D�"��=�-^:�u{k���μx��<z�("svO��p���j�g�l��\sӲof>����O|+��eZӍ.�1|�˙1�0ׂd!FS+ߥ����ku��Ò��ޡ5���	�l�.�pb�_��`�B��� ˟������a�X#���քa�9"���xMsP�S����7$$}!��3��0�p�*|O�5��jy��t�L��by��s��II�����3*R�������ٽ_ENdsǺ��7�^A�w ���b�Gŭ*��b���v���nԼq�Y���G��1Z=z9��{HD��,�s�ؙs�8���Hq�D�CP$�(3G�?�A�@��=84��y�b� �H��7*��U�bE,�5R�S�AK�8�#<�(��w�y��q����-���?�`�b�: �g�������1�)*�=�j<q'�Q��e��rpCV�Sz�O��z���R�;�k��ʆ^�6����&eU��աAX+�g?���=�)�n��~�Hy��em��eR���O_1�@T��=c��J�A���=8��/f���c#!>� G��#��D��x���x�����w)hZ.���ZRz%�]��l�E?uM�꽍:w"�&)�gW����fD�e��LƉ\,YX�җU�o� s6�����m��:�	̓V�/�x�䳣p��u,���6#�b�|��à�-q�BlH x�_�s�qd'���ay��]!���Ex���� Q{��ά�m���"o9ym���x�x���5����ӷ�1�"�j�:O�`�CyQȡ�b��Eδ2)y�m"��J'��R�Zi7D`�S��%��&l�F(�0���-4��y�D��Hz1�>��r��|��e�:q�*<�|a���3�D' z���]��1x��I�l���/&���cyJ�5��s*Ɔ���1�1�A�<}�c��#�؟���hA�;��"��D��~��Q�1���f^I��a�Ѿ���7i��Є��J6͚;ιv�렎���;SVVq������|�CBCb�=>������4����_{���w	8�[�q��tNC�4ޙ#d��Ɯk���Jr�x�Px�$d�
nQ���E�\���R�(��:�U�S�0�ä�^���W�\�����Ar�ϙB��q�P�������kH����2y����6񩇾���8�(�7mg���3������Xu����'maN��۵���t�.d��[P��m�P� ��<X��PhkHPXc񰼡����75��P��U���O��r��9����8rY �9��D�v�ЁE͈R�{$�o>�+��9����Q��~ئ�ٛ6�X�����0��-+vvE6o;�>�N|��Y`��Ȕ� ��p�GQB�YsgV{.���Q����3f��5�#�KC�f����'��]�vj���܎��*�F__���:��q
�����8����j�����K)h�xgS]��Èž�n��07A2��Ƙ�B×`�Q��֗�^�&#��]�a�6�#�}�/����)������'d�u����hv=~�?����/��/����r��_���9�V���nH�!r�d!������}0	Wl�Kѐ~r֌DT�$" "c�k^��A����&Eu:�z𧧈"��*A�ю��B5@�����x
R@_�g�S}]��JMN�M�MX�A���&��Vm��gB��X�~W��Z�Ed��Ν;��駟��v�Ԃ�
��,���5����xoBa�d�Y�P �^X�M���H��<\ϵN&ꚽWz�k��uxٕ��X� (R 2$���9Ȗ����V& 42�����D5����.ϛ:\�\PR������
m���<��k��	C8=��c�W?V����}5K��x���Zx<1L����3`�Di=�$A���Y� ��d�cX�{��m��m)*��?�T� �ݫK�b������Vím��gz�:~#'F4�+=�bJ�8
��G��0W1#/Gn��ع��(&B�>��Hp�d_Օk^�� ,3Mͅ��,B>
]��>s��ၷ���z_~��~����ٟ�����384�c�%�o��Vù"�4�n����M�.�IOEYZ�z������1���[�D�i�emQA�f7uv��S�F�		i?j&ee�^!��M7�݈5�)���F��Պ�T/���b<+7ؘV�X5�O|���T
F�# bR���H ���P�@�|�E��t�}Omٲu��}�o�8u���fޡU�2����#t�O��F]ց�EZ˵��F01?6�����H=�4��B����n�`K�_ޗY�a!g���,<D�TE�̚N��}��nx��;\6��6� ���>T ��W^߀P5�B��<�c4�C^�n\BR8j���9��@�p�^��	@��<����F'�Q2h�d0v�������#ı�5�G%Hm�}��#
�{D�PF�K�z��<a)F��(LXE۷�� �v�F6C��p�1O���� �y����]�ه�S9pm��s���37Y�2 �x8�A/1N8�a�UE���i<K�𶮞�����~���!]��e�e�g&���ɔ���<��B��E��|��|��3?��?�u��������,)*l���t�1�f�0��N�� ��Opj ��u����&Ѓ�&6��R�:|
�V�w)�{υ�|�E�+��D��t�
���H�!:�7�)����{����Nɍ9�ʪ���}
m�;��ha�(�UWS�T�V%���%�H��Uyݨd �:������O����G����?�?/>������nY�[��"斵GDY
�t0��l����Zpʤ,�I��;]��4N�+��sy��[C�X!|�M���� �-n"���A���Â���?�$$��#�xX����n9���#�9�����G���+���8-tN��7w�y�_��� �=�緥�&�=[�ߔ~���Q������T����N��1��=Td�}���	���sT/B>�2[�ɋ�P ����kauc�Q���Y͡�ˀ������ `0�p\��˝�p���گՂ�1E+X�!#�c;�X�Hd!��F0���(�`�X��g	��2X�|(,����V:�S"~Iy<wJǦPW޸~���/)+VTf��_���Q�ڥҭV	��W��Hh��z�ȃo~�i���˿�+�~��7O�<խr����9��2BN�"4�N������j殀����k�<r�I���pM`T��b"R�-��9g5��<�ʕ+v�%�RG�#]�G��K������˰o��m�m�k^�!���*������0K��I��J�VL���b���N��J��}�\��ڦ��q���
5V��cG�u������}i�ޏ<��Ï?v�?*��� ���72�F��-%�A�s��Wh����2��x�/Bn�pJ�ּQ������0����l���ж�/x����5΄g=���<� ��m߷r��?0I��Q��� �@�����	r�f�8#=k ��Mb~�;�Z���$�Ͼ��� ��m�@v0�c�<�_Q^|P9�>�i$'r�:�Zyf1�0/����5�T���0蔮��B9>�âf���c��c�m'X�`���AE�3�)�s�U������
!�p^c�c���!'���1$0Z�\�kH�r��ZX'4�F��U�$)�Bq	c�S���s4"�yyfxpk&���>�m��z꓁�UTT���'/�������T__�SW[7T__7p��w��@�����~��~���_ڗ'���%K�<�����
6k9$�!u�I#u���ȹ��)#��v�{��e �V��J����H8�A�#1_�<����q�J�
~.*	��� 0Kw������{��ݫ�'?����'+�R.���S�6��ְn�*���逸�����y���;vq3���?��|��{/^���՝�Z_�CLީ�� �==p�!aASBk�-WB�0�YX�p�MS�t�ի� Dh
u��w]萫@m�<���4s��yA[f�V83M�-���0���E�lx9Y$�9�ؽ����@��+�B��F��
8�0FP����G+�ӱ��1(����4}��M0<��b1���F��f,x���~��h�q2��U襫�(x̤ ʭ>~ �	�y�Pq*#�G�<8��#���w�>�DV���ok#�(%L�6 `���i�K��#6"���u'ﹴ�����n��q���\VE��]�(a���輙��Z���W�����b�Vu��u��1�'�>#��:�f�f��"sE��A52�?5<40���9t�ln��emǕ_�������.in�"�J����;w�|�5�:,d?��?�����+���=5s%s�[RRX廒^��v����jnI7��@]�����=8Y4��Q�W�#�=�H��p�g�>����9����(�lc�R%\7�C��*S@��t����^}��g���_����.X�;h;���fn:j�m�B1�+ۀ&������O?����x(����w��SS�7���ҋ/�����ߩ��Nݸ�x/Ɯ/�2!���[X@�9�W̥�¾�3Xn��|u�A^��� ��Cm �{Wy�����N������1�	�N��$2ç,J��¸��[�~Ķ��=ʽ����G幅뵗�e��P��4�`	:�iQ��z�SCm�<do���#x�O<v<�~�K{�{v���I����7�6S��|��zfK�-4U�ޕ嬝&&��;��2���[��7O�V��H��;�:`N�Ĵ��Q������0ў��O�x�]�7��Nу��{��S�b��`�����ι P�#��%~�QУJ^���o�kx�|��Yz&;�A��K;��4W��J6 �ö1��#���=�]ݭ]Ǐ埐l�������]_[������xG�������l�O����C/��rI}�{=3�X�6�׬����1�
B@J%��5cr��J�e/�R>^�u��I�z��d[�N윆�� ���cxa�$��|RsT�6��T�Ǣs�݀^��&���-KϜ9y�Hiq��1
a"e��m����O��*�o<$˝�jS�@�]_��W����S��{��_]��Ï��c|�rl�L��v���"�-�h�۲����%;0̇���m���{�/��ڽf��iMϪ��jƧ\$%�x��qX}��9"��!��2�h�"x#ۡB��Ӎi���o�=s:ΐE)�u1��5�1�̸ ��׼���g�-n9�z�+�n�y�941�:�{�ʾ0X��-���+oC!�%7B��6^+� �R� �	���6��&B՞� ��@R�VZ�G�^7`��q����`1��C��ΈB����6�.�25R��+)���v���'��#9+6�1R$@�o�n�*�`�k�sb�|�t,�
��ؤŮ��7�'r���	׆mیD.*�Wu"h����
���Lϔ(=Q"äI?��x�?���?���~�ܙ���������湖e˺T��{Ϯ]W5D�k��?N���'��7U�U�ZT$��D��f���3�9�-�PFʵ���S�pJ`N9$�OdDRqµ�ơ�p��D �DR,Mb|�ǝp��|�@��*&���&B�+W�k�w
��n�o�=�Z��ce�cʙߧź�xqr�,�,�,�q��8�Lc���gΜ���㏞A��ך���?��?�����G�9�N���]߿]�U(�o��G��=�AOnd�i�a+�|��r���� �b�O�Ƌ������{2J��'��#��9��G|͘�b��7�"c�u�r���F�"d�Ǻ������T�L�y@��lب1�'���n�pMzk�˹z��Y���mT�7;��GD^�'՟��-*T�]�c��MB��R�ym�d~ �p��HS�\7���1��m�H�8u2�p�����c7�}��v�k��uww�*��yg��a����"�:���=�Y���$.򰻕Tq}�<뉛:^4�����3_	ɦb���̓7#`��n�̭oY�
���c_?�a��v�~��F朞)�<5�n�9�c23�m�=�}}�'��G~�q��mY��랻�M?x�[_�����WG'&Vj�e̾ %@ڿGRB���u7�0�P�$e����]��II�*53���L�D��յ�QII'י��8f�]m�X��]����,����fR��G.�G
�����inZ������c]��߯r��9�Ŋb������\��kv�
�����x{����s���o�`�כ��߿���{�<����~��'N�x�4ٿMa��hK+��I+I��iߒ�����n`T�9�y!lK���и=�����C٘E���&:�����H���+�)O��%�@&�\�}��颅 ����; �#�g@Λ�������Z���X��g���g駇r�޾n�0��QD<dB�t;�5���D�<�7����,����`��t@�J�BY���q8�p��497�s�9P�K�L;�n98�׼9����Iy����ԑ&�3�a���+�����e����a�8�ǐ�x�/��mV��nϚ~��[�N1̑<�rv�����y�	|yDm�P4����w89��p��.EZ�LU�˭P�y�t�<=3���O� �}����J���C�ɴ߱s��}��������s�����̕�ͧ�b�kp�1D�ޭ����/�(J"����!�Ȑ��o%hz��1h`�b���h�Q��}Y�v�i�D�?-l�=�L�E�k�7p�W�+)�_��L��O���-�]<u��3Z �)�[����o�݂v�G�7��=�w�r���[,���z��ԓ�~��<���v|�]��>����{_>~���"_�_�ۥEa�	1�z����@�a[`Л���6 �u��K�^�m���Y�Y4��/�f7,<;v[������F�3�@�\(P�,^���6" �xY�����x�[������5�N��;�ӗ�����8�F���s{� 9Mz�s��F�����>FFd��*ߋ/j�t��MhD�S�ղ����#�LG5#i1����,7�AB}36�m~��l����I|z9�O������8@qlB�'���g�Λ0/8���e�7��;�|Q�����w8/��p�WC�j?�@2tc���&>�w$6Z�R�m�7op.)/��w�����!��wl��>���������k�L7+t}���ȷ�=}��ٳ���?���ϯ^���<4��R~���\�r��ѣT��u"��ژr��k�69\�����)!3��8v)ec�#�d�6 M���Kx�He��h[�j�"^V����A�-��٠���";!7�pnY�������z�7i1��o�K�2Xֺs`3��qWV   IDATR*�%V���/�vC�$K�?��/}���/~n����dN�G~�B��?�W���Ç���Bԇ$�@a���������	8]���V���vӒ	e�ԯ��,1Oj�pȉ�4����� ��w;*	!<h¦���й��w�VM��<���y ��ɰ$�*g��a�{I��#A�r��y�|���٢GW�3-x�����c8!�����H�*�
`G/r\����#�(���^�	vOܙ�D"��Ӻf�^��f�h�C�3&���Rc�/ێ�T��12��{�*���������5F�Ӷ8�\����8Cn��J+��94���Q�uɷ�w�k��o��_d�;�:�ZqT0R�Z!��Y���Gw��&rK�$�ƨ|8b�X�D�+�1Yr�4_:\B�a(f���ڡV�LI��kUE��W$��店v��K/����G����Ukִ��q׫������a��}�jni�RT�Dt�������k���LN�0D)�l��41"��sn(͝E|������H:���P<xǯ�4����F�xAA���"Y�S@_$'�f��;n?~�����[)��J~��S �_���勹/P!g�����?�W���ȑ�/}�-�����}�?�����9x�������CC��n���9˴(K�Ɩ�,"�����T��pC�<�C_����A�P����s�C����8�/��"�<��!GϹZN��9��I�B���
[�j����;�[�|
 �Q��pf9yd 	T-[���B�qtl$���t�i�V�Q@���ͼ��cBڴ�n<7�L�N�@l?�	 �$��a����4�ըk���h�7X<]`����c] 5�c�V�6@Z��z�q ?�)e6��R$:���\�����5��6���䭔*l�j�1d�9����uΕ*�r,?U���{����g�Y������EN�]�F���K��W�7���!���ν����v�8Y�[��<�*H���m���@GG����/|��e鲎w���ف/��g��?|���ݻw�y��UTXP?"���1E6�sa��t�7-fS�ϵ�$��0)_7�0X=b�k��U��-T��G���c��)W��I+Sc��ч�ߩ�TΘ�п�	M_��f������>���^z����u_�"���U|1��les����g�U��3���Mx�Ƕ�~�ni��["�f�����{�ܹ3�W�\z��� �k�n���W���},����n�Wy� ���{��Ic1Do!�y��,0�FzX#��w7�}�w�E�~���G�+wT�����U{��?g�I�x�`��c�S�ĳ��pd�P�m�� ��� �=Q�{��K�3IO�z��<������bFWH�"���#@
�z];�q��&ؐ>��1�5y��<wo�"#�H���aV��5�ƑW�j�E���M�'x�+]�eu�/���DK�~�3j��y�F6�Ǚ"ҁ�{���FG��|�,�a����������ތ`e/`���>n3�B�a����M�Y����'����c0�'/���Mʧ@��B�����0�k������t/�����K�-{Q!��M�l�>z�X�ɓ'[�y��7�tu}���{t��
%��y��~ޤ�3S��"w�^b�G5.W#D;�%��j:Q)d~���W�'�Z���|*�C/�k>�g۫M��!�G�,��߹���5��t�I�c�γgϟ�����F-�M�<-�����`���.����R^��}�/���Ž�}q�{_���>�A�ڻ��{������ʕ��������57=�N�F�Ǌ}���a8��#���9���z� ���mo�d+\�P��y��M
o$l?k��d��������yoc�u��
c���G4�8+X4(�Fܴ�9�p��6�'��#�����ڀQ������!��$ŀ?ȯ��t�(?QR��GH�E�J1X���w)M�'�m��,��a��-� ��(1C�yB���w�Z7:ym>ۑ���Ĩ�X�6���NO�ȉK�P!Zs�0¹ ���p[�|��-��]�La����ES�b��:�r7��������y05-��ɊDLO���y�$�Je��/J۵/�\�f�}K]�׍?��h�>�{�7�Wt���<�Ɉ�666��S'O�t����|�/�?��SK�Z[�4<8�K�+Ľȅ�aMrt�*V.�Т9.�ʵ��l�y�vP~M`G#;�Z�\��N$�4�M���v�l;{�������Yt����_xO-��S@_g�&ú5�'�����'�x��ߡ���eB��rpq���8����q,u����������|�/���ww}#Ӻcǝ �e��_|�й��O�>�Ez��)u�]ZV��ۢ�����57 ��3�����O��=x���:���Ogb���k\p����B\�"���h�~��uB���y?3C��IC�jV�����=�o��hޛG��Ӏ�	�y^�uё�dq��ow |!a�d2��f ��E��l��|%'<�@��Zc���7�(���^Qg6	���k���l�N�0P��d��aa�ӄ�1��Zh����C9]L�0.#���R�I��i$�&�	����;z���&��׊��y�v�
��.�pysc�+��\ٮp�A���2��"���,l6P=2��w�wc0D���+�$��#	\.���n��Ӆ�ŅKe�-՜����9��Sub���4����$�����S	����߼�c��qރ��\s�-J��L1�!e@��2r+WF�>o�'a��n���n�z�(gB�謮iX���|\�)�_�������w����������S�7h=�1#y��X\ 	�Q'�`��=֗�Oz���~�����[��?�;������73�w���8��c�>v��-��m? o����{.D9{�0{yĽ��@� �WF��R��vD�g�X�
��zJ�p�7n|��%'���|f�"�Ƒ��<]� �g��y$�礻��\cK�;3������&<���������rwP�e���Ѣ��0�B�CJþ"6���`ю�R~��t[��N5t�U���i];������7,���Ғ2um+S)�ۼ��t��^㬚�@��!\#�F0�`:o�F.A,a��.-|���Z��~8�'%���g�n0L��**0B�%^f;���wff�����`�	�@�\pF����ql>"���YuN�@��Q��nLr]_�x�X1��./-N�*˓g�X7d�;.��� ���h��.L�/P�! nO�8�n\eG�ߧ�k[VE�Ss�1����S�I� >_a��\2&��k�^>�o�_)���s��q�������?����$yi�{qOy�Њq,�ֹ�(m]����-F-��#���/~y�o��_��w����7n���ί�L��o��������j6J^�{��߯n�<�R�
�_��u��O�o�`#K[��,�ءX�����jp�����m+zKN����t�e�?��"!,�O]���y���Yy�<�l�����Z�\3wl&=WknZ]��yB�o�ռ��>\�a��+�?��ޜ�=)�W^�wz]Cr���2�y �/`T��V'LT�vb<�\Z;��˗/�&��9pA�1�?�H��=q<B*0<��;��2��9�1}�ٵ�y������O}�1�w5Vg4pI9��L?�
���*ߏi7�i�{���������{�#��|�h��E5���7#�l�~]D���o����2�8�"����\������2Sq+�:a1�.BZuu��.V'/^T�a���[)e �M�I�k�ϗ�e���w\�p���	!�v�U�DF���El8V��,�0.0�گ�gPBF}~B�#��u>n��lۺc�������f�H?�E���E>K�ᆴ�\��&d+��b�CD����={�4�����G��~�;:����]�3`��/9p��+�/���PHu3JtƂ6��C{4�}�uB�{k>�.f����^sۂQ��_XDM`����<��>�d��^"�G��Mc�1:x��k�n��_�au�@a�-���Ǔ!�{�Ga �r�ћ�9g[�-б)�v������#�i�&�#߈���� V/�s#�	v.�ST��0�{�=kG��6ў��s�;LJ�;��i��LF�W�aG8� "��3p��q��*J��q��Ϲa��|a��t'N���+��iJ���=V��s�8��w�߷���3�MF�
@eD0o��K�87�"7a�=��	ׄ���x�F#�K}�~�]� �|�H�U�**Bfepr�8��Rt��H���X���L9bZ�Fv�)�y��h�G4��9��P\L0�7BuC�k�q��dV?I��0�#3���OO��7��Zkjk���b�=��r&n�q����z哟��ﾴo��B�/��-�($8B���eE�"Ѳ}�âc�Lnnaqn�]ʧ.��O�-��{��oy��m�p�U)5y�[ޅ�޷�現���<}��}����wjqi��J��9��ZXŔ�Bw��k֊Gl��:8�B�y�4g�8�]
���q�vÅd��	�{*��C_��Ӯh�$  ­����R��x�x�E�#�1<X��V����a��6D5K��Y�7�u�v��G�ZU�i��4��g�C�#�%���qfy����Ng�����og��>�9����TJc���tT��xo{��+��P�J�<4�f3R S{R��ǘQ4ʤf�}h.��.�qt�=�=ftU����sT+X��߀��ͺP)R4Sc������.<W�mz_�9�;�q�V���x�f)w�Ȋ���L�<�> ���H7v�s�pF�E�.J���T�r��?>9w��y�uv�@sμa����y��G0�����.��\�����m]kF���9�$�c8_UU����_tW�Я�\�[�&f����N�����o�=s�^�Nʻɝ�ql֖��|��Ͻ�m�?���"����a�e����|��g6�<u����o>����]�&������n�������>��#�-!�=�"�i��* oԂZd�f���å�0♯Hv�v����D��=[�,����䚗�`E��y�fXx���o�6��}<pcD���L9�&9W��1lo�r�`9.v����0�JC�~�΂滀?�h� ��
S`�7�Q��J���;��;��
���`����{����>���� r����z�h�`�y�x:�ɠH������}շ9��9�� � �T�d�wQ)�>G�=�&5s�p.�gK�^�<T@^���CZ%�i��0z���$���/S�P�UT�^�䕭�܁�b���Ĥlɛ
�En�Ѣ��6>�*��H�s�3�'���fg,�t`��k�R&�[�� �sr�\��
�[$"���`<����ֶ˚[�s��Y���\q38�賏�����`�Ղ�sƭB���2��e��c�A���UHS[��k'D%t}���/+-M=�J���3�5f��80<4�
c׈!}�����K[���Z��{�X|���nN��}���%�h��>������z�C��ַ^Ubˇ>��,���?v�Iu�K{��ߣ�ޝ�M:�
��q
^�U�8? �L���F�
�lp�ڗ�����������ӣV:�{_�e�rhM? [è���+H̟P7��h�=�%, `�� |c�.Ԉ��r��#Lo>Ԥ��u
��x�f�lIQ7�¢m��i �wA���iO�7���b���~+K,u�xL�#"��X  �ov�ވI��5k��o�7{�r���� ;v��͙4�Zw����:��%�#��)��3�Y)�� 	�4��[^����>�`/+��G"�h����jr��|�-S���V4�1���D>�#���T��R���CU�O�Z�j���Q�p]�+��B�)�ҢZ"���E%�����F����ι8����&������\��@�nXs$�k|�h0�eֽq��_�HbI���Y��4B��A:�G�W�*��7z�O=�7z���}�ض���^����}��% �y��o����&���lCF:����`/[x�'�7���I�ɷ�=sj����_��?��M��}��<p5O��[�McZ����s�/�?�p������<nT�� G��r�(���7B���<��N�!��vR�h�����Y(�ј��~��|E�^�7n9dm�R�ˍ�h�H؆���F��M�.�z�R��V^�OR�����׌Ǯi0��%���:	��إw"4^?�^b�!������V��ܐyv�T��W�����X�����hqq��e�ĺd�脭!�q@\o�a�i�H�͚��ׯ������f����+@imr�ԭ�>�Ԩ�F/ϒ��g�f~�5\�}+W��:c�wvj�~l���C�{V :3��R��p|>��~���6#�{�m���x� ���i׏O��e�v�� �\�;����[������`L����v`�G�E$oZ�A���'�|6H+�C�+�q��x��m�OΝ?�\��CZ��J4و�D>GԲ�'��9�Ԗ�,�����5#j.��M�7���$�����mWs����J�j�f��oz�����}���S��Q7�Z#~�Ǵ���{��9p�͚{�ӬVT�����=r���'����_��?�u�so}��7y�Fl��;t{xz��/W_�t��������k�Jtv����\�Q���J��ټy	�º�y�x����G6t0��c�ü�g>�쑀H�h@��	k~���y�"9kF��|���"�ѡ�И�5�r6ʔ �Q��9a^��:'��eT�[�x-ge��3M5�B:�� �"W�mf�^g�;B�?k�	����17x��姼_:�s�P�z��~vvx����ӗԋ\g�~dk�\��U��ꭧ�K����|X�u�9oyxg�yO�  1�.�m'=@�>��Ѝ�ro�q�Ok������Q�K��Ȋn,���]����I;�A�E�p�	�S&(D� C!�W�7tyyCH�Xĉk(_1��˵1��%��8;>2����<�L�$�Q)#��}/Z�HD^�����m�m=�����ukG]c�ό
�x��[�zFF������ot=x�����=���_���-�?��>���Oe�{z���b��x[�c�+[� ;hw]mc�1p
q2n�����Ub9P�!�Z� e�J�n9v���'�����|j�Ν'���?xU�_��z�;Yx^���'�z��;��*U�S�7�נ0�m���m�~�ˋ_:1=]+ŭry��u1W�,��yS}��<<���C(4d䳹r[��jnS�k'5Yd�<x�\:ԭ%P�Z#�x<W����-�/#��-�$,l�N��
^+����I���V���D�Y�#i�|';Σ��C�ׁ{w�!,=.O�1E�7�`E���+�P`^_�`��q�*�k��{ C����G�c�?osp`H��7���gD�:ɛ
l*�1���V���чI��<9�wKs�I��}~�0!�!�`�Sj�*�[a@���.�KF�Cu#(�W�䕭ŨE= ������<���e�i�kZ�c�s��-�@u� ���j{�S���o1��X�vp�\t8�o"ܬ�;��w�y����"3�Uἃ��v��:��H�:��g�M$k�L/�w��p�����|^��i�b��)�w�$J�b7���.�=,��KK���E��B
�o�D��ym3�-oW�c�~�sO<�����Y7�-ʺ?Y^ATad�C���@8#�;@�ʚ�
X` �i�X�Ȼ�U7����o��h{�?�Կ�����=�}۶�]w�7��F��>����\�/����<���Ry�%�}�eZ����v��Sr��F�w��l�JXW��*S�{��D�q��^�Lm�Ze:��i�,��?��̙�1�ҼL��U�V�AyU�E%%c�����0���N���������ZCH:����*�-�XUK�5-���zQp�}�#��Wi���!uV_�A�cARG7޽{��Z�Ի�9s>ֹ��*����-�tE J9��P�Lda�]T���ƚ6�sV��U.Esm��cBr��%(P�U���'���N�UK�
[��؞B�!�O����MI��	p���_��Y��v�ftyD�y!�j劤O�������x�%ʟ;^��5��֣� ȅ�;s���"�xY�t�N�o6�5�MmL�GQ�x@�@�����B�� ��cDk�e�8Y���-� �@�9���0��]����<c�&�;�	��/]_jUKuxsCQ�6*�\k��G�0V wxV�RF\k��>��-(�Ϛ��j��.T�.Y�|�I��U'F�^�*�~:��7h�~�Ѳ�y�ΎΟ��z���T�+�������o�]P��I����G�,x)!����3�j�S@5+�M��9!&�n��߲��s6l��y�=���*����ɱ"�~�D6� �I�r���Ԥuց1Y�B�̛3�EW��\	�̙���2r��Y8%�q\����M[�b:v�"E�?��8 �9v��]��=-l�Y�<��b�ɕ�X�y�<D�n�yhhR���=+��D�,��fi�C��c���M���qY�Z��6�y}fDa�'N$'O�2�|l$�bg�f���9Y���Q�~�0���E��$-.�֝n����?<z�h 2ƀ�,���5��L�č��
r�$g�jj�5/�<!�=�#b��7J��Io;�9)���Wl��lp�L�^�����?����ͽ*�=Sk#�o�z��� �
��P'	���><p1�*u<555�.s�P3V��y�~a��8�(?Cz�T���Ѕ��|~�H�w���h���\�	y�O�V�dģ)e�c]��J����:� "�����'�B4)�!�M=�;@t�SR2&�v׮�l��;�Z���^FS@��3�n�����O��+_�)���45=�-
E��QA̺0R5)RJ��������bg��*����	PWC����ia��h[紝�'�[Zlܰ��-}�V�W�������t���7���omoo�E��-hu�FE�՜	OkM�j���I�Z��0�/����lyrL���27�Y·�m��h ] '�&XCi�<H-�D�Cw ��λ)�i�nkoO�J������X�����׭]�475eC������(���,��6���$()�����WZ[�3$.@%�č����� Q�Z���%�x�J� �A�ՑA���̸��c�~�������gƼ�jy��#���B �2</��!7�cD�|od��@�J?���[�;�eϸ�/�㵵5��#a^���\���Da~�%�̭�ү�8^g�Ƕ��޻\Q!�+�14�դ)iWJ� �\*��2z��&"�����80��1(I#uwwZ�$��֚�����I��������,[�(���4���/����������~J���Ʈ����B�c1���}���C�,�[��o�� cn�� t{��(�EN��̀,�6�ђ���-K�>�b���C��y����]�o�X*>s���gϭ������]��V(ۤymԱ���0W�5c�U�΀��=u�6^g�u����/o�'�y5BdF�ջ�k(��i#o�7����g,|$�Cc�kN���9%��z�j�]î�04���X<^I������2�� b9W�"�`�wW&�p�p颕��"&�OH���DF�Q�s�h�k�:n0 ��y�����'�9��}�2N3� s�����2�'^~̓s�U��v��;����w�D�?3��E� 9㛄ȇu�#2����ݢb9�؇ܔߔn�����^!2_������^q�:�knt;s�5�R�Y����xTC>��z�r�Dz�c8u┄y�����~��0DO��C���vR�LG� ��!J`����k֮�����={����O�9�z��O,������������+bY�i��3O]K4V�1^!Ņ.Jk��p��t�0�}���DiLSڒ�K'D�h<X�uzrX[���+��ey����<�p^����K�o����5��ZO��{�)lmo���h��lk_��׷Y�q����:��[4K���S��a�����y	�	��R&�����HN4(�m+�/wr�@P��gދa՘;�"/Q�=��0ʠ����I��Mթӧ�:�G03q�@tbE��_�.mI��\n�+1�j}̍�Eh��pB6��0r�oB�mOI����Z��z�>�2��xR^�κ�$���"�5����w��<C�� !F�:(��G7l}��0*��	�
T/Xw2�̻�@��=��F 	��?#ɉ��������v6g!��缳܄�����32j�\ ���L�	ۯ�B^SS���+���1�k>���-����� ��آ����1���>�< ��s*k�ć� S�_g{��t�y��N� �L%��5���o=��:1c�'\�Z�+C��a8)���{��'�l��ˢ}���hOM:��7���'��߷���?"ڡ:�B�D*cE=��9t[(����_<|9����� �`�а`��xR-������,hZ�GF��vmC7}������UUV��(5Q_W?�E{B!�э�6�.�����D2�%Z�K�:���{� a����6���P,���^�<a�̠2�}E���"�zxz.�{�Cr���9�3�䧈�x��5�l���Fh2��k��DB%VL3`�e�f�����'��j.��h�W%���p��'�z�C�ޮʭ
���ĖEO���TN���I5�0���	�s�ޜ_'C�qcй��(�y�z��d3/�r�U"9�}9&�·U��N��&Z���f��[�r:������F%������\4�:�C*C!mhp(���"�C^�Nc�Q��"�v��N�?�b��#�Q���L8&�Y3����6�U �T5`����9��=�3��T*�^��]+:�DmH��ёxx�Y��ad���5�sS�f�9�(0ކݣ��\��Q�?��S"4����d�W�1�����F��4��:���'�k���ˠ��s�����3����?mnZ���h��ȑ��u7��~����J�W+�w4�b�4�d��\5 h�ٞ�=u�qbB4�D-4O]�I�:��1G-huS�c����%��D�@�2����k���_[�B3����⢒�ZH;��mZ�z5�	��hA�{wJb'-r3Z�f"J�	0`Ҿr��ܱ��B�[����g���x�<�FI�.�B\+ϱ^㮖GU��.(*(�
]&9f�Uk��,��it}����â�u�	Iǚ�p�,�EA 3~�!m�+�s�*��"�R�tdJ@�E�}BH�Ղ�/e.m��xB$�/,_����5k:nݼ�D�?�����K_��-ޛTvv���/ӷ�th͞��֧r�rՒo���^/#�������f=(�i��F&؉ ;������Di�.G����މM ��4J�h�*Ic�e *p�a�[)^�X��`D� O$va�7�ع�,�M��I�^ۍ1����gL�t@Όj�-�cr�\����͸y�� ��h���7 wi^�.X~��������-���4W�'/<xX�U�[`�x�?��������^���v��Ε�c�Zx}�P=) ��(��s�� hS��k;x��6ל5�	��]�9E��8��e.�ޞ���;���7����žP��b?C���������Jy��/�?�l�g�7�0�a��yP_������)���p ��,��gq�<�i�������S�2����	I/.�sx�S/mLi>Xiu�B)�g�x�>��.3�Ѩ�,����[S��u��r�y�{-� �)�˝+���Q��B}��B=��P�Y=��Wx��p�K�k�#a��f-���c�4F
��mG>�l��o;����c���6-4���>_�� V����0c�]����ꏉ���5�;����c���G��	_&�@A��91�'V�X1�HE���>�Fu�?����Vǀ��M�`d�\��~�{�ǿ̣����`'�Ã ��n�'򶔓�ק0��sg��fy`�:�h�������;ax��^#p����92Ҝ���ayݑ����R��A�[��#'.nc���GDރHc� ��촫���F�y������g�r�����������zɇ2B�u�'��7�l��Ed�[Jܢ@��T�*1M
6�����;�C)�n�{˫7���PҨV���]�R}�]�ߥtF��!�|��k�4���d\�҃o}�����t��~�����O:�W1O>�D��O<q���~B��O��D��!_Vl�hP�fL���C>ј�ZU���=߳��	aybқ�"/lд��.�[
��^���f̻Ѣ)R����Z`�Bx��o�ﲣ���4��f@����KhmgpF0��5�����}��$d6��d�Mȃ���w�-H��4f���{$��x0�0��g,t�㋤.몆4,�N�(ɗ(��?=;uFcث��/�^���ڵk;7�����'~���[N�>��t�\[�� ��	ss�ܡ<b���9���X�(F�;��׫�&3�]@��B���[�F.X� :�B���<O�5���7e��1��ɑ��a�cD�ʜUi���9��^�F�Z�2;<|�K�9�� �)Os;�����K���� ����ucFD(�и�F��x��GT���F]��zy��M�Ͳ��\I�")�w>`���������͌"�,ʦ�Q��#���0~4�sbBb���0�
~zm��ٶuۏ�{߃�^�Rt�?��5?� ����_��J�2���^�6���/��+�L-�+��,� 7j$� �j��ñQ'�� |,h��@�
y���uAc{� 
`aPc㥇:g[ؼ����w�W�\�N��Y$������y,�ѻ���vsA(� e!pF��mF�焍�gVCܖ<l�6�0/��� E��w�u��R1`%e�a�y�����3lӟ�D{�y��'W�Z�qϮ{���u�p;��?Y��}?(���ծG�9['��.�j�;�w�;�o��gM��4x�V�E!�1T9�Ig��>/\H:�:̃e�.rS��\@g���6x����� �v�TU�<w�<����8� o��z���Ґ��
2�v��:�?\;f�"e+�t��F^/�_0�0Hݺ8?Mm.H[)yu[c���<����D��#Pd:�Qߝ��ڳ��șKWX�9�ߩ�7�O�X��\��m�g���`�H�BsL���ι���_z�Co���e+�����;��c�H�y�f�𑗊�y�[N�<�o�� z�c5@1x
O����bHZ�(�FB���ֶc��(��wොc4�k��~���0������1�l@�v�f��1C;��������9y_��mnƅ���v�tf�#V�V;Z��h ;��zt���0�"�śL+yq�R?#h�|���6��-z�;  .ڦR
s��9�p��U�_Y�j�y�u�Y�.40�.�ǟx���{������W牜{8��3\U�G4V��`n�Zs�A�ח眭�F��嬥��|.��L�� v�r��b�C��ܙ��&h݇�)3� q�'Mk��-�.��u�5�|�ܸ/�<�q;"k�3�n�z�s�����m-׶��3� �h��".n��u�5��Y;ny�L������׉�r�,:A��y���+My�{��d/4�
��D��r��>ce��'�Q�}P��f����%A&#	"���c�/ ��*d ���*=��;�������w5^�-��~u�3��"��ݻ��ٳ��[Ο?����=�eiN9ejF���8[�7X�x���x�F���:ؑw��>��9�$XԽ�
�k^��{��������vHl�������^}6�Hg,�'lˈ�� n�����Sw���6�@^3Q�({Z�D0�K�eoa��a��������n��BϨxYng^�k�;�+c�r�/('���KO,_��{��-�D��w?�?oY��Ex�r�M1z1_)�q;�P�T�q�Ir�p���M`�B!L�a�쬁Ȅ��	�*GN�F9q����p|��Zɛ �o��P"s�#�M��'a���w�"/Noy��	����<�G���^q��y5�B3����CU�,��n���s'�GN]�:FdAc�[�x(�3�������˙&У"*�@T�rI"AǮK�G�z͓�@Ծ6*z� /	䜙����r�M�O�+&wn�3�8fg./ij���>�����o|�4-�U�#�E{jҁ]�x��G���߿�ҥ��?11v�©+�n���9U��ⱛ�����P����k���=��u�,�k�KG���c	e����1b��d��f��B�C�|������e��>'����F�ˆU���>��{�?!X۷������s��r�&�<U�ae��A��Rk�����0�	�
���k������p���˗��cǮ��q~��m|�/�|�={�C@��
�n���T�Il��0n9se�#,q�������1L�e�QL�eC\��4�C�� ��5�Cpww�i<Xw��n4.�4�и�;�����ܻ~�\s�Q5�j~X�"��.l��We&�f����`^�1���:'�3���K֖m���*yJ��6z���Or6�?	a�o��Jd�����Rv�{TT��;���nw�(r�0)sHx{5v�:�%���T�T12F)�}�������a5U�G�:!��n?�H��q�FF���	W'�A{���N����S�a�J�Z���?o��W�V�wy}��cWU���2�=��P� e��d%,���I+J�����7\L��'�uoT�ۑ����zx_8�K(�~%1<�#;���.���T[.=�X˺kVl.aj��>=	���i	�!x�����yk�w�*G8�5?� ������������v_@2���g�F�~�k�<j��]@��l^�1����=������i{��-`��*���<;�X��y�E�� ����6�Ғ�8V	�)l�98k7?�Ic.;����y�Շ���)���(k�6F�[���ʶ��a���* >�4Xi�L�BR�؁{I�*j�,�N���ަt�6�d0^toe	a���@��YPn ����./�=��jӄ��aׯh
�H��c�.N���<vn�.UX~P�ٚ.�5Q��d��J�t��0���cI@��=G}+��¶�o}����@M��n�bd���|ƒQ�y�|���
���&TEߛ["RxT�k�.�s=��,� �R=U�_�
v��7�i}7?OQ��4ov�Y�����hG��]�Nb�x��t���?(�%l[/7�d�ɇ/�����-�;jW���-��Ov
i�����Ř��i�b��(4䯟Lue��]��A�۔Q���㟽I�r;]?k����m�l�}.�),��X�)�_}"�����~���-�&�h��kpm>ߩ����^�/s� ��21d9�ҟ���l5E�e)�&�٪P�9��!24��'F�Nv���k�}>m�r�MmP�B� S*�v�P^�,A�U�Qiw����|dXK��,#�Ⲓ���?��w仇��'�u̺��*,��%]&�q:�wk �ע�'�<�+�/׬*��i�n���w8�5}2���C�w̖q=g2�����s|�:�U����m'�_w��4�9����w���W�R+���ݹD�2�1�fd�����"��!��J�������0^',}�t]d�,��
?Sۗ�����B��h'���g�1l�B�|߂��z��g&Rr!;D`�Nys��9������V��[{$�j��J�	B�ȶe���
_)�W���J��.y\�~|���@�����a�j 5Ky�S�
/�P�+��^�$�ن���Յv�u�� ��N!R�3����|Ӿ7�a�B8�Pm�X����n�)�p@�{ׂ$/�!�͵3�!*��]�F{d�p8�C� �Ӭ#|z�Q������*��	�q�U����P%���4 su�Ԡ�Q����{�-��:ʃ�'�mɛ-��$���^�'�������(���R�n!�*�& ���/�NP��[��%���=��0�3�߃�5Qћ��O|O��O�ԕMe�1�k݉�Z�uv����`��l�/
j8�(̦��0��l�o^.b�0%y�˲W�\jꚝ,w�䌽v���3*�]�ѩ�&�tC����[!�2��ڼ=��б@�I&ZЇ3�� s��n��&�I� �ʁ�w�/��!��]��P��/���� �
Kc�+'��Ff��<祛̞����7�t?)��+�ɎEi|��"�ӌ|?;_�~G��bJ>${:���6�>�����x���mV�5���8<%c�xm"�2�h��xx03��n�U���S��/=�<�8�k��fEe��mJ���Bp��R�i�qV-��f��t5P7�L ���j��-a�R��ѫ>��!_L�kB�q-s�`��n4���(��F��WL�������f���A�a�@�����k���t�@��?1��]rb�m�z�d�m]��'�d�P�c.�r������]^���O�Vڷ�m����N�y�uz�[o��=)����A�����ciT����Ħ.	C�6 �
Z������bLw��v��\�d��Mc�%`�<�Bl�E�a+3�����R��{�pˉ�%V��V�?��	*և��F�o;6�ȶqЙ�p���a6�u%�y��QmK�n�O�w�Jⵑ�(F���}n��r�R����Ɏn?��1Ry�b|%��yKFũ�C��}��i��Ipk���*��X�]T����]{G�)d�Ѷ�u�H�ȅ��*�gSlڑn��(�d�C��H�����QʗI�<{�g��<qK?�uɘ�_ ��û`� z�_�[y�J},��ji*OBIkn������vb���W�`~O���ZV�?.Q�K��f�}K��o�G��e4U�W���� 8C�)L̬�m���RK�O3�t%/vV��#J��*"/:�}�v,� �����t|�tZ�B�4�g��<-\�h>��76�BLS�x��v�)}o�0�/�nO�w����©��#��GW�<T�	��PySDF��흉�@eqv�:��,$#]�0S��������MKKC9���w#?7e����d��=�z�;�Ѧ/����78�-�e;�iW��*�r�P��9�^���Q�S�SQ�8f>_�}q��|����:@��k�p< �$[�ҟz���y�Ј8��L���_2��y�����}Tnd���N�H/#\�T��[��U��<-dx3JfA.C������a�a�}�Cl��	3��R�z��/���8�7��B��sv>;{;%�h���a�3R�O��؄�~�c)㿤4�-R;U���O��U�<�ezîc��%w�{�s:����Qo:Tֻ�Ҡ���YY'�q��\-�T��z��6����FLl#Q��d��Q1h��si	ٸ�*���������Pt�w��_�a��/��bOѮ����Yb���A'��א �ö��uW�@w��yyݓ��(�\,Dje��c��F�]�*B�-�����~��3
|�0�����^�9dS���
_�wЊPr��n-��=r/	�TR>���J-�X쩹�NEcz���\�rP�y�E��ܗɚc��?�!.�j-I����c�@`O�����~�{��Nn���o(�c)'����ǞCX>��E[+\�f%�(�`��"A`OP2����k?�P
WE0��qA���L��Đ��6���q��k�䚄繓�й�I�>gu+Rx�:�y�k�,emm-��m�0ӹ�fx!���G���m֭O+�:�$�X'�\���=��ol8}\ߥe�;�����;�k���.^���1-\qq�B�v⩀����������ȵ�oC��'=������V��sde�$����M"��/���|���Xyw���?�;���C�l
��T�@@�n.�	�@GOL�UL��[�T����.�\�����4U^TUx�J�P[�GB���B�?�Nk��w��q�p��j��e,��w�mCTC_�X�ڥf��l�IGG�k���mZ��a��V��f>�t���V��͸�#�B���}zOW��3�
�0}N�pR�&�#�]��]�<�Hc�7��]�2+zO��a��k{�O_S�Sq�2��k	�������H�����LM�Z�s�P��5%+�>�H�8�G$�:0�?�G����7�\R���s��.F5�,��&31K�Pd����q3Խ����b-�Y����m$���Ŭ$W��jr���g�h�U���՗�]������Vm��Kc����gTD�����P�dϛ �v�w��
�uY�Î�e�\SI;�G����H	���*�H�5�꺇�����y_��J�XO�%F�d�񾋺=���O`6lƒO#���E���B�	�Q��������7;��˗+/Ma?��0����;��.55w���$MfUr��	�*!lc �_�l�j�gXEEBm�2�-L��L[&��	�KFt=�Պ̅5�����,�$�W(��Y$!&~�u\UWSw�h&p����p�c�מ���77�����̘	�R��]����h{�|��Y�e*�>~Y��)W˿���7�FS}�� �+E�w*�x1�	���S'���q�{����p�3X�F�H�*��F:^oe�2�\/"p�_��g�Ex�U�AT	o�6�[-!��I��p!��a���t���b���c�$�r��_
���`��\���$�1hmH8 ��rɍ��&~�K��vjvC��M����۞Vӧ6E8���¬�~1�
��.�K�;��(oe����h~ F����p|�� �'�(�)mN���{nv�ӌZ2b�����x�[��و;������m�*C�0r�]� >^�i����E�U=�� '�9O�TT1�ohg� b��S߃?+�%�j>��ƣ#�=:4�_`b��xE��GAQ���:��Q'�h14~�)6��OzO�c7'b�\S�ŸŬ��2Ŝ^gкNi�����r����T ��7 ���(ҙ!�e�0�-�B���c�}t*��Ϡc��y6Z�%��S}�&�s��qFM{�Γ�v�7I�K��k������\��?��!
��}���C>[;�Q���DED�	��L�E�2���~�����]�n����W���s $���1��=%�t����ɨ�򱸛5���W)����hB:�?��u*���v�3N�°T���_�L
��F�L��Ɋ�~2��G���;�]�<&޳-t���7��_�z^>����/{�sR������#ws'L�/�~��0�l����C�Y�8l���>�4uԝ�?f��}�~j�_��i~}��l�[�"H?��̟���"=�����ì٧.䔃�\�i!L|¾-��Q���g������p��e5�W++�g'�}��"��+��J�oD� ��G�K�2CR�[�qO~!)~�j�ʂ��|k�#��a"%q|g=~���Z@�քTq�@h���]��G~E�G�P��jМ��W6��w���Z�J+�2�A}_�BFb�Ŧ$M��5-��M����``����wX�r������(�}\c*��D7>ߜ+˗�yHy��W�<���%a�e�1��"��-�~c/�h������o�T�L^HG�cV:�!o�-������`�I�fyγ��]�92�-�O���9�@}�S���1�ЭT���7�\����c}dw#D��I�s�$�$��z��Y�$�t�LN��Ƚ��-�l�s����*8��I�kA�[;��{�A^?��,�7�d¸e����%�����yz�F ���. ����D}��ܺ/g?����G�w6�{���/�ߺ�րH9Ŕ=�H���o��P�쭐 �Q�k�|����I�;3l�|�G=��Sq��������y�y�$M��r���D���
�<�*��.3��G#�߶̶+X�j�� ���	u?�� ��H;���u��_Ĭ�Ċ�({כ��6��4�E80l�ŀ���Q����ҿ�V/���[ �Ètǂ�s�å���(�<�9Eu:�>w��d	����VDX͈��s'9f0eyM l���L���T��{�����Y�wK�"NG�0Q%��n��tb��v�ڦ�m�7?su#���CA�}�r��T������8+�������k��I�����E|^����6]]��g��w��8��|#T�_<�r�$���P����-�63A�K��ڴW^�'-����p铼O�`TR�~�O$��P����DՕN5�\��o�%�v)nb�M���#���Ϧ��ݫ�X�
H:�Ġ�/��<��޳��2��2Q|�_�ƍ�=-�=��75�����br_s�G�v����F��@>Ω����-K��;#�4�S���݄G('~k2��la~
q\j|�7��|�xW�S �� N�kg]�>�7'��O�5��A�1�L��^�,��|��
�vFB�MK�Y�ы�,	/���;�d��!m>���>��è!����X-&�iY�4QoEjk�1Q]TJSq���+0��z6�QgQ���p�Y����8#��n����
����f�ߗ@l%����	�ɮ�����mW���\3k~@l�>��"�w4;��	n���Л��|׊�GV�M�`u��u��p�!:7���kbI��&��k���|�u��w��΄h��E�#�2`w{�o꯯����@YeB��
����9��`�%@��>��� ������Sp���0ꊵ/���0_w_2��-��J<N����J�Rg�>ŉ�Q�c�
ቁ��Nz#vފW��N�����D�A�Q]�����Z'-�;���7���Kh%'�?l~�����``,{�K�'��x��uS���0],r���jh����_(�m�
�G���C�����c.5o#Nt����q�"�3��?�c��.@T���&qDy�q~-�ϕh����8;E���0���zdE|����0��8
�)�Z$�D/�V�/4��{��+��E����!����Nq2Qd����~���J,���I;��b.㐒=���vm���l�X�d>��Ƶ���'����wG*�ȧ��^#�oӫS�� �堯�.1�<<�];K�G�ѧw��0��ѧ�L���S��U����=r�u��˾j����#������5��d�j�&���eǞ�1�2�,��F�Z��w\/-y�g�G�P���}#""D
�Ώ/t�����j��ʄ!�<�_�Ĺ��!�Bp�b�Q_���~���g.m�w"*�X����M��m�����8ᩨ��O�V�O���$�z����˅,$�Z����·#��HG�~���$��\j��������2o�)Բ�/��e�]G��_V�_�P�VF/j#`7��,��;h�����VL����L�J��40t��mee@@���t�l>��xjj�̱"Y���l�_ �L��U�����@D5^4�|7X�e=W�N�{��*�l4����'cz�g��պ����'��g5�Y��8����'�(� h�-l�8��5ch��'��-�x�O�u���m�ߞqtD�\�� ��'�	�,^��/�᧌#8Tѧ(,�vKv�@B�YI�ަ��ê�����d�e$ŗ��X�����LG���M��������W5U\���Q-�8���!���T��i�M��1�
L~|S���I���f����Y{&�>�����;�Ѽ:��Ͽ�)z+|�~�c��J�P��j|[��#�=�����)�B_����s�M]�a*�#��^nb����@�2�C�5� ��B<1J�	b��4מ_悙���ÃwW$��h]u�7���g�z��A�>c�=���"�k�t3"Z�"%�����J@�)�l��k��c�ZoY�l�����3���cG}U���������TO�!F&�)�y.����e9�y���9���^.�!��֋]U���?V�o��l��'m��K����2!��
�Q�Ubb�&�����D)o�l3�2��w�d�lG��8��.��f��D&[��9л�� �*���:����+3�oKH>�B��YM�c����M��,�8�}t����T��﨔���L�_ùY��xSj����p�[�vZ�>�:�k2`.ބ��
_FZ"
s��Q�i(3�y?��?��m �l���RSU�S��`���>���_K��̃}��ɱ,�� b�%摯��BlOD�a��z�y>��*̷,<=��|ٞж �'�L%}<L�����,Zxu�H�Ay�0��*b�~@�#��MR���W�FV�N.�d�����s��N��a�C��x���_	���T�󿹼����=~�0z<Ѱ[�Q�����x,x
<#����~^�nVZ����^�?B=dP��ÓߝS�K������Oa��~$��ϙ����|+�Mg�V&P���;���1
A�-gh������Zk/����X�ZV׷4�X;Б-z����B��s��9��\8g[�]۵XRv����2���{��	�]�8��W��/�_�g��F��>���D��ᐮ�2˨�Zj�#�6�0?ip�p�Uh���`�Q`G6{W��_�jW�^�y�߆�h��Ĝ̷\�����z� ����:�K��%�̾hY���!���߼���Z�~[o>;��.u�ִ��*	_͙kM9��omW��������gA$�����Օxk�\FҲ��F�n�2є��t�p;�m��i�?�	큂�MEl����_~��	��h<v�����tu`y���Et�Ĵ	���L���Sn�rP(e�P��|�_a�ǕKI%~���v��c��Z�ߔ��?�B(�z���T�8Q�;_5�sOc䀥���f����씈Du`��pR��v��>��ˣ�Ӽ�>$������*�Qp�~ۉ�d����a�`�x����榥��!#l���'R��9`Oa��7覀��KWhX
ָDs�Y-"w\Yo�-�t'W?���{/�g��H�d�����e_05�^��/a����m'u|���i'��|�"�����iy�Ӟ潪_i�:�x�d,�s1m���R9�u��HHD���5!垢���2���|���򀭥=�3�@^@����sY�5ͱNm���8�]V.�[�U^�l��t<5cڕ�`�7&c�!�k��^�o�8x�}9ik�4��8>��!�C��'� _i��e��楡z�E��҂���P���i7u� W[��o�����?�B��QP��m�~W��0Q�y����)�٤B`���U�=H��׼M�Wdp^ONߦ�!T�7�c1��Llv?�k>���,�x);���-�:5���T�]OM�Yzmu�7k����VY��0��8�@?<��<�4{#DQY$�c����_�2C��oܽ�=�D$���gH.z}�4|�8�����Bs�^YI��V�.EX�ͪ�����z�����U�6���J�Ύ����ؑ�+�(f���^ �^.R����ރH���nת����Ɇ"}\���en��_�9�af�y}���S�tt�f@G%�#\���\�m�BH{p�_���G�-��&H�����;|Ķc��)��a�j䄼=r�W��s��\��� ]� ��e0�����֦����ߊ^���v�>=�x���u��{�aV�Ờ~�@UL��'_Q����iMo��>tQ���pX��=ǔV�{�۱�d ������D������/�s�2	,,j�Ϸ�p���s����0�H�g~�L	�R~{L�Q�#8u<}`�§dw9,F#��PX�������v�rp�@����G]"���}jr� �Bt&�[��8zn�G�.V�WI�w�Syc���d��Ȋ�дy���b�XG�Z������ūgʡv��ܽ:}N�C��ȿW&Z��>�<����E�lT��寘(HH*�SR�߳?9���J���q�X?LTj����t�m+�{9YE�<��.�0(���������Jmg�h%$7�L�a%&&ƴ�W�^����)o�:.�7>.X�mJ����hpbSN�H�ۣ��'��5�����TL�|e�O;�\�_ �c:�<�i󘾦 ��	Đ2��P0N��R�	����]8��,�İ�=]����N��ݔ���;��S'kk���:��#��M�����ڢ�#�[�e�e�4��[Y�Y#5��O8nT܏ͽ��v��{�=��:�8�5?<H��L�i�JM��6sBΥC���m�W�p�
[�����i���Z4����Ex�s�n#g<#ŗVf'e�+��-v�O�p0+��>���[oBOXDj_si��;�~>����yM��y��T��}�`��y'�qr:��
h�7[���2j&8������R"�؛����*	��#��|�p�����c��rV�m���>jz�aԭ�8�rD��s�A� oh�Ha>A@e5FzX?���ߠ���<��
8�S�L�'W�[�27�E��[�f�\�����	H�e�>�9xx<��$o��o~�}�/L�RnqTLax2x2..��k��lhT!M-+��#uS��|���׫���*�w{6�����Pq������<�9��:�@^M�@>����苆�[}�������,�2��U�5�)�q�]ف��+�e�*Ty2xd ]��s\'���~ۦѷ��9�*�9{n�u�.gTild&�Wt�q]��߬��T`�o7�2ΊSU�p%59�����S��fY��B�d6�˩��ж����n���?���0�#�S�H�A�;�йbK����V�L��6PJU݋����ȶ�*DE����z���`�߃9�j���1�4Հ'Nr�)Խ����3j�oo�%vģc~���:���T5��P����#u<�o�D�6�\�O_x+̱z"5vf��ٿ�UX���(������N�49�.����Vs�<K�[#\��5�<�(Uo�Y��b�3�<�����(CCUh�t33���
�Ih[_�{�o����퀥���q�����@b���!Bߡ��V�`��}�g�,PC��{����:�;�J���e�F>�)NDN�Ԍ���n�D�;��<���dP���C�.�
qY�Xti���|	x����/3?cJ�WB��vn�o�u��Q�>@�u��}�ܞo��d���*"��S�Qb��>L������9�!��W��l��z�����*k_+��}�*��h��(��1e<d���^�S�T浳�wm��`6ʹ�mLSK�|������ss��V�wQ��t���a�Vb����q'��H�����w+�6�K�/,I�YQ��27_�\3�����蟹J����39ٶ����LyP�`
&��D�1Z�fd�#1ŭǂ
*�9mO�dQP}�A�(EŜ�xx�i���"�w������F�6�*���/_��V݊��<�2��b7��NZ�C.μC=�W�������1�9�xT9�ƽ�oo�wv��l�%R'#�bԺ#�
��T�n�����ղ����RO�bc|t��d<�r���U=&��^���a��$���}�����SR}��SOEi�N^D��U7a�q�F+޼��������B��~�n�>���W\/QY�W���O��B.�����������&p��wg�m@*tufBذu�;uk,� �RTwv2cZK�6���6���Ļ�Z�+��s^�C�z~^#JL���f�4fOj����9��\���G�V���vz\�RC�'�|�����N�������
Z;έM��J=��,��M^�p	�ER�U�؅�6��g�k�,���Նs������D��������	��s2r�M��Ҡ�8>�n^�՞�e|y
�eU������g�_�M��[�-�I����c1���[+8uR��|�vS��x��I���c.+=m67psW��J q�������������թ��
�����3�3{�C;��U�4��,wl'���O�K�hˁ,c�ܼ��#��}9���O���'��Z�,kr�e9,VSA�Xe��V����{w����|OG �?#�"޲�׀�qi����MH!P�n��d�"6TI�7v��;-��U���S�kjj2>�)/�|oO|R�����K��F#�Lf���U^.��̰0dF�����p�i����B���WZg�: �?
Z[ߕ?���i�%�&ې\�gfn��0�3(���E��*�8.&�{z}��o(Ӫ|r��]�Ҟ�6~���}����0�,C#���Z0M��3I������Nv���֣`�q��2j��t3����aQV��`w���իTN���ͬ�r&��ʯ�J�_TT��R	U�v��ʗ1�F��rHwr���jFF�6�0��b���7��ᇚ���Ŵ���n�=�����ݣ:3�p{�\��i�r�@|.A"�>��篹���A	�+o���)��A�s��#ü��; �wpX�R��ù8}���c�U���?���?�d�z���`f��$qZ+��m��|d���АiMk����z���p$B>�!�~w�ޱM���ǆ��=a��$8h=fb}Ts����p���]TTT��)�'�P�[Ǔ:�HKSH�p�nʁY�`=��i8�����\��}��O�Py���R��%KΛߺ'��,
Qӡ���W�RPwf2���a��w
�g�r�R�vw��B��s7��!������]]]M�v�G��ttTWW����U�!�����4��L���������3�#�����~�������{�����x�5u�P�� e����=a"̟��E?$���� <tWz_���-�Fޫ㜂(����O� �/6��cR�/,9{i��s��*���έ-�̼�����=�jAi���q�Q�q��LY}S�	]�}nOy�g�6�)	��5܏�G#�ó���ϟGʘ���4�u[ur��?��O&mtLL֤S�O��c��Y>��y,+C�uΠ��g����1���P>�'�"���v�{}�=����C��e$�����̓������g\4`[�5j�s�a.�{��ݳ6������5N�s&:	g��T��׉>�YI�M�X*��|�ģ���3$�f�9����"^^���������V�����Ծ�w�0���Һ�ˣ�I�W�#�J75����Lj�8�t������\�a����8��' ��ج�.��P.?�#X \ܔ�%2j��5�
��?&�������-�T쿯����L&�74b���0z��u���-M~g��W��c�����͙y_����u l��Ru�����ϸ1�'�Ku�v"���kO�!�����
����&
���siV���_9�r�^O�A�y����$��zFڌ��ć���B��m�5΁�h�\�ȕ���ߑ��fQ��x�Qv׀~>��:'�ƕ02�y�	��)ՄH8����ňM�oC��b>�"�k�
�[�Dy�X���|NfV!>8��>��!�fk'�h*�ɝ�������
������g̿OC�L�o�w��d}>��0ukp��a��£#��jF2���|*�d������U�D���D g��%�5�3�\�������!��q��+��C��wYe�]
S��c���Is��:|�O��PodT�ۀ���IUlE�Y"��ܼ����Ŏo�dˊ���a�M�c��.#��N�Gv�M7��CS6W.�((�|`�γ:������c�3�ϲ$n�ڃ�ȼ��3�^��	�Q ������l氛�}��IW�=��� w��r�e�Ca�әtF�9�<C�"�d�u=�D,As�F1/dB����(T�ٽMΪ0t��̢�~q�qy\�>�x`��7�dG�����R �cHe�'Ӊ�F0R�HD�z�sҌ�톆���3�Hx��v��X)9��a�g!3P������R��ƭVJ�+�Z�VUmWdvK��<��@j��}�����y�50L+"��F��n��?�i�c�`�[=�Pxud�GS(�?{f,{L�B1�n��I�p�-�z8c��FٝSԸ� ffj+㠸K���Ky}_�X����G��ǐ����<�cД��`���H� �:�.�/!lJ�ϱ���%�ok*�J����:�Y�r񅕥,
����_`���zf��/�����vt��'�ͮP-৿�i$"$&.��T�{����)9��d��J�3�hoe7�%�����>�Ԑy{5Ż����U{j���)�i�PS54�\9��_�#ܙ�1nv��m���,YfB`°a�kxn�k��捩�Mr����I�@f���W ���kd���{��Yr��3g������s˩h�+�$�+?��jU$zx����d�:-�Ӕ�s^��Co5�������PA[�����l?��E~�n��!�����w��筀H��R�8`����q_;���(��yNTjh�wk������7�����6��v^-k�*$7�=�\\\�~b3"�f7٦����$�M�-�Y��u_G�(@��a���� l��9�^s��y%�j�C�sFS���߮O�C��D�7�!����ϗ��zu�B���/�E��o��gsq�췆A0XOxu癯���K�Z�`�>GÒG�u��I/�]�����2�/��q�XXX�f�z�2�$f(Ѥ��Mٯ�Z��7��LE�i���jhM�'�D���e;�iU��AXt�+�i��������������۾w�hRN��LMn�t�~��°6�D^�{P69�o#���~D[湔� �O��G}B�-�kKK�}�Ym�]��
��ǫ��X�AL�Э���-��XE��aʕԲon<�7eZUￜ�M��yև!���d���~(�_m>�-h.�>W�gL��nФa��V�TU	j��=����0��t>up4=��}�N��/s�7C5�<P*a��a5@7�����e�/MD����֥7_c�͟5��O`-��힊���{ڧ	� ]+��M���<�,+S
$���@���g��)�wjʠ��Ċr�����c��[���#�)ww�Ms���x�k�d���x��	�d�$3�{HG�h�/�K����Ǟw�!5ة�����,�駲"w]8i��)��W+����)1t�3�B*ًn ��%Fr`�箂^��f�B���K@�#srV������%����%�k��i��<���p��޹C 	��''uzhR��*�1�,p,K�z�����Y���Ϲ���پ,�� W,� �A݆���+ã<s�u��d"SDG��?'�F�w�!����Au���H6�G�' 3�����h��,K&�C�gf�/Ҋ-�U<Oӧ�|��ä��/�/0P����.�OSu�_��d�B����QƲt��<��]NW8���aG�	'���'t܇ݐ�r�*��r��^[۝�3laO<������Wψ�(������h��y.��o��?U���C\{$
��ON~�ywе\��*P�)hr��o�g���-]C��'���D����q��Ԭ�Z�@���3�86����Y��C:�S��d�ʙ"��ῖ�����5�"\j~D�j��$��m���t#I�^�KM{y�qYe �#�*'�e��������_+�C�T}�ٺ�\=���4�"�i���5�9�ҏY�Y��:;����%jv��+�T	8�T_![-��e,L<�Y�3:�+]�Ip�����l[N���B�3�� �on�8��7��T�vv���3RG��F���J�� �N�J+/���O�j���ڿ��ch��!����q'�a�ո�v2�ޠ���j����zE���
y��#'���ir�`�0'#`T�VM��m�Ad�����Gθ��B��F���u�5�x���pvŌ�Sؿ]�RI�� ݕl1)�l}e����A���Or[��R#3�וK\U� �����|�ٚ�r�?�P�a��G-��B�����8ODD�\��"M%C�Ɓ���
TP��Z�o<�(Ю8E�ke�
&(��[oE^I]�����ϡ��^A����-���V]%S��@JG����HKe51c&�d�V&v|�G��M�7
fB[����R�3��bwN"� F�$"
���DZ����j4�o+��UL�Ez���3��m��y��=�լ���Z~X4��1�,���gt�
��Դ��!�e�ʟet�.����J��#^4*����N-}h�A��%����K���r?9��7�W����#K9�S�R��J�^:A�[�*t�ӉQ�,�S�h#���<��v&/8t�l����O:_!;Q���Y�^�`����&��T�ϱ���܎%ꌳS��4����[a7���kM���o�X�(�|}a�B|.9y��?�NgH�P��4�9��������P�-��$R��?U*;h��}���������SRa�E_����圁HDB>(\�q̌�z��]?�IU�Һa�S�LaD������*��?��n��{�Q���ݻ�PNpZ�U���u/���wyrM�QZ��Ʊ���L ;J>ҵ42����s�E赛���ӆ�>�Sr���}ʫ���B=���m�z��T�H�^'�r=(>s�anK�k���
������u�֋�F�!�r��m�s6�$���H�#��cH����v*)��4Q������c�T��xmuq֎��A�}Q	�X��p�
U0�4���ɝ�R��Zv��24I-gM��K�c����2V��C��)@ֿ:������فҒ��-KW���^L�|�8{����Ǟ�Ŝ��w������A����@	��ٔ��2�T�zRA�~y֣c�Č�:G��zF`�8���
C��)c ��ޟ5����b}��S��d�nZژܵ�1)����^:!o�2yPjnnY+�HΜ=��x���u�D)�C��
��N�>c��ܲ&���g<�P�V+!�S_��Qa����d���	/�W���9�Z�*<΢2.�v�����g��	<TUV%�V�N�߂@�=�]wߓ���HŤr�
(7�c�9.��<~��jĀoom�-�v��;� B��:����߷#�j��Qf`���52�߯+����[�{�)N�7ׂ'J�V��D����Ëi>R}1��t,��Ï/o=��O�O��%7/S2�7�H�T��¿��s��L�?���4#��9�O�S�T�$y�zSOy�ꌘ+ �9�+A���z��f.U���@����ʓu-t���]IZ��$;��f�jz��={FZꛌ���9�M/��/|�Z��<sj�W���7ޮ0z�B܈��V��}2�$$-O(�: ��]�f�/=�:�������I��bϞ=oF�z�yZ� l�C�&C�r*��zե�X���ϱ�Y$�-0	\ͮat|���TQ.�Oo�8{�l�"m�D8-�t��w-�9��/]�J^'�]?-Օ�sH�y�b����ٸ��2�u���Ⱦo��{OAn�"$����Z�t�]�g�_�21�'�1 �\��"���D��z�i�jre�7�1re��\��2�����l:�:@[WS�����n�֧�]M�N�s�@}��WK��ެ:������)_�z妕����!̝�{˥�N�UHh�.'O�����H�f����1����%F�B�cSb��;sA�"�;�<�����P�<��/��<Z��̊4�gO�DQ��"����b0d��~�ҥ���U7����u>'N����|pvvf%�BU�����Cyҗ�|:�q5�g�I�|f�_垏�7�/BCKIq���y#�⑽[f:�����Ѧ9y����l�Wj=J�����6�&�q&/yZ�B��c�	1.�5��r�'�)mK�k�ۖ"��aɋ�MV,)Nz.�&]���W%��~�Ս5�p�|rǎuY�L̕+V
�K�Lcaۖ�Imu���W�\kL�+"��,e��
ߟ1���+�X�n�3�a[)*���C�T�0,0x����0a9�i�w�u�wk�jM劅��5�5 ��=��1�M�VY�θ"R��ƴ套�n���O��'(�pA��pee������)}fR�a	�(Ο>�X�3 2\�������
U{n�j&(�z�[����S�"����*m����S[ר���y���x��M=��K��?��S��X$B�Y���!�nq���k���T���_�*=����_\.OS��+��_��<;B�0�c�����jk*�����#I���IK��d��[��l2�h�6an #�bZ�9�c�'�r�tƹNy���*���F]㤞�f)���+��˕��T7���<�*	���nI3��I�R7�(�+�W��"�-T��U������;v�R����cڢmf4��xW)�c��ee����Sb:[$�3���>���xsKˤ�5<84����[����Ϋ��i\w���	����"���_ֲ������o����;::6���BD���8 ^�(u�8v��U$�<���s����k�Mc
��ܤ�i=}d�����E�lI޶�`����m�2�7���1���d23R<KJ+�
&�hF@� ���z����0>-B�DW��f����d��5ɯiI��#OĢڗ\8ޢrB�� `�	���4ע���\�::��Un}D�NO�ݎ�{�$YyT��(%���5Siij1`I��9�|P;[RV����E땎w��+�6���;�Ҹ�t\Z����)�^&�ڙ��ii^	����#ݓ��_,��b�
 b�r��]����
'$�9.��Ȓ�%c�8HQvthbrbtIcc�����[��^gmM�E����3����S�K��1 _��Mz���������=S����{vff)�X����	�SjJ��X���zdˆ�𳯼���Ʀ�o~4Ww)�_��L���@������Kg����4a-RگfY��i ��y>V;�=�t�M%�:[#�T1�i���]|�M����-)Bi���j��1$F{gR*Ϝ`�ҕIۊ^幇�Ɂ�=j����8a�Ȳ�>���yc<w�8G����X���&�7?|��m�X�q�����[�j�)E[�	
dzfJc����PR:R�>�������K�;�m�m�,��$-�9�_���z��]�Խ�(6���J���S�_��Y����.c�]��K���e+V��jx�^�?��+mW$fS3WZV:}�̙	.��Q�� �&4�=���4G����~�<.�O�ӄ<F�������>7�0�����	�.��+7��={�V�9�Y�]��JD͢j��[�]!x�:��F-�[�E�.-���۰�E���z������M9��sǖ��#�p�n���P��D�M�s�� ����A��	x���d&#�v����yDm���셗ݻ�{"�.@>Q~8���|�+i�VX��L����7%��{A���j�F��o���b��MJ�t�=7�|+?1DȗH�u�m[��oGH��|@�{��k�k���n�3Q��H�s��H(���qϩ�����}��f�&dzr�Ho�	C����ҧ^��?b��q;;��J'k׬65<���	xդ�|�Z��6�����nٲE2��]�{�H���s�j�
�9(�x�B�榾E��cJ[0&���/���DПWDc���gL����3�k�_�������G?zJT��*�1��˔�WdT"8&������4�S�*_��w?�l�/��^�+�� ��� ���!��) 2�G��� �5&G�©�i��<.���8�)�/Ƴr�i��t�K�|����dY.�����r����_1��"�뛁�-��r��h�S�B�.�� ������̳@�QX���0���IOau�ccc��Pf[�J�X�Q��߳lq����w�.Ĳ��[�lٺ5y��g,�M��ͷIjv$�F��_Ug?-ag��(��^�X�YQY�$u�ˣf'O8����튱��)E��t?v�h�����i��kR�Ѓ�^ v~`��]���˖&�~���G}T�N$oy�C�<�߷Hlg���w?oQ�[7oJ��ݫ�"�ݪ��1���u�N)ש�^���Ү��2;u|��V�����4�4W���At�U��9�*1�8�16<<2^[[;"��po�y����.������_ږ�4�g�+CkBF���zB��|�H;@9��q�����gÃŅ�t$̷5��xtk�jqv�t�aau�OÕ��ƿY��V�E�H}ѝ��k@=��ǆ{�]&��9#�9�{ފ�K9J�D`�EIT�j}�@o�ڙ��I����{�K���[	��x�U��`@�����Y�ح�C�`G[�R�����\#ɝ>}:Q�Qy�%��ǈ��;B����y���[H��[oݬn�Ɂ����G�<��7)�k�sd��y�
�www'��#���e�ֈ團��cu���:�ᕛb��g3�����*O��h_C��%w��K��煽�ƥd��QP�w�׾�M����6k-;<<����oI��y>9�>�Eт��Z�n�~����-���z�����dtb4�}���ܹs�JwI��`� ���x'ٸy#�8������kWW^�x9�CO�"&�*�S�@�y�Ҳ��h�r�RF�2&@�w�#�������]�W�a����G�5)��)y�ӅE���Skډ%�����|s�W�h�}�ɥ��~1�W�M��b�3E
��*�~���B���?�'��r�r_Z�|���3����Я���[|3��qyeNf|}�ާ!�B[�����۳�_w���B��(�;�h6]Qj
lΜ��C��ؼ��Ibϖ�-����ȫ.Uh�2:�|&�[�1�/�0���,�ZZ�R0�)�j�@��ٱ�6��ΕQ`�9�$�Ǟ>uZ*q�f���0�x��M�]�Qm���\
���Q���4�B�}�}��dH���
w;a/���}S�μ1v��wɩ[t����N0|(�뵼{����m�:��O[8��{����ߟ�ر3��lۄGp�]w'G��>~׮;�C2Z��;��*��8�� RM�>wW����'gՖg�K�Ly�|��w�B�^�kWr��!�ٸi��͞!��e�_�I��۶�766��?��~����yb2`�����qB�>,��:ߍ��UzbT�b�Wi��T�����u�5El� �/~ä�9N��~W�`��S_�mx��¹�O>�ĻTz��N���Y%	avȢ1����c/�A�E�_{�z��y�[����"<)7ːڎ��s&Ӎ�t�co/9
�|���O���փ.H�eZD���������<6Ƽ�oA��m�::������q#�M�I]�@�h���/�sZc��J�$G�3DYP~3�X�2rw���89l�Ve^vF_9i�F�3kHD������5��%�8
��&�^��� ]=ɥ��wNc���9S
���$��A�P�k`vJ��\M�i
���	Z�������F���G�ޯ�>w�ܑ�ɰ���@� ��_���}=jz#�ٻ�g��>��`���eK�%��s�<��&�K�~��}�o�|.cc��v6�*ߞ={����������Æ55��ַ�֍JYd4��I�*8�#jP�{�����W$`�"w_3R�9o��RҿW'/?������q�����z}T�߫��T�A�/��/��\O��>�DYE��<�����6l\��o����y���2��G��2�C�T�p/1�v��9�(1$=ס���I)+>]��K.S@�Y��Ep�}m�jg��+���Զ����&������M�] 8�f*�\g�s��&b�
ž�'���p{6�>0�f��db�3Ɍ&3ŵv��Ma�K�M�m6���>*p0�E9WB{x�� ��9�� H#:���hQ)ؔ�늑�`�S�N��
��O��屰����6��U������WFE������YԀ0<y�+j��5�4�[)4��7�H��H��Q�Ot��j��o<߂�"�����-��Y?v��c��w�|����=m��ҥK�*�.)\�"�<� ���n�� m�m�� ����S(}��l�9�;��'N+RP+U��3=�Ͽc�v#�]�6o�9)�1_��X�R��w��@F��(��'O��>�$>�3G�zEZċ8/�2�8^�:~�|Ν9{vB�ҸB���V9ޠ<�A��	��_��_� C�*:���ʊJ��+3�ȟ���<��Y��뇡��z������^�����r��hz0m��b�8=E�p?��q,�����������/.[�tQ���I�z�Jo�qv�WLN,��X)�!�k��d�0����<�#�\7�: :�z�܌Bdܐ
uȘ8��s3�y)�u�$˃�fJP�p�g0.�^��/bX�ڑ�����l���dbZ^�>�Z�o�,���r
᪆|�R��Q�N) d9~>':�Ǐ�з �;��Xyظ��)e�W����_!��9db���E�8�V�L~�g������Y��Zx�T�,V � <[4ݧ���絸�t��|3&e$(\YQ!IY�`<T�1a `C�X"dOnY�Ύc�T����q*(2>�[�5��ƍ�l_lg͚��&�&]�&��x�[��o�]��k�Nӱgηo�݈z}��;�3�d ��$�K���v��.<��K���IM���!�꫔>�XҘ �r�;�<�Y��geUUζ��KTX261^��Ҙ�u{_m�$2�fT���G��z&:;{�E��a@M}�����^y�]��W~����6}�S�����+�d���{��Zw��§�z�}c�#ߦ��2�1�����<��R���9�H��քi�!�[�|��[�v#d�E�H}ў�`S�չ93�����f����	�D]�`~S�b F�?=ʆ���þ,��a2J`s
��}���@����+�4��]�`c�`e^8��.�#�} �����.m��`j�c���������Y]Ke�@F��
�v3l��s�ԣ"�֪��H9������8:���[��f��U HpF���*v���T7�\��и�T��e<�=4���1��x8��)k�~>^<�m_��2�|F�ɶ��A��R���U""T�ϋ�n ɜ��3 ���.R��P*�Mn��y�������0�ߛ����豣����l��6##2��W,79����9�{�ט��r���^�mc� �Z\���U�c��^���.㡭��"
�J;l�S*A�:c%�J�`\2���Q�6�S�~F�Ϥ��1� �O;~QQ��">&c☌DLft�S/�5,�O�\/q���e�c��"�h��9�'�`�F3kQ=ݳVQ�tE��$�����wδ���.���Ww�c�˝�)1|X��Cp��n���u��e�$�aNݔ�Ӫ˞�W�m�;��G��%����kBN=��,�Ny���D?����ǟH���uךW�����^)���G�, !v �E_�V��H��}_QY�v^X	K�|G�-��T2��OtvݹKl�R�BZ�V!�!V��zj��@	������<T��t��*�K��W�*�>}��Y�ВgL�����X�7��$d�@�˝�xf�TǛ��_�4��B�ʭU���1\��4��YX���Bs�i�2�a{Ξ�	��O|�����1�D B�ce��GT�D��*����[7�j
|��j��a���c�@�=w�R۶o��50Ч^��57ef���<�2F�S��Z�{@�Q�;�I��u�m2�TR�������'ߠ"3�E�8.�O�<���Yt`��F������,��Q�#�HeuE�W,��չ��(_535s�������
�RD������.\h���t��j�r'�KJ�**���Q�~��(/����v/?p��ֽ��Ȉ��v%"ey�.��i�^�9D�t��R=*��^�f���S@����n�5�@�œ�/=򙦢�9)9��z$��|3.���5`�m�`�|@l	�V�Q�Ή-�m�Ùg� �Oǵ��	�vQg}����9_���t��I�$O��f-�>�P-�<"�}�B� 	9 X�zۄ^�Xx������ї�	=�����#�� ת b��8�8i���;��E�;�y��٣z�ϥt��K���K��]%�mO�06���@,�����-*�9�c�-L�qϊ�@�:��`0mx��W:���H���^~�@�<�"K�E`i	��w��������9%c���r���������+��B����a��!uՐC���D�[���4�U��<�����gp�<��{F"@��o/#_��d���e�2�?��.�(���< ��W߁���y���S��Ԩ�P�9����
+����߽~�����U<�4�hEe�Jg�*X�A��S�3}y���u�����J+{e5��U�����OV����L��낽��O�߻g��x~��J�M]8ƹ��ɡ�PhKlyr]W�~��u-�r@���5�����H=���n�NLe�F֔�$�FD�hjy��q�9�2��&��1g�%Am�f��F]LYM�c��A���s��R9�qi�l4�_c7�7���&/�8'E���<;����ɭB����E����X08�_@o�<-��ejɗ~tWg���J�£��	�kfb�r�3��	��lA�m���9+Ւ��g߿m˭�D'�A�G��Ήm�����~�'2 �7N�Kw/�<�����֥ä/0��\���H�#�(#@%��#k����l⑕��[$%DIlr9n4�u��|u^�X�A��������:��řpJ�i��9�,ڶ@��р�`nJ} RR/����(�+)/��9�U���|mX��8�O_�B��"#����'�>,�&�AX�J7o�l�����]�lyr�]b��7C���_DU��B���ʫ˿���ߥ�:�o�j�/hl5������`�B������U5j|��t��������LEY�huÆ�����le�`YQ^_yn�pEQ�В��֥u�_:?z��t��(or�8?wX��S��L�{J����.�k�r�����~H$����S�A�0G�=_�4ר�cֵ�q�QZ,C4/��=:��њ���e�V��8|=,�)�_g����P����Xja�Z��`�Յ6���;z���h��1��u3� ���zր�h;������z,��JBj� E^~i2�E����Z��h�J(V;� ������ B����,�*�<��#�s >�R�x�Z��R-H��5x���ct�8��E#�=��9�η)O����#��K���b`�"�jnj�7�<�r�Ӑ���Sm�0h�d��7�pt�`��k��:(D.���`��M�faһ]M^���!���Z��xb�`�"�vD�@8y��7�<�F�U�v�տd
`���G��/w�]JɟrQ�%�[�hː*H9���b�_!2�G�Z.'���O�<~ ��:��]���Pă�9e|l�yV������z|�gr����`ꀛ��'�ޣ�����+��:k��G��a������p2����0�Ju[�����������hD�����#2�j*d9^�����o���_���gE�lw]A�@IA^���p��0wT�W��+�|\�����֜L��f!�������E��w��������u�����U 7DM��.)̧�J��ez�j08õ�{�W��ϮY�������~���l�
ea"��S���C��=�w�~��2�9z����c�7I�n_�7��1B.��3�7tq`��T�6����G���P�Gɿ�����}�I��}��\}S��ȭ�x؄�	�G����aR�,|mak�%�" ���Y���#G�r���+���j[��(4����ŕ�yW�}�B���zdP��뤀��0
\=DlӸ����,�1r���ԀF ��Mj;��x��H9�Tz��>����۶G�j b���8A���V(C�$g����fC�g<��~�	W=����&⢜<���N��\,����ǮM�o�ڬGc�s+�"" ���`��meH7,_����T@�B��%e�:`�S��|�/+.M��*MS	ё6;O0��H8/�L^��B�/U@r�����G���j�)�#o�{�s���6��1��M�\i��d,O\�e[�LAK2*�tD���S93�I�������+Kƒ{V7'�˦3}�9�D�\���99c��E3�u��7���-�aH|�n�����N(�q����]�e���ܫ��l/Q��C�t���?[�h/ּ��Z$�)��Ki��F1��IM�	��R^&�<*�[���n4R@����z9��r��V�'�	d�����γ%Q�Dp��{~@��g4����/����ͻ��(��	�]��e�m;Z�$�
y,ghL�zeR^)��Ay�z_��,|��IB���ٹ2���%@QoY�Td�E�?B�sj7g���Ւ� @J���ʷ;����ǉ�� 5	pi~B��A��38<`,p��N���IJ��`a��+�<yU
੏(�P����Y�`��hTŻ3��ֺ�䘯���,9}"-0�1\��Õ13�㛙�0`G���7���P4p-�X�6�#_0��S�3���}�sM����S���p\����+���	�W���1$��JL�@���Q����=�:��X�2<��70�b�� 
x�Љ �s�=V��N���̉���I��}���T��-�����L��d�XFԚ����6טf��Uhߺ@����ɘB���˿��,)̨l1W���
Mo����z+ tJ�HKXF�;�N�u�:�?��x
O�:��ʓMK��_�5����\��ߢʇ����٩P��M`�s�q>��y כ?!�:��j�jv�pC��߹�����x��}�����\��oj��'%�1W�Z:�Z��\%��?w{C�:���[��܄�(d�h��&ܫR-Nъ ,��&l��6�&��Ҿ-{,,�[��S��Ŏ�!˿�
ԋ��U*{�hӪ��$7�v-��}YH�s��o�:5J1�<�陌`�����8�[�C���YH�\��JW44�o۲͆���[�,���mp`8i�kJ�6/S����2捖��@[G��!�E��<��Mv���$F�W�/x�r;�s�X��q{��!�;44j/��}��2�:��cw�<�m��{���NX����hULY��!>� ����2գ;�N�4��jB�s�� Њ
=����I^٤���ock]�4eB�
�_"�X�
�?�G>�X	\)��4`�4��'|O�$W�7*�2&4F���r}!�AC+_�[��v�J��Ym���D�ߢsU���ڮ4�-:@�[��4�4�1�7K`�}��i��\��2 F&f�6�����Lr���|UO���_�0�����iN�eF��\�K�n]����8'�Eh�����{�\2��Tf�$�5��c#3�3���4�o�.g���x��������kzs���:�~�����4�[L4ƺ�yJbd��c�C�gTl���)��g�T����6o>�M-r���)�_�IOwi-|�|rہ)�e�p5�{�ʣ�K;�OYv����l7�yB���<�����|n6�>�gGaQZ{��"4iR��9y��ʕVH/�@J _!O�.[p��k5��E�5�5";�Ȱ��M�Rs-�8��b)�<C�=�H�]�I��@q^Y�^r����z����,������,�m�_B���:���Zw˵�ʠ��fD v��
�
<����,���
��+3���240x� .~3�o`$�f,�=
+%�>,�<^#��!��'q��y���S�դ|7c@9�hA��YG�$\���0bDx"e! ��4�y"�j�f�/��	��vW�yW��m�}�1�4\����ijz���9��.,ga�^D�N]D]
�K%����֯vNtvNzbu�j�.�~�J�J5��g�u�\d�+	8�x�kF�ݟ_�c�I:4�I�8� ���j�r+u���79�ӟ���M�5���yE��K��R�ʊj%��o���F5ԩ���{�7���4��������������N��֝>}����/�����UXP�
���+Q�v�n����<���������܄_\�v��֮�8�z��jo?��=���^�Y\���+�q�T��aY�^avk����e� �گ�;��|�9�绡�-��<��������[]Ⱦ�\}�.HF��._%QyN�N/��T'�f; �QYY��*��	�k���4�0'�t�� NɄ��
y�X���H�\� "O�rF �O������ ��cyym�������_�~��|Y��ۑtt�xT�O��}�r�y3�J&qV��3����8'�a09��i�^S#�T�.)��9_H�)��04 \X�,� ��;4���Рr�}&�9�c�9^�j%2�`ף�OH����̈��9R�yV��<6�;�<ra�'���C��ǌ��#c�������O��"_���/?�{�Ý�F�1�5��r���bxOٍ9YVw��pFs��5l^>�H_�~��F�&CgV��%��Q�ye������]��=ׇ{���^���!(z?mC9���q��J��9g5w�l���Ye[&���i�@d1뜮�K�����Z����$G��S.�v�AF���ַ/�^�ճ�f��Ί��d��{NGeE����AЮ����V�D����Z^�^|�[��w��� ?��CLב	�`tZ;T?��R!��B��+:x�L}�Q�{��6��{����(>���87� �Y�����qG�Jw �jn&�by����L	�����"|v��/��lh`a���Q�!�|�!-Igs��h�+���7[��C�Ceh���sm�:X�W�����Ԯ�X '���'s�p[X���� �����s�^Q�[/ֳ7{qrϴ�p��eۄg����#��=��Y3-�< 
Hs.��>^$��<ȁ�Ɖ��g 1r�,���23��!@�R<�ۖ���{<�:����b����d���7�C�v	���K� 6<�Mn��֏W.`�v�< 	�6����ɨ �25 b�X�\/���ǔ��Ȋ\W  �t���O�W ��	 /�yo�GeczϘ�2�,�>5a��:�83YQj��y�y|�g ���Nx}�>�6��.�(��ki� ��/IP������|3e5��Ph��%�#Jg�SU�`~�@���9u$��I��HrZ���*g,�֭].�޽�J5Ź]$Ji�+�c������ <Osߓ46/IƺF̈#�AU���,Q��T��ŋ���'�xd����J�/ij��	f�m�� �K��?��ǃ"�S׏Q��Ii��i�(J
�ȗ�8)ȭ�U'CX"E*�*�d��-���9����]��Т-
��\s�l�����mDv�fao{7(�e?�� tJ��˵Pq��R��� �Y@��ǝi�$�> G��	Y|�f�7l��LV�ߑOq��5D&X����#�����ʑ�yY9�A��A; :��e 1�N)��~�B�4å�&O�E��:����f�eȵZ�bF����x���Bs	>� �B�_�k#��GvV5�MK�a	yk�]]�,7��|3 �_�܀�x�<A�xkDH�Sn�)�~�HĦR��Q�}��ϩ2q�T�����Oh�:sʼ[�� �G�3O�B2������~.i^Ғ�P��1Ĺj��:��@�B��yF�1�� j��">���h@^�f\�8э*��Sy�g0fH�dE^dѧd�˥V_0"i37xx4�K����A�! �ӊd&�Vxu��<]CtlOb0�v		�Y.b"�
�܍ � ���az�FQ�k�E��1 �Ļ��9��#�e��
�W�k��$Gex�扄�ms<%�:R	��xQyrrd6٬HM�����vۦ�g^L�D�����(��|�?�Ayy�y�%�j�O�8��q�9�i�KU���������K:������i5�9���ܧ�|��66�{�*����NX���#5�i^o-�'nm�ə-��T������*�b� ���/41�
c"3է����mۿ�z�z���G
���y��G�0#i�It�%�i�e���%T^_�[;����K��8�3�۶=�n�(H�ͨ�,�-�,���V� ����l2,�bx� �㶝II�Hn��ţI��.&Z#�Z�v� ʨr�x��oii6uP��z��9t��J�F�]�͇v[��.i�h�{�;į9�ݏ����vc�6�TdP�pK���
k��5��A����|�lB��<��3g Wv��c�M0��ja�j�y��U���׃�]��V7�Q�Fޚ}���^��P��J�\F=��-�A����39&p�|����	y��ͨ`�A�ynl�n�Ĩ���N$�^�,��fMsh,��>LɜDb�4p���Ԁ>yj  � +��7>!�"2��(�L�f�B �x�<0� x��	�����`Ml4����N�ӫ^�o��ǜ>7+��\�H��Y�g��&k*c�r:0*�^
���fW�F5��Tby�R��Q	g�B�S
œ����(�N���v3IC�T�t͞UY��۷ۼ��%�W!j��R Dx8o*i�����W*<�5F1�k�?��'���$��-�?v�:���k~�W���ӏ��" ^Y�|yǖ���x��|��R�H��^x��o���4�Tj�q �+/?�lQ6�u;?0�ԉ��MȮ-���c�Z/��-[�p��m]�����|���ˢ���	��������T���/�=u���Vc+\�k�8��3r�8�������}�m�S��d[r��hݻ�� �U}bV��E�2i\�29�q�=Z��m+Y F�u S�O 0�S��-�m ��!���u�[�n���e�ڠe�X�x��� t��X�q� ��{.y��ߗ��9�
���ΝU����ݧz{@�| {: �WM8�v�Z��5�&<��m]dF�7�w�o�/�imW؞�)�.Mq�W�`��Rg�'��"��fF �g�H�(c���LM����P'�m�m�3��j'{T����~)�uZʀ�m�F��vy�{�Rz���ǸB��-^�y2|��<���W�d �$�ʹc��o�����7` E�� "E"�aP�H��Os�qy� rEC��AvDoT��Y�5R�/��Dz��j]�
d�1���[�:]SccqA$� #��wH��18��1~`�p��������H�ǭ�g�ѐG���0�E�["o�i"/��O2
MC귺�+�$-��O��E��_ #�Z�#������EX�7��U��_�z�]���~�N�� !��6�u����K�?P����f���������}]=�t�܀������ܟ|�c�q�ϯZ��mxt4O�xM�����t>�{y�@���w����Ǡ$B�<06�k���\/�M�zs�pp=œ�"���W֬]������K��jCO�z?����K++�$�ت�|F�4��<���r�; {��ZN=|ž	J����`'_��š�Sg��/61�/�.(eK��7z����E?�/���Y^٤�����S�˗)�i�Ay�P��6D��X���1�5 r��P3��]w�'@(���A�bA������"#W����=�-�ˢ�`�X�r�y�u
�/SY]�B�ݒ&e��W���,���)
s,�Y�*OW,x��)�@%L�ǘ(RP���jW�X�6�OjLK[���jt�~�ÂN
Uj��j&#�5�X*lK�G�DfL��yPmugW{R]�/���/��I���j�)	�6�P�ԯ���]����-w���Q�1 �lǝ;���$��8:������i��\�� �c T�ؐ���sȌ��9w��ɱ#C�9��i ���"9Wv.�M ]|S4�Z����)��O�\�&��x��<�=n�N���pma��������*FU_4�,�5wa*� ���H��
@���;���S�x��X#R�|����a�t�x#/������W�����\�b���
Qr+������&H�8�	�(�쿲��ٲ������ޭ��8{����W��4����m��,Ҷ,j�|+�9�Z���Z��=o����2~�R�5�~z%�qat�NL趞zT���������u���l�)��g�:<���
�Ry��$���[��lhq�0�n����=�>��xn���Ey�H��[ԇMXo"�3�}����N���o���=��X�ᇕ���P���Q`~6ɗ�FN�E����zf�!@�qr,n�g�� 754��p������N���dj�	/�U�u���,��E[�1���~?�<�B�& CX�8���b(�Z#�9 i���k����L�2�I�h�,t�Go�"� +s��" ��+ c��T2SC������~��H!ԪSY����)��%u*;"]��.�����	O�1��󯮮�5N�Ȱ���:�w��FÀ듶���|�M�t����D,z�}� r�.JЅF9:4�a<�2_�w�����%]�
{�l�l�}CDA0ڔ`�h���x�p>�p=4,�PO���5����j� �5>�:B���/��<����1(x�t��eq�v�~��!��J�r�a�-D[ؿ��!Cj.�����M֪����z����ȏ\��O����uK�4[$�q�!�m��g��4X�b��g;wȈ:v2�HU�o�4f(��T�� ���Ϛ��ɚ�a��eƃ�bS+��Ϣ��Z�˂5��&���M��]Դ�)]s���*b�um����]�K��r
�7ʙ�Ύ���l\�� @��9)U
JC)�-DDm��}Y�	vr�~sGҚ{�|xZ5�3���"�,(ݷ�(���^�����l��t�?�J�P��䌖��~-�9�$�}<��7ko�:�R�Z����� �T��N�?!Q1.��c&�	�2�1-�������h��4�	��ƃ#D�m^�ۦ�;����в�J��<$�c������ƥq���y���(���n�ô���7�w��l䄅�E��;�j�3�d�k��p���k߄�����r^`�s^0�dH��ϑw�`N�Kt��֩Z�+�U��$#�ojl�OU'j�G�v�7�<��J��k�$���z�K�n�_��.�f(RЩR>���Ƞt����/C���(�>���뇌�тZ��V5�a��	?�6h����	;[�_��Ij}4U�D�#*{���ӧ���>�r��)�떬n�B��D0�)K�'tQ�G(X>�� ܩǊ�ĵ+9����	�����e6�rN/��diF�����Ъ��jI���`�ݺvtx��w��m�O��o�`��vxp^1l�,Ƿb�*u�7������=LS����E��gO�" ��Z�\�,�I�Y�~bH��N�:����s��F�L�k.\(��i9��ɹ����K�;v�Y�f�5���Z�w
�Wk&���jX;���~�s�nLw-�A�]�<,��_2č^z����<�Uc�o�Y,��枳��x�����2���a�� Ńp�8�K�-ޗ����lO�'�}�i.�҂ަ��.[L]X�YZk��4��g�w�7Y����HR��?�tɣ����汖��}߹���ܙ;��r�p�Fm�6˪�"Mm+��?Z�@�"�?mЦ1��(� A��u��u'2$Ɩ��Z(Q"�!�ې�}���]��{?��wΐ�kWtH�C>�����s���}��{���}�x�F��d�J8	F��� ���a�>���o}�[�7�K�s!^D��8�~�Sa��0`��� 7\��vK��ʉ������\ۨV,��@�;�����4��0 �칳!��'�V��6����F�umצ��,!�M���hغp�e�)����g{�c	�̬��;3*��E&F"��_N���$C�$w3��{�����F�Z�t�8�C���/��Mc��������!�G��n���?N��4G��Z�v�2D��
�m���Zɐ���ѻ�\�: 8?�@@�"�s6�SYX3&SSW�=}�IɅS���M��Z�=���xJ���p]NF��E�Z�.��oaq������]m��Ef��>�+ [��/����,N ��ՖU&��0�4��˻��g��g_?Cf��{��U�e�^rE���.g��g�N�Z��u�xq�Ҁ�OV���A�/���xe�Z��Ϩ�E�H�~��#��ݔ��w�ǿd�|�Y��̗�����ЃO�h_͏O����P>��D���ѱ�u�|L���k���T�F�D�5�{����n���iJ�t1��H����&�kN@������Dko~�`��T�֨1��U.�چ�41�{��^����s��4�*�nk����^�RHqkQ�566uV�㌨N=w�����|���|�U�8�b��[�W�=˸G	[��M��k�M�.aܬ�^�@#Աe*[W��yY�WLF��C>��ݍ7��y_��{Q��=�Kѓr��7�]?,��Ǿ� ���I���kЕ����=��r�pEw���^}{��y��E�q04��a����xǦM��t}_��Ld\�!�x4��+j�L��P�F�u���1�V��73�\G]����jl|�uZ�<�}u��3W'�Sq���u����#��q1�r5���r��S�p�\d|��V�j)�r�U^#nmd= 2��a�%͌�F�<����M{��\xa����[�g��#m�NX��QB%��E�۬i�HO�q_Y:�n��s������}?���w��W_'Z�F��B��ԩ��+��=�p�y�:u�c��[ɗ�	u�,��11KfF%Lt�j�W�p6C�I�MNDφ�Ȕ�Ώ��������V�m{Z�n�2Z�W	c�=e2F�K+��G�w�<�s׾��1�s���P�^o	���ǆ�_~miq��*e��^,���Z�;&�/�����ӌ��,��t�����L�Ŧ�ƻƻ��ţF��4X�5�ڛMb<L����V&f`n3�������l.3QS�w�^XӮ��T}���ڶ,�L��GIkU�)^�z-HE��i�}�����L�OE���[g�>��¹4Q����jD�כּIX[�J�C]0~�կF�����L���j�
�hh4JۨW*�����*5d�늼�Z���x���&��Q�mɈ޶�`sS�\U�|:���E��lC���r�G��jǾ���a]��)_{���
�q,1�F��bWF�F3����C�o�z[s�~~���F'� 0�e�ZK`�#f�����e����jۓk0�l����d����h)�̣�f��ߦ1�/�~�������(\q�>4����?�l�5���d>�o:�:c�5�Zo�����N7�z+3�f}NA��WI���`�������n��cн蛨4!BӀ�z�s��߉S�Lǁ�﵃��s� ����}'�.炠y�����f� �sN}��|�6�^��p�.^�0
'Qn͛�Z<��5!˱�,Dc�#�o���j�k�[Oc^E3"z�5�����gP��r⾓?y?s�:�[2A�����G�z^xl~�⧚WV��CA�CWi0���Z��9�}���D��#7]k]\v���x��bՃ�U{���
����5��(>r��.��,s��cXLQ��FRsz�ru1�g��cD#��c�21��++ZC�1=O�k������`;&r�f�_����"��Ѭ��.DJٍ�����즙'�0g`���-�ʸ�j�u<�Ik��0�D���Y��I���5g_?5�����W'��5m�����*%
b�'.)�V��|Gd%/���R���W��R*�ͫ%�Ī��;;0�D�J��߸a ������dC� ^�mw��F���;�L��˯�����%Ox��NgC��k5�^��&r���h^ǥhҗ̎�wu��9�jbjK^%�Cf�pH|�F�s�>y���c�=�c���Zߺ�jo9|���.e��5�֨m�
'��h�Ç-xW���ͣs¹�� =��5�c{��
:q0� ��Eߊ�'Q���O�מ����|]We���2����*%j������^m���R��N��� K!���SYp������FѨǑ�� �l�5�ٻ��p^,UX�����q	�z�w��q�G�kZ��4謉�:U�������'iuĠ��NKeE	���.���تS�z|N�̭���]d��Z��h���_�ү��v�a��J��^�"��t�۹�����k���4կ|�.\o��ROwS���~�j�j�e��:6E'�I#P| ����=�M�=���F���Y�W�x�"�k�>޳DEhv�(I;�^q�i6P�
��T�Ge2k|hЭ'k�� W��������n�i��3`k�Q����a�;E�c�c?��CTL���Je6�yUֲ�rfd+s�ګ5k�l\G��9�n"Э�����fdܻ�?�F�5#.�v:%HIJ��@�&Fn��:X%r/�u�\W(BZǉ':�D�.�r4��V>{�K� �"��L�n��*Q��o�b2��I�2n&��@�lE����ђf��L�-k::/��b�4L���
#�W��ǌ�n��^F��ځ'�rFj_��%�B.���HU�޸v��jx�)C��h-܂P+ӡ�x[�dM�;�OgfAb�z����$i��^|U[>���I1��g�2�l|��FZ�t:�/b	E'�LFK��쑏VV�� �°u���	T�i�Q������Q�o��tB������~��y+Y(p��8]�[���������F�Jq�F3)%�^��^�qB��{��54��$��X�wzux�m�B+���|��#p��Y>{��^2r�xF{�Y���_>t�~���\|�o�i���W�=~~���v���Qp����q�?�~X����-����ˍ^�Tg���̋���7�Z���WS�)Ʃ����|���Z{�Yj�\c����[��T��(�����]�ؚ:,�\e�n>FKF�a�''J�5��5ʣ���(�{FH�[c�`kX���qb�m��(����n�c7�i�b���PeKkj"8Z��H&HgDKEӾ)j���u>v��R�ss�˗�pN�C�ֹ�O5������0��u�j��P�=���FR?�s��]�h�)wO�F-�H6|%.��'����D������7k��Q~m����d�Ջ�k]�����#�1|4ң��,}8�v]_ei{)C�2W�5��#��o���(X˾@	�4�Ƕ��sݸq�����h�����x��� �h�U�<�pV�G��
#�I���1kbm�����І73�����"��?0������)$E	���ft��J��m���$�~�0��Ӵ��m��K�LT�t�:���B���KD�rCl��\tV��@x����҂)��V8�{�A�̾Xc�$3���|�f��yT�a(���
ϡ�	'��6Y�4�P���|�����{���������Y����
���z�'��Y�/�4�D��ЕJ����N������k�}5�Ñ�[�-E�,Zk���ln���i?e4Mavw��D���3Qw	��(���w6�H�k�c�pci��1y��!z�1@��,ͣ�d�}�
��R6b�X]6�Q�@IL6�xbS��5=6}��<�G�����t3�����$���+����ihS�Fi��n^�����k�t8�q&L���秹	�v	[��֫O~ꓕf"L�U�f�SQ��lll�JkjL�fJ��7R�n�F̦�ݬ��C �hmÆR�i���yK �}D;6|U�J&�+i��ƥ�9�F�V��0V�)�+�*Ǡ4«�T��%zX�����w2!,�dq����C7���x~:?�J���(�=���%�$ �"�yc0�)���j�4�[�n�!2����bP���
�{��%f��s��S���C��֥No�9�;8ceb��3:�7Ё��@��6�#r6��#ʵ7�[_��0���lK��zZ�*��yb��Jz:�@u�ѩ�C���m�ef\��0#r��a��Ǐ�����ALa;x��?��I�Ȍ�����"�q�.F١��y�� �T�g,��&�j_��4{�w%T�����/�\�1xl��]�w��}�l۱�]��~�d~IߤA�%��}���_������.��m��� �a-ٴ7���˔]��n�Q��)7� �ųJ�D7�0g�^.������x*�3D0�H_hh�\�Z�\� �ۻ��F�B���J][���[��� 60�Cl]�t���:q'��k#86b��F�M��[��<b7�f[����x_�d��!>�t�ɨ�������1�D*c��{{�M/;�LC*S{��)'����J���%g����Vf���}�qU�T��e6w#�5걦�cd,��:K8 W�^	��E/����`		lK����?Md�*�d���t���9��棾n���aʵ�>i{��,�lV_U�s�h3z䥾�eڙu���R�Yô1L�.�οi���x��f2^u����t4��f����0\�l�x��=e�Z�(>|O����4��D�:eW������L�߂	��[Y��~㏾9��1q �^��4N�"�c��ȹq;!�����ǭ������`�K����1��p��rvklC����2����s��E�̖Ne��M�5�qh���c�I�׽/�*����+�?���`�?�����~�5��o>-��G���>0s� �:b:/b��4s.rt��)W>/�q���"�۪t��I�ś�s�q�\?�<�����>����>���v�߃�q�F��~��+c�խ-?��p6�U����������9�X�K[�����J�<lb5m�7�]2�U_����E�z�%	���y����c�`N�w���wK��YR���k0�!��)�{6Ҧ3|��ݻ�V1���D(�	:�*�4c�fU��%|��Q�%�=�>�;�t&"�ԃ��N�k:�����ꪬ����Cal�t|U�6"�n�n�w3moj�/��o.��A"���%�;Lݴ�<�x5���4��0�f&<�E�x���z�'&�"RӠ�����ϑ��٭���Kk1���c8�H���6aԯa�\l͋z��E9`*��R�5h��F���D"`Q,�����ILO+5������%}��u�� 0�/������̀�-��Q*wk&c cjZYe;����;C�Fa���D�֢_e��g�U��]�z�v��1-N���/m�j��jy�q�u;ޔ������R�r.�ٮ"�\�7Q��b�X��|�������~ �
&�6x m�����ŭ��)���A-*�9|����ΝG��?BV|k�M8�8X~T�k�%�*��|���]
c�c�^c��ᰪ�P�57G�2
��E��Sj��ћ������� �K����w�)�>r���鑿?u�ʺ����n�+�����V�t�ᩳ�,Z7�a���䐘��C����^���0��W7�ȃ!6s�9_������#�̱��Ri�nm��~j��ڥ�kZݶ+��
�h7"L�@#ۢ4 �)6��H�	�	m�>��X���)�Bew�����``�̗��N�r�o2VF�F�W3#g���xS�a$�x�A������QV��5�1E�y��pbz��h� �V�U_1�&jU�\�*	��H$�]�9T"=ĹJ�>gצ�I�L]�Դ\y~��M��\Ű�~f-�����1��4�5l6�-9�H_�?Bt��Ŵ�f��"1��٭����=�v����}���<�u}2��6�q@4��J�#2�F��U����4��q�J��d-�:��:Z�6��Q5�N���5=��5�LB��{�;���9rO�!�_�"ؾ���+�A���o�j�j�}g��G�=���u]E듆ڟ��0��#%o��Q"t�:g��~�1���r��w���a�E)����cҰ8#~=W��tdM�_`[L0�8�9��}�3����Y��~��RJ
&{!L�A�D,Cb�'Cc_J	�3*�j,��#d�a��W��:d�%'���'�����_>x��];���اӠ�(�{�;#г�����3O�<���z������ߓk���v���"�g�|�@=raq.����<�����믳SW�����Z]��/�/v�D�R��w���rc|v{G��!#l�M����)��y�ψ��|�QG���o.�8S�$�]��H�E������~/ڽv�����\ݩBS>��J$P��Z�sh���k C�>6���Z�j�mT��W�8c���G](�ɔwl�i�l�b�aU��:��"�~���Y�< [�
A�R�Z(�i5��\+��5�2o'�'��h3t,���أ_9��1�*�a����o{���㉋������n83��s8��Tc�����:־7q~��������g�#"C��	𔚭�}�1j���9��=/ڬpl��~za_�(?�ȝ��U���׋���^S��p�����0���bH��5�i+��QtzL�{_L�L�	@y ���4>�A*��S��Cd�\89I�-2\_���P��X2Zovzio���j��i �m�����H�>��Q�x��l!������h��d�uxb����o9�%J�NA$��,14F������$4�&����J�f��0�g��G�7����Э1x���L��M��m��
��ۻ�@ߦn]<���?����~�w��?��а��mnKsD��X[4�$��)��aU�-8F��4��Tl��H���5���K�ݟ$�q��Ezg�+7��n�	3������|e+�IO����'jQd�j7u���]7�ڵs7���ڶ�z�I�c05�Y������Qjڦc؈m�3Zq�w(�$)���o��4�n�+�\�ҪSz�cPFͤ�����f=�H��*�)eZM�~�#e*���\ԭ�cm}�����*��΂=�3�>Վ��yR����7m�if�D�O�����5Fv[��]_Dt��%�@9�R7�{Y<����E��Q6�5Oo2qc���Z�뭁{:M��ꖰg4o�ii[�:��k4u<��D鳴�Y��qR6u����x-�{��9*���)���1=�s�����ڽ�g����<1<�%W���I�uCf��|�s�·#h;��j�t�jΥ�	�	���䱽N'R��W$R+AƻM�д���[���� �9n��)�G1K��l�"�� ��tb0imTG���J3�9�i2_�ǯ�NU
B~�ʔFYO¢�5{�Li�u"�a�O:��+0ͮ�u�lj�^�*+�2��C��[`��Q�=j���u�#K�gTnL�����Y����0�X�7�7�?3�q��~����A�K�~\��7�OO���O��{��Wv�~xnb����kK���Wz��;�[ڛ��V�So>LD5Z�f-/��h��ǿ��T�X��Cݵ���"�z�@��<H&|��v"R��ǘ�\Y5@�mDi��2Y7T�Dc�~�� �L}����xIA�`���?y��OF�id)K��:�ަPa+;����{N���s]�m�7EՒ��=F��A���m�j�=5�F�;q88iӯ�k�rvn���|k��NP5&�ހ�,�*t�e�~{S�F��^��AK^��=��U��`I�3�`�����N�5`�O�&i�s}��F6R���S 9�@��:�0�18b��5b�6/�P�n���[���u@d�G����2C��x6���ä=�a�c�!�M�h!_��pb���V�t$πs�l��9�C E���7?�(��{k�FŵK��s=�k��ʂ77#�Qdc�	����5������h����P�f�����έ��;z�ŗ$)��:�6]F��Έ)���s�YL[���8�=����k�YS_^���9��-�q�U�k����&�6m<������i�677�o��ß� �o�\Ӡ�U����
�?�7������Mܺ�;75�1==޽0=�ie~z��������kK�����ז�������%�nTF��WA��	�d��Nʽ�B9�\����ʫc�e�N��U�v�J�Q��F���.^�i^_g�6��٤b��)�Y���&�a��4:s�-7�˴8��m9���-������ ���Ǻ���.��U�h'����>f!Q>��֏�����h
�����C����g�3��C�&=j����
�%en�?S�"��51pN+򩞗B?�X��l�時��k�����)t�c���0�P�ᴄZ���tĉg�Т�y�C2�$�(�i��W|�f�@k�u��b-�Gg���ڼ$��NF�S��[L�3����ԕ&�] +aO��z�k�S�T��)��i}��5pC��M���wM�����y�~}֎�1��p�1%-3��a?�p����zR�-��M{��羱��s֖�*&�����F��Vᡑ��`�'��8W��]����V�q�� �h�v��IXDrXiV�7;7E	dW�2i}��N�u��Y#+!n�I�|H<��Y���Οƻ�5�Xz���M5{�:�,�vZ��|��}��o��������y�}���Nm�i��)d�}�6xȈ�gD!nO�����B���L���L���d���D���L��������-�h���<�d-���@]}��V� ����$��_��.5}j��2�\%����fZG�����#��è�]�pm���m���q���/2��R�`9N���s#��Ei�n�d�xW��V��|�J��]Ӧ��(Ԥ]#��X%j6:����:2�M�j��ػ8���q��3��Z�W7��D����/$��׀�Y7w��������榔���"9�iЊ���c�fȭN�kd|��1YT��Sqm�g&C궴,uC�Rʴ8��*Wk�k��uz�p���/�G_<Ƶ�&����;�nd���D�5�7�s�1W|��J���'�5��?k�3�O"��1�e@N��b����4�Ό�����*7�n��q�/�������<t�{%J:j���k�NU�V�5��s��)C�8��=UB��*��x��'����:Q:1���jL�z���F�N�d�9�g�G��wp|g��`�ްZ�j�!t~Kωt���U��lE-N��X�b�itbׅ����K|��)VԐ�1���ղW��E8�cE����{��������&ޖM��&i�?@��r�ݽ���(�U���g69|���mi�V��䭾���-�ej���Fn�>�8?����U��+uDq��D>l����[� �e`k�hJ�~}06��D�A�ia7�ÇG��ѵ�^eu�m9�N=�ӍO�sg/������v�ptETxψ���#&�� E��a�[�Ƽ��0Ƭ�;�����:Q�%���	��^���y:"�Ga%w9錍xdl$DTJx^�mPㆁt�
�8��5�
&��ip��K$�n:Ң��?;#�Ԫ�U4T���a�m�jl#j#U=ɱ�o���i�{�`�+ƣ�=7��$m�TH����^��GÑ�� �>���O�뢵�����Q"�@K�+ur�8_J����k�r�ƈ*ej����u���L2�J}�q?�_�~����S�ܱcT{�7�._��`�Z��ԳY��)JL��#R�J����<2��(n�H�%T�pr�c;���zY"����G���m2�'�Z��-.U���6ʇu1�'��P�j\���0Ў���Հ�R��G�Bd�����|^z�t�?��߉���+N��O~�S8itG�|U����Ǯ�$���H���)�[�Xlnoi��z�Б#��3_���0�z��x��A�������l�k c��_#|��q����2r���&�'�x��W����+1��8_F�ґ��9�I%RMR�u�5T�U��&g�p�]��Vn��N:њ�'�xڲ�sw�(��ׁ'*��Z����B5��1�ەg�KC�N�e�ۻZ��ڹF��֊�%R���j�=7�\D�����%���sS�G�#�k��y8j�1��k<���~�q]��M'�������qp����`��![}��EO���pe���H}�w��u}=�Q�m�646�ź<W�t����yP�9�0�؛��hf�,w ����	��L�j�C�'��$�Z�#�%�N9���qHƃ f}جE�Y8�o��ڴ��{K�q�F�:"���ǵ��4�f��
Z�2�f��u
y�_g@�Q��� �.E�n�[�X����<n����v�����[�!Lr�UҜ�m��̭���Pg�e'��8?r�W#5o�d�����&"~�{��{�蹏����=_�?�y��+[(')��V��4���t0�#[��a�`#�+�n_ơx����y&$ҏ�z�L�?~����;w�����/W������dޣ+L���0�����[�͟�z���l�����C��::9�K�1eɶ��]{+�v�(V�;�!W�t���,�Q�uC7P��52��M1ʆ��UYG�/�:��Ͽ��R���%�i�4F���$wi45�i�8����x��-Q��Xc@���7�^f��)�f�mQ�I5��[�W�|an:ƹ�ۻ-�BQҐ)��Z�������0�%����+Q#�e��ڴ� ǖ�8q�����	��v�y�����T�� �7�=�*��1�۷m��or�s3(��/"fJ$:.j����@��Ƭᰕ�kҁ ��a�m�̀�������krrCI���\K'�ӥ���	�Ҝ�]�tꮓ�P�W7�ض�i�m�&/^�@<�5v�%\�Z�4�-^S8q>!>��2Ad�
ډ��
k1��i_8��y�h_š1[����63d��c�Hʳ��{����eF$O��sf ��
!nN�9����"ێæ�ҽL'�� K��ޙ��=8_�W��� j����I}�қ��l�gO�4�,�))L��z�O�E��������	wbr��=E�1oi��6(����9�a��/�>�~��������ߞ<@�ف��u'�_�k�Ӷ�b4�lU�b�!B�w��^6�H#b�e�ٽ/"�[�02��������+D������ �ᅮ�lr�����i`���f��Lm�U��1��:"�j����Ij~��<�9�ĈI���r�������c~E�p�~s7�2�M��?�v=Fמ�ן����
�ΈmdT�Ú��F��!��<�kg^���~2NE�@���gl�{�N W�(�V��� ���QkI�Г�)��H9� �[���~r��l{#�]�i:H�-�i�]��Z�CA��D�X�ێ����~�g�#���N+Q��(Ư�A4�^;G�^!�n���#j�^I�;��Ժ-fN�k�La$��{�:o�g�߈�d������
ID�:��6Ԛ�gK�t�����w�ERf|�6��Ʌ\a�C�FTi\�)�P��&����(�VPi����|8k[Z#�1��ُ&@�L�f�i�B"��#&�E��'?�	��/}�KEٍ/���V�ʏp|^i�^7~7�w�ӠߍW-�����#��&~����W��hk�����.ףHeF?�x��,#c�=�P��@;V�Mz�6c8���݆���`�FI�: e���$B?Kf�s���Q�5�+g��ma(GG1�u�(^C��Ո�g�p
s(")����#$�q������(H����:;~��ǟ9�Z�;��^8��Ȅ:�0�j5�&�k�#3PmO;���V�n���)-X_�E3�v���jnŬϠ71Ƥ9"�����V��d��ǎ�q�?�G�|���Ԉ��a6m��V�.FJܑ�=��ci�0��'Go�u{�r	��,������8���n4�bY�Ѫ���=��-U�)x-4��7��(���k��M-Ł�,c�Z5fs�:Q:zF�:}D�W�]��>�%M��,鬴��R�fx<�%�����W�E>F��6�}�tL$1�xLE-�8{�`���M�gb'��t��"e���R҂�A�q��έuz��}���͘_�΃:�־;��۶نùe˶�p��{.�zțO ��կ~G�`h�[�7����y��eiO`�!���B �;�l��]�@�Sn4�/�|�w�u�?~�莐�d#�\$CW�
����'�Rf��
��H�o'v��6E9<t�2ID��v�3yU/R�J����ɮ�֨��K�;u�ԝ�5m�ԍ=���4{̮���k$��i����G�f�)ZSަ�%b�'j>K[���}��Z�W���<C*��{��z��=䞛ji�і��F�>/�A�)n����6
ڮL�ߞ(#Y��z�L��7`�^kOs`�
�&��_�����g�ވ�`�;2���ipF�[�D8��hu�b�s[�T峧�2�����{C�#sq������m�	�V$�Ŝy���`[��XǄ8]��"��(R_�
�圛d5��h����"Q��p#dC}��֩���[;w&��W�]�p��g"�=�1W@Gg�T�xY���4�����G:y�6��;���2�Zi�㾂h�}�2b�v�7�w,�Vvv�T���X'�ܳ�,��
�e���H��9�����8r�ѐ�Ձ���Գ�$c������U:^�k6��t�i�����~g��|���30�w8��������(�/�lI���F��MN-p�Ѫ�ޅ�O"�uQ'l}�� 	{,�B��M[��K6�'�$?O��1ٍe:��j���k��0*�v,#<�D����fl-3��}3H_#�_��_�h���/D�x'2�m�F�E�SCk��2lӬ���Qs��S�4���ù�=F����mVCC5c���COf�'1D�Λ�V�sB�Z�r�bZ����6���{��0��݅4'K^����%: ���B����Q���Se��P�	�`,nܸe��l)3#�����m� ��:,u�m��8���G:ש�"��/�"(��u��3�����s�'�� �5��L��vM�;�T�E�5�t$=w��3�p���K���u�d��?K&�ɾ��@i���2E���Qr;���N(�"/sZ�J��@_�q��UF����/S&z��#�~����*��/f����ɠ��V����~+���ڼ��-q���s�����H���B"�& ��"y���C��)��+Q�.��)�/|���|>Py���}2��jO��8jr�E�����T�y�G�tI`5��F/z���y��Ն7E���i��z���Q72�I�=�E�1�k�M��כ�5�,J]��-��g~�� �}�#	����W�����{̜��:�����Ā��G�������Z�L��L	� ���k��I��l�0B�N���l��`���m�������C�FŵY�0B��._�h4��8cd.\W�#�p}4.:�|��m����%��a���l}Z��~��:DN����ƿ��1�S�	U=�?D�ez�3۬'�"[޴��J���Q�n�k�^v�	P��,��q������!@��({�ѭ�s��.�7Gv��螻ٖ �� ����f���iR�7Ȑ՚�J�{D�M�M'!��C����6{�u�y���Le�v�a��ѹ1�^�iJ%�#�3�3�Ce��}�^w������߈�A6��%ֹΕ����	��X�lWOo�����6�;p��݅@[[��K/?�g�C��>�=?��ZD��d1*�lkHBۉ�e�K���lTb&;��~��^�HA
m��M��Ncl]�uz�M��i�R�ĸؠ����T�l�h�h��Մ`4��c��N�F���' �I�{��G��\'�5���k�#M��v~����Ԫ�!�/a���������nlD�c��|��o���'_�)��~�guN�0]X���8'�^�oh�_�,_1��O�c�R��Q�x�����28�.��1{^E6ۥ�3Ű�~VH�:�
�g�ر�#���@�U#3Jy�b\��t�ˇА�MQ;L﷑��H�'��>�%5
��s.�n}��?j�3�4e$A^��̬������̏9���[�Lh�g���	�)o�+O��sQ|�2����;`�5ϫ("��5���p$� 0�:{`Q��P7w<*���V"{�m��DeO�@����<F�҅�ܬ�e�w���+S�:�����!����
�WKD�e-d��������iP¸����$NGyB>�1Ҡ�c��߭�v�@$�'��c;��t cSG4e���&���(xÆ����{h�TƲFy%�xP�d\ �3�lt�ߊ��*��聖Dd뗏Z�}63Ѭ�5�i�H��l�e��_5�����t��k���%B|�:_���?�'�˦}��J[�Jl��q0҆�N�2��r8(׷�ɮ6��'��G4�!��]㽡k�q��n4k۞)wyf�Q�m1��X�1E���~�uW�׾�z"��*�l��_�D�<G���Hic�I�0�6?8x-��֍��	���B�X�E�A��6���ӂ6���hi_�(�S��L�$���*Ѿ�I���mQW#u9J�޸v��ʖ����2�l׮���h�o��5n��.��TУ�������'6+�S�8'��q�t�p�4���!쀜Ќg�t9}�5/�5�3z����<YHr���e{٢%�R�I�\�Չ������fj��3���Zy�ٟ��e��[����={����ű��ͺ��y���ſ�Џƿ�N�ߙ����޳�ջu?��֝�n�Z��w�M;����7��l�De�bl{v2�L��xD�lh��d����FT"F(��p�Ce0L-�-S�L�J&s����<�3�M��Ѹ�]l[��b&�qX5B�Ƚ�1�$�+��b�U"�{9[����a������[�"��#Z���������(Aؚkhl~���O))LRz���9s���.���7nܴ�c���>��d���� �3m�S��:j鍝��q�f$6Sb�#����9l�<�:4��B����S�KY�2��#��7�7%=MTކ���䘫��X��<?&��m�����MM� pv���<��<��,�um��W����VB��PQ�CF��Q�c )&"� ��P*��t�0�@b�F�`�����s����/��{�}>������� ���s�ˆ�_��,�#�����ػ�+#��U�?��r�X�G}sU	�Q��M���I�0x���Wwp}ih�=
��L�*\h�C[�c��9���`�o~����7#�4��o�781t6(�]��O����s���ޛ����"��'�ܗ�i�R�~L�R��+^���A�\$� �D�)��mb^_��1t /�+��q�W'���>��rór��!�H���������1W��� ,��e���<��io���L7q����Qs�{�3
�������7-!�ʆ1��tz��T��[ĳH !9�nwx�I֯:ُb��퇬�?�.s���O���ᖴ����P2�x�r�Q�uq�$޾A��PI 9YL�'G����~~!碠d"��L�͇>����w8a0J�������84� ���2����͙G��Q�\�b[QD�כk��?�n����6�P�������F!ӏ
�laT"���u���da*k�l���-׶�Ns�Б�ب��
P�o��.���C!(�IҜ����Á�z�W��lEI޵zBׅ��(ns��V�1O偰Z���	�i��p�.�>�4�פoi������t�Ӂ}⸔eN�΋�utk-��"&�p�;{�9�����R�q�=���C͝ �:�h6׆��A�f̤����_4��5p�2V�U�z�#"~�:(bo�B���9�c���X��V_���.;ZW����\�ظ8�S����(�w}�ϕZ�ʌ�e�S�דcCi������3�<�լ�q�ʼ����b��E���b��;��}PfK,�'E�}�[ǵ34�e�E��I�\���������17�>�~Q������뎷���q�X����3��e��G��{/�Ȗ)��ه�"����x���z�mQPp~�>~��M�>`z��EU8�$����a���h���uZE[i��q	�ؓ�әAֳ�,��7�%q�q������	�A!!!�S��W���,u?��+�� hJ���2l�p�Q�	���w>����U]��yiQ��6�[�_�49�l~�]v�����	�ʺP���Y��Ÿ���s��N)m,M� �+��`SE֘vBd���W�yԋ��H�8Vv�Z�#	n��1��A�ʖ�ZQ��mNЩ6j�(㭶 �Y�R��3���ۖ�9�ُc�����╵S���L��V��|���4f\�����.�eى��BC�f*�fZ[ׄ�I��~z��gL�ɹ����ͯټ�E3���/ww����^T ��CW����xoW��M��b���v�몾r��E�X,���$�9r�B�Rk>�����8�*~Ln�R^m��j��8��X]j��mՉ���pB���#.}M�iV����Zτw����� ƅ��2�N_������K�+
si�����ഖ��g�����=�|sUJ��e�}X�h��N[y��?w����w�wo�V�"�ź�]��t����	W������X��������m[�ŢN2%�KH���u%,����?�~���LRn��mB�Z��<��k/��p#��>�v�V*:bL��� @�w�v"߶�E�N���(�n*:�:w
+�\�LCV�7�>o�@��7zQ\�WqWL���'�-h���c�²M��C�d(|�X����A���0VM���ޞ��U�0K��C`�)&21D�R^E@�;��L�'�n8���k��^/�4�(ͻ��fS��>'h��j[��b�/�C�>Z%߮�R3�	�P`��:z���������M�P`��џVg�����sh�%����/���r�[Ö�b�-�O�R�a#@w��<K�%0���&��ֈ�`�Zs� �-��=���ϡ�?�>���+8�D�Ҳ�c�D=�wo�IBKvs�8ԝ,���+�!7���N��T�D�rď�����+*�c,���c�n0��ԻG��M���RM����{j.ʈ1?K.��W-��g��d��j�td��`�&BN�� z�����]��]t9�Ӈ����?	 �����b�Ct!�-�&lO3Oh\,Q<��,��_xF&r�]�"���bYc1?���ŝ�w�+�5��������N���n~�}��hU�#_Ͱw�\J*��P@��]��w��;�KA���J�e���̶��"s���!3ͨ�eK�vN �Gess֧�-ӡo����
�8�VW��;�&�_�3�VJ8m�bڋP'���2��U�SJ�A�GS۷>Oߟ6�_䰫]6込%�c���Vq����{P��������N^���uL��ܳ�������L��z8�� ����%�!=c���ݚ�hg[<�w�9���|"��;�ޕ7�\�e:F�y�-�� ���x{�[��EQ͝�]/�8�o�������5��Zļ{�ķ#��_N������g̟R��v��y�d,]ғ���)�%'�g��wjS8\��_$�`�������\�p���e #r��+qD���M�u>1%=��H�9YRlZ���EMf���`�e��d1�2Y{���&��/%Ә��q��u�*[�t�JC�z#܆�J�2��|��31�Hn��Ԛ�{�Y��O<�~���d.��6�,`���,�&O�{Ќ1��<��$�W���9�N�ࠑ0qRp�Qu��t�rR�%�h�(����~�����ь��]��xUN:�z߁T�(�+Ϛ@ۊh�d����]�)�Po�ݹ�����u����;8la2*�C��۸[���e1�-Q��{�`<�5|���G�3���?����l�k#�N���!܇͋«�XKz��l���Pޮ?c�ٽ$���g�χ뒊vt�_[+�z޴�:�@�1T��AX�ނ���h�pZ��d��Y�Gj��jfK�;DV+��%��T��)/r�hŞh)������D����C��+�L����]�jJm��t���i"ZIo�	�=!'�wd�MFu��^�FC/���Bk��+��YU�o�M��PDɮ�� q[X�D�����ɵs���+ب+<��~���V� ����@���ߴ�y[q^r\kr�6��0�!����ױ�����&�z��^eg���D�o=���[1��%��v�dCűO�`nM?P��s��y���'��"&k}�a*��u���s/��"/�ē	��ڷ���-��B�y.�>�Tl�q&��V�����Ac?B�uS��-c���9�41��4|�'��,�[�ݻ�\ۇ=�G"���Po���s����T���r��Ǥ�0kU���������+M�	(5x���UMg$�%E'2�rC������k�b�ҟC�rD�p�D����Ĥgs@���O�,��v���~�#@KH%���:�����ޥ�)���~)������I�oK�(�A�c�������,�(���8�qgJ���b:G(y��H0���z�\n��M��`ga/U^/�8:� ��=��x M�.��D�i����-[�y�ٟ30L^�	�u��hQc�J(XK���u�I5Wj��.���t��|*`��n�or5�e��.���=Y-}�j��ծ��ݿ�7CuW�V�9�ڪӴ�~.�!y�� �6�Ɛ�`7����^+g Z!�յ����S�A�2�5���pa׮3��T=��H}��}��[P�����m���&-!R��R�P�:�'�2?5�r�7mR�����l�Lw��%o�ʗ�- �j�I��C}'�B�1=�2��L��E~��yXz�S��!<U2����a5�_� �>�Y&)�0�R�f�G�pM�4��s�8�£I�Ʒ��Ы�#�o��Kgz��AÍ8��z��D�k=�^���E��u���5Əύd�s,���\W1A�G�7�2�]��fC;"&�#��PH>��x���;0�_-�m5U�4�*NL�Y� ���,�P�߃J����C�C�֮�g���Lj�1���U�u6�ֻ��򀌴�;,���7������f�l�K�d�S����S��R���OrF�C5���hy����wr����)'ɖ�2�,9	(�r
�: >Mc��	����)�@+�xx_�`������2-ʧ� �3�nx�4ᤰK�׎�;�٭���i	��L'A�/&5VݪGv�[�d'5Vh����ƫ��φ/C�!�����0�H����$aޝ�ؓu���H�,t���O,+�D���
,z��	���d�Z��ژx����?�*���8���&zZ	9��눈���k�[J�c��654M>��֊{����!T�$!AO�f�(��{4M�� �[ᭈ����R��u��oX����9ݗ3�`˴yl�K������
>\���X��\;�N��33y6^��tC���Ή�C!�2�2��Z;��J���`��ߵ��I��G(�P���svZ��GT�{���8��H�?S����W��e���l��ky�Jq!����ʹ!̬��s�jA�V�8�b���m�Ԥ�f�F&WSm
�9���|�b�1�=�Ł�`.|�,-�4�"��߂�b�h!��r�� ^~���67�U�Q���h!�[�2s����L���Y��j^,o�hP�FP���#�ğ��:*���h{;��a-AVE�����;>��fOop�5ƿ&����K�N��0��\�\W�,�|ݟ4�H�E	��`/��r[Uj�X��/=�VJrW����2�'���O��R�T�����%�u��xt1{|�U�;�Ã!�V ���˒�����*ݚ�'z�#�^&����yج��n�<�7��>��-{��e���I�Y���}>�Gؚ%#Q����`�]^�J�;�2�������w��,W��S=��ۇta�&��3y�Ѩ�E1l�R��Pu8ٛ#BJ���"�bI�ɝ���f�J?>����-}�sX�I&�Y�p�����a�a>8[0����|c{ �/�H�=Tm�|,���A{
��N4{nLV���+Lo'���!���UKu��!-?���(���6����5ү�pB���U3�*4��ܨ�����{� �"���]�U�DR��fA�q$$�������q�%���M��jG��Iӛf���Ϸs������[h(��p��قT���P2�9 �z@w#z0���ny���6DE��Lf5{<�"賈���m���K\A�U�Z����w ��Æ�@�WON˙aٔ��P�K��t/��?�M��.&��*���!;$-��m���̓��
:\ڃX����$���mp���ꀩ5����`�ҥ8�6���<�O@�,j�:xk)����k6GS���@�ɴ_j���;[m�SG������q[��<�r�+Q6��*~&G�	ym�a}/CҠ��N]u��82�F�����l��Cy�p�OdK��� �O�xr$��TxWQ0��L!�f9}G�{��F�(*#ɭA��)"1I���t������)��`�Z�?�7E�:��e��R6b��L{���w��`��`l�}m��!��HK)E=�O��O&�����E/��[vA�Z[��4�<���kT��QS�\��h]�]�Jo��VWeG+A�	�
��+�;�\	�U�F����L���8�����Lz���wk{�қ�Q�38"d��hS/���W)�4�	�0�`�e�]1lo�$>S1>Prl��]�k�7��~�}��7[�Ѕn׾z�b ��,:� ���-�n�B�Gjg~�}�+f���a��\=�d������pI�T�jO&�j����{�D���=Duu=m�lk�ۜ6P��|X���C��)Y_�}��f��D�}\ʶ�y/�QF'n�	<���.�s��m���J�$w����7$%%����?M��B"���xr9W=����D u�m�5�c2>��޸�ȿ������������qz��)��^S�kWW���� X��.�� PK   �cW]*�Ļ� �� /   images/5241023b-b430-49fc-8631-1e6053993f23.png��UP^�%<�;��w��$�M��	�:�Kpgp<8�!@pw���n����pnUWW��>}��n��'%<lJl  ���,�  � Ȝ����td�  ���rrZ*rr�Zn�6�߭ ���L-]���c<d�"e�.g���id6e�wX���!�rV�HK����<�lmd���l-
����٠}�����ڞ�^_��"ޓ������� RM��_ �h��m$���6' a0�Y��<*" _~�	�u���E�����fM` ��D�LL�>���1�R�:�:�w�GD[�3��&GR%'cH��I����Ï[#�� ~���#��"�-!�����S���H�J��r�T��Ҝ��#����#�̜>n�$��o��f}�^�v )�<���{��f�ş��*c�_�E]?�ơ� H�p�s,��Y�b�$!f��7b�t�9v�\+�����g�]Ut��c}g�=���cTE�3�)ۋ��t��Ɉ$����\]��n� b�l�@��D_�DX���~{oz >����xU3��L/9���n�\jW3��>�̡�ޝ�c�S�}�4���g����=	�*��J�$�޹�������n��b���rV�1ďensq)��/�ߙ������?�RV���e�+`BP�TВ]��0���o^�X��>3����s<�M=�d/��!��L�(8Ht���L׃fb�x���˘-��Zxw�([�E�s��]h���z5\�%Qݦ	����h�?����͆��[�#n������!��E�`��PF�Z�-Ӣ��:9)4-L��=Gۈ�+�p�wC��g���e��]qyO�����%J��4��/ �)tj`i���:+�nQx����,6[a�$EKg^U���s��ls��V���<�		e\yQ�g��8!M�AI�4�t:���C.��\*Yd�ė�V��$Ne�k��|��9�$+.�#+hܟ�l�7�¤>dY�;���k�?�Z��@▋�F�$
y��B�Y�\[c�Q[к�$V]T�����E R75��	�c��B���AV_uYvYɎy���D1�C^��/%K�X��^�������̄��iϣ"?���G��T?�J+�(I0c�+���S���B�*��P���.����n×��/�م�7t��Ե���p��M��|�.��V-��ӣ�dn��K�K/���[��A���~���ʘJp�l��g�	ڂ4e�����C�PS`S\S�x�����q����'x}NeN�a�*q3G�z�y��,�[%������E~����ܷ���B�̔	��B�@~��9A{a���G���Ăau��xq�{O�L�,�8�S�4����mV���+}e�U*n49���#�d$��;�b�TNAE��sܦA��Kn�d�Y�@�m�-ʭ5��F�V	O������ R%�w7*�&ކ�[�R��L��E�[g���3bˆ�ҕ��_��K�SM�7���c\c�C��b�y�6�s��h߷��-��]�[<ZHΛNsb���u%m�8ެq,UnV.��X��m|�ǲi��5!bĺ��Bp�wz�}jx��l�|}Vuz!�E�L�E�I�ӫɃT���ԵXl��:p��2hp��%yd����0�O7�mYci�5�o�u�ڇ�L�p��\3=�rn�����g�kv��
���L�ZO=��j_�=/�����;q<���Қ�6�D-�|,�f�vY�=��F�f����J�|�{N}��D��!g����EE�p��^ؾj�\ߦ�,|��oo+zkt��ٻ��+��\[�KI%�
1�p79�(i|�1�'O/����������(o�i2�x�c��wW�ii\�܆b~A&7Qo!Yo}�5Nc������m>����${|�o��sL{�C�C�qj����a7�
�
�����0H�a}�:��v��KG�$��lq/3�%��GQ�U�V�J�Ja%(�)K���-V����Ο���?��Z�R	�(�(X+w]�˝R�yb�J����Vs���2m�Vp�܎�-=LlX�>,�B��ҟ\]ov,��2�3�M~7���6�Ʀ��V3���]��h���ӣ��p���=�"�'S��&�x�ւf�v���ڞ{�}�����V����~���X�e��n\.��l%�0���6{5�}��"��u5-����N.��@F��{�:�Q�ѫQ����zSD{��XGM\�7vo��M�u�5�:�_v+NM��w�����U���vl���f�5&�����jU2dg�+$���J�x���7m���=����_�Z��A�A�!0�3OOO�f��QP�۰��?���.ja�
-��\��y�z<��W��=���./iX�XUs
��4&�'�2�2jS?��ni>;�@����OU��.�>����F�C���IV��h���4B��}M�ݴ3`�u6�kxe�6S�ĵ���p-t�Xʯ?L���O�k�;5�{t��
UAǹ���6�=��W7ļ;����?��a� ����ކ�c�\әӦK�K�_J��!T��Ws]�]K`E�����G�;:S8X� ��o^��0�����MU�%�y�uu��զ.�u�e�v{y�4�d�ص���ђ\��z!�������u�"q���H�����h�5��*YRXZ���`�@beF��� �Dv"H������9�Y�0�O�a�-� ���.X�PI$�A�b�2�m��?�o�����n�B�+�>���E��Y�����
Q���M�'s���B�v���  �z>�N_�S��|7c
���s�#|i���bN�+�dl,�&8u� \.���T�%43`�M�����#�&�+�ff��4k�E��by<R�Dz��,툜*~��K�{�)1N���qTl��
�����U`�m����Yϝ���?l1� Kѵ�n��^���B�7�`\�B��LLh6��O�����[$������Fһ�ץ	�=��MA�������� ��i��v�y �|�q988���#o�������It D�Ĺ�n�Y��a7�tő�>ĥ�����<M����/��$�	�Ȁ`Ϗ�Q<&<�G�9����b빉�A�l�����uo��,:�7$P�o/Y	�U��(�u��n5^�5�"�_���?������h'AdS>�YG��y�0�]�,��>O��K%󩯨��1�����t���St������,++S�~�988���qv������#��l� ��OLka��S����FJ��"=�~���
�|qϊ&�ދz����

{,L#���^<�t��%w���,��{��+tR��
U^vVV����*�+y����I��X��?t@��2�Q�-�<���
��~��Na�^�����LceK�M'��|���l�Bv�����F|����i�z��D)i�BNN�%Z�n��9�@��GM���Q�T���y���>�%�&��w��a�~�'#q��,`H���3@���-E/�����}z�����Ȱ���.Rl���ڍQw��Z9d�If�
NW�޽@}H������?I�yM�0��<6��a	z�6u+MH=��^w%剹���SB��v�/3~5
��.�W��a��^��E���ʽ!qH�}��uji�\�l�K_?���8&�0n�Li2���s6k�{��p��B.WVV�#""��E#E*�8����Y��TK��;��+�s=$�l�I)��#�2�,�%hܽP�	�>B剱^�C��C��Ł��L���2I��s[@�H*�����;��kV���(:����	B6���k����B�������8ɟY������X����u	y���E�<oCR��J~N��bXuS�^��2���Q��{^�S�$�`j%�=�&�o��3�%˭�f���G�O�5@�����*����X!F�A2���vu]n��`(+�k����`	��'
��@��:�-��2�jP�z	�~��M�w�z��ҿ���E�K[��)���x(P��<m�='v?���5�I=\����<"'�\Kp��1��F�pO|��!D�E���j���0S�@�F"�;�$VMt��l��^����5}�5%P��e�	�9<k^�?��c�ܵ_�Tˎd*���� H�쳈�F�ވbW_����3��K?uc��M ���о+M$h��������0�C���C�i�q�6���ż�M[�F�*P�.i ��j�O̼Q;D)h{�XfV҂��n������I1���OO��	�����v�+j�Uz�֖a���8�s�p�du�i`3�866�
����sL:�a��g�����cD=� ��]ƣ�xHB���PF0��Keu�����h6c�.����'*�Y =�nY�I���~-}b�mӅ�����p��]P��;{sβb�4|�py[��i�3&�ZӪXn��S��o���Lz�����"�Mp2�$��h��X����t�����ܻG�a˫3b��y4	q,�R1F�{{��{ZI����z���&�����������8Z|5�������(� }t;	l�K�r�>�.��'t����<��8��T/��e�M�샗�#�W���1�E0��-�	�p��ǚ���v�g������m�\�*0E4���.Z�+����@��3p��*�?�䝗��iG�'�`i&�-��a��C��xz2�\;o�FKd�S��&��M�Ď��+�?=jHr ��r��`]��H���Yy�!�HyPLrs��ϕy���9C\i^�C'��]cA���N5�o&� �B�Q������M�S���+8�͵�{�b���5��V�c�oI%;3�e	�R�_9�����m��]�B`�)�B���A�j�2�m��6����j����B<0�},{;=H�i�h�Z{yNSN�2��ߵa�m�0���-������o���ZX�*D�LM����a)������=&d��9�\�&��-ŖUp��	6��oO72�	^��4XR�C6����bg�$zy1P�#8��V-�a�Ð�W�y{�9[��Dx�*s�>�5�Y�4�%����/��0=�.	(����".d(�P�|�)��n�` ���T����z����YR��'jڑt����9��ݯK_�ø��\TS�pL1��(��)����Z�=^r+,�CK��d<��˓S�{�Ḁ�f�f����=¿=��0*%9*���!$L��������%m��7��D`?���TNs�@q����!N�A_�#�S�:y��S^�����B'������yh�T׶�9Y��6�e��������R�;����h!
�,=�㋏����ҧ#vQ.Ruf��Z�/�C�3�_�w�*\M!)?u�Q�1�D�
��D�c빹+�)�:ߪ-����C�����n��#�r3zNB����֟��e����!��|���XsJ��l�'��+gd�2����N�l���:�0����b�����'�h�6O����9�E�_E���$ xg�@��:����#	�[)c޵�Ru���כ���l�nz����~�"K~IAR,0 �2��Y7�a�'�6��6!!}���M�u�����FAA�&��.�-#��/h�j��D�`2-b�����+a��2���w��<��WU�/Te�!ߦ�A�^4�Lh·< `4�2���ueh¥�Y�[�������!���چ�ϰ��|i�9��v�����d �ov�"���B���f?�&�,݌���%_(-��ל��<i���m�TJ���_����gm�'��խ�?�o���|)�':�&��`�C1`]_��������y���J=?��ꚓ��5��G�����3G�#F�+F��q��3����b3�:NMm�Afq�`�эH����R�4Bq�" H��x/�T8ښ���g������]�����Ȓ�*��I��W�-OAN�4*���)aF��O
�UȲM��Cu���Ľ���2bH�R.���d�?#�trǛ/C�����-G{��O��O6�6��h����PE@�Bd˥�
���mb��|v&;=���"�]�yͨ�ټC�#��jx9]�ُ([��]s�����P�����x���p�v����AQ���k�O����].(��~Z��)�y��eq�0<��C����-z۶x�	M�����P�	��/K��h����	so���A����;�w��Nj�v��+KK��$��C6t����λ�t�Q�ݮ|�*�ݗ_A��cu�W8�O�w�M1������x@��r��w�B"a�Y�җr��������@��5`(=���E�۸:ԻDz�g䐾Od(��8�,R���O��f�0i/͢ �P�G�N�ԋĭb$��ϗD_ك��,� �@�9�eY�8�WG������ѫ����0htʉ��u|�Z����
��kW��SY0�Y�� =�S���ŭj�����1��b�O�m)'�MW&+ːS��-]�Ug#}�l��^Sq�31a�G��)ΝkZc�6�������x��a�{�����w����'�j�i�Ʌ fR�4t��u�	b��gX��[�mmeu�S�b�(��^0��1߭-��^6w�8�����V�o�)̆����or�.%P�:;��J"#2�+?
^a���� r��w�����D����q�G�x߂�����R#^���]/c�Q �s��:�;{�4���w�)�d�=C�m���ooh��|�;��]�T{ߤH�A�l��y�2'�kΰ�l�������4�7vV���=f����]Wq��<���ׇ���^]�7��̦@��s�{���gXKWi���M�*���M?w]���e�:G�]�z�e��c��F?��)�O��)򴯭7�d��4�Z��Y���n�s[NH�D"��˷
L��-t\��6�6nu���9\;L��Y�s2�M.��U٧+�g���L����$%2�	�j̷�r�!Z�89ګ�w#D	8��^�T�_�{�:Ԭ#������gH�U�r<2Q�s�_H�_݉�'}'mߍy���{#���yG�_5��P���HOH׾���{��/KϹP��/������+q��t�X���i�iu��Y�U��1�Z�-���O��:��}=�t�T��tY͵ck��b�H7<���N��5�:[�HCn�k|O���V>:&��i�g�ιL����РG�7��6R��Rs��?�pf��_�O�W����l��������n��~9sNP�˝�WE�M��B����0j�!M}�W'Anߌn���Е�+���_֜�g��+#w��_+Y+����������ȽQh0��A��)���i�`�1��Z�QC��ٳ�)ng����;�q���u��_�g&B�� ��\�{�N�Kk�� o9\�'C$�iq���۷G/�+�k�Wgs��,ݾ�Jx��Pg�#��M$¯���>�>��wp�n޳D\X�-U�k�FgC�JGwK�����svk��H������M+�דC��h��\���&���95w���$��(C��:�LY�j}��2�u�����Cgd�Y��w���f4)5�������v�L��B��V���Z x�%BGA�n�͞>u�{�7>��C�d��Fӈ7�3Tv��5Q�K(���x:��o�WdX����ݡ�4X��x|c醮�����m,���W|�u)ǫ�һf��M��R�sD�xb��_���<q�:?X���+hIVC⍤�j;ކ�4v��t��=�����5��%����L�������;'g�L�?A&�9ڨn�нB�96Z86�'����rij��b0��]�5�ݭ�w����������ӷ�-�RQ���G3����,SuMMr����j�ݥ���o�&�l��!1�ґ��b�z�����%|�����)º̢]�ڊ�Omޥ�Q�s��iB�湜�,$�td�|��؄m;^+aQ�&��9��W�	��l'�h�I��Ɖ��aAu�iL�'���M#�I�b�,1��=4�����pt̶�f�\���c#���:�!,�3wjb����1�[����9�D����\�.���S���qU�Hz�v����	�F�D�7��m�ϒ�2G�.V]���S%wo7�T5������I�,N:��5��f�"�,�#�r���������A�D��r޾MQd3u�
Fwoo�;v��R97O�x��?�^eJ����ߺFgCl�m#�0�H��w=���ZO��ADM�#,�e�c@��e��*s�~��Xb���W/����T��Sh�MCd}F}��T)x��>��l֙;�v��,��P�[ĸ�.@�6�G����-9���qUh���.���϶����V'/�X<|�{��"�-��20PXj���ň��$
�~f!���/"�bw�	-�9-J�+"���=����1$����t ;;�2�K���-����2�[�����C�k1��ø���AZNV{�_U���f�H���̥�����0�;	AMMm����Y&�a�T� �����=.DN�s�NH��Zʇ�Hw�N i�.�CC��ȧ�}�(���v <�R��W��-�
eud�~�
ҙ�{ڸ����̟P�7d(Ͽ,a���xkA-)����=M��M�����L�(��;Қ�z������/'�rO%C$��wȧ��U�9����6��Gz�v��ܡ�y��Ȅ(������	�k�]���+4ܨ�חp��]p�E#<���g���z@}"�C5��Y�����nuk]������z���\�ɜne^22C�A*-T³)���H���6!X���5I�V۳k[ƀx�U��_�
�!�v�#�/k��/D�N3���]�1wqq����B�K�iqG�-R��?r3:F��i!��Fp��ʓ�O&��p�����3��n�BzBiW�)�h��@F����n͗�57��

�
���qk�v�=#����x��%y.�^�&���m�D�Y�Km��>�X#Ņ�
��\WdduI#Z����m�Y,ED�(�R�(+v�X*�/
��?FwDx	�����$��v%KJ|���T���x5H�񮋀S*���B��bpϙܜ�\W��\�2�b`Y�#`���[ѲX����Mv9����i��a����*�T�z�?� ��S�&�&��4d����}W��Oy"Ǿ�4A������
�zy�4��\�0ڒ�ƒ�h��S�$]�yQ����B:���ůU���Pu@�0��k1���&�|G&"Y�#֍��04x2���A	֚�����$�4{xv�����R��V^jnvjGY9�Mf��9 '��E��k��C�RV�\���'1��I"�1\o�/e���_|�����J�FL�4D����`|�7qx[��+}=�T�U�+��K�9�9�]Ik��0�p����>{y��)�eg(T�J蘦��e�xゃ`��=��S����)e�]�M����)H��|$V�VX������)��Y��װ�"���A����r�;Q%�yF�rj�������rcl�V�N$v���`����t�q�"�T�9��l5��ږmQ0ġ�X}�O3�=�b��gbbB�.nLMM�W�Իwy�ޣ5i+��3���G�+�G�S�u�B�����թ��~-�/i6��Iϭ%c��`��\�� �n9NpU!O=�i~�k��w[��'�d�`ma�SJ����uw�qUper��!��Iy��?a�%�<���C�tz�w�)������'M\��o�=(Kn[߯Q�d�gb���4���'�R{�}ֵM��	�����I5��3IA���J�N�ػX��&�Bu`?� �#�-��E��G�Ly�c1�!Ѿ��⇮�`��r	 �͸�� %��
��}�F!ߪ6Z	�e��{�P�fgs\�$�b̹T����������9k�娇�&�óz9�
�0��!�]I�aIur"��}�>Y�Z����̓��c��������^ND�ʦ�L|�m��.��-�r��ͤ4rh��Q��7�
�th��Y�CH!��
�G�C��k�x��ůW�5�e�Y�W[@]��/�*���@���J���r(5H��+���-]�A��qll~]5~|�$��Z���i�f#�V�!�*�*��v�y��w�ǩp�PJ��*(�-+�[��6 ַ<�����T7�H���cK�8�p���z�;�~���������s�h��; ��C�� 0�ޑhJ~�Q���T!`Q2Y���n�\�)U�'"�4Q����n��-?F%��e�a knVu��ck�F����"/ўtꨋ�@��,yB���s�:D)$9�(V�<uVX�N=,�(u}�)�!�G|�l�����;<��v������x
�qB�S��
��T}����΂mD_H�廅����茔zj@YJ�:�BlGG�J�$�nm���8L�v�al�;<���P��(AвaV�c��W�P��o�a�F�Z�O�#w-'�]�^b��k o�R�2�"����75q2a���$�jV��]>�m@��N�2a�
7}�&���;Ri>oq�����F���5z�k�H��/�*+02����/�?�<BKC������0赲^;YT�T��~Q "�	0G�hj��,̸�s�&agAB�2����p�����׫�X��$�0�0u�A�x���v�nK�����z/LF�:!����X�)�����Z������Uǔ��o}�4�+����5�}��ZO�g5���߰`Run|i�2ϙ��e�b1�im6lu~-#Wr0h�dS���q�6t�,!�s�"�k�'g�N����ϟuV�#)��*z��m�jh��uBL$r�
'v�1 �3�ƟB��A��"�v���M�M�*O�3;4He�&����n�}�u�G*�<�c�P'T�"k'<��}�m��6���
��Q��EH���� ��!':xgt ���:��Y5��������I���1Tq���'�7�$�+e;v|�'����G/3}�DIZ.9\�'+.�Ҝ�6�gc��G4>ٰ�u���vMh���u���+���k���䫿=��\�du��[!��R�|
O�?�MԪ�M�}���j�װ���5;�P�Uc3�1z,͏�u��u�r$��T�c��M�]�=oR����n ��2��e6?d�:�ŗ?ow1�m2����zx]\�{~�^�~$�����z�g<�.!�����jJ����U���k�>_��i�_1�D�0�
�gs�ss�1�m,3��Pg*��j�Gf~�M.�2bTJjMd���t�,g����m�-'B&(W��Մ6���N2Y�V��d�r�]����o�����YA@7�����{����*1i.�5�li�7�Aߞ�t�^6����q��l.l��D�y��s���l%�+���B[�y��%M0۠:��
�]|>����wM#Jv����ô}^�&��(�f��������b���:�#_1�6e�e7wp~B����T�q-�-��q���[����RI�A�WUo��C�p�nY��VW��Y�R����,[�X� :�36uV��獮�]�=U+m�\sq����}w���Yee���S�d��U�ڥ(Jr/��3����oI����Rḋ�?.�"!Ii���3��)�ʔ"'����]՜�.gl��io� ��J�+���$b	�T瞐�Yî"���O�����AQr��y���b��%%�2En~�D��V�^LٙH�3Κ���l��Ly�n���N�ȧ��@GY��i����Z����e`���ݨ^���͆�����f�뭘]woI��$�M�1�V<�c���#�+��+���vĀ�G�Z������A��4ʹq��H����a�s�O���1�v�pś�y�	�ܗId��b���Tן�����+&J��
i����pԧǉ�PI��r2b�K��� ������i��UG����\�VZ(�m�
�?�ۦ����8\3-ܣ����%n~����Z�ܘ��Tc�`�
rИ}q�	�pR�ȟu8o�{)��0�^;{�`�F�N��U�!;���Ҁ��.W�@K1� c���༼�꺦ڤ0��'>��.�Oқ�3 ����vƲB�sҚ��o�v
N���.AZ+J-9sr?�`�R�݇��>���b�/\�.�[Im���B[��O}Ѻ�߼Eb(�Q��.��`A��jԿ��!�dUm:�D�6ԭdg��}^U~��f����U�\��S���f< =�U�|��ɞ��Z�BB�d=	γ��x,M��8� �]�u���N��l`F��ǛT1��"N�'����
�{_eXV�R\��5�kd�� |]��#�U�T�ۮ��GLH�=�Sշ]�����횉�c�Ϯ�!>Iy(e]�B��Y;ᙚ���0#����'h�&��+��D%�|���)�,�-��ExqL�wZ���(���_��p��NGA��7`(���o�_�J��Ϳ4�{t$�L�`� 'B�[�~�����3 � Y�8�s��bl��U���y�:Y�88�X�kg��5n	��\XG��8<4ɤw��ͻ�8��|�~D5��5�:c�<�Q����Ž:ޮ�rg����M�	�/���r����^|��Y���o�v��U�c�e�+K#��-��� W�O���8ڵL"o�X���;�_!�V-Edlh�����F�:��ػ;h�	���D�g$�*OL�Ħ�韩�kWĆ��9z�5�=�3�[8�,zx�}�>���w\��i��Z"�k��� �����e�Yݽ�lyς��O�e=*8��OTC�R킾{2��&sL�x@�D�'�=���Ck�llG#�#	3������}%XkƧuk�z�ŭ#��(��/�f�F�6.#����y���GX�(��ߵ�إâ��ŋK�]4S�K�|�� �=�D���m=��ԯ���B���|��'12��f�<?�2C	-:W���Yɽ`숅5g��8�B��,�dkTّw�)����1)���\~�n{�j�L�q�w(f�F�#��!m�����@�
T���ǀs�B�(����Q@�{X����&?��%B����:'#X?��G��+^PY2�ꭟ캞�Wk�A�m�&��}~�lF`[��T0l�8ԝ6����(
��n��ﲁ��n�����]ږ�iǐ%�4��~����أ�~y)��	pV�ml*�;\����1M��I�& )�8]̈́+�}�aȱ��lRY-xK����k����P:y.0h�@���^�ԡF�����#1�`�����!LL��W��d�YUj8��P���;��1|d>>���l����FBϴJ��*�$k_c-���|k���<-?���n��.r(�=��C�.��n1(�`"�l��î�$��H\��zf���2"�3��@��k/�joj���{C�7H�(�Q��yp�@�y
��C��	�x�D�[H_Y����;ϕ�m;�����ϙ�o�gQ�wV�^�����5�'���Ǔ�9��~���f��`+g�?OX�Ԅ��S�ts]����J�,��1���}��YS��&�MƊh��z/e"�%��dC��W;�XD��.R:�4TTIlj(��rJ�IX��T5��z��Q�,�m!0I��x�`��]��m��b�,��(,$�$5*]�`!���X�e-�^��p�����N;��R��r� '>�9����Cӧ��,i�t������cD|�ݼ���[	�Y�t`-O�فe�/7�l&Spr\4l`ڊ�HO��'b���ï�C�9� ٩�̔� IO;��`�!**���{hp�w��L���eQ���̀':�mD�e��ɠ�-�N�:���ٖJ�X��q�	͈o�4RO��4��9��x��х^D���s q��x@�?�;�������s�{ǐ��Q�%�]m�jQo�?�6;��u��>c���?x/�=�BN���!��*q�[d��b���˒��73P{�m��$��/<F5nn��O���
4�ć�`y��:eʺ�$���:~ģ8è�xn�Z[Q��)�$T����&q�^b�7gp�HIiܿƞ��I>�f23���◆(#�㮰�s6�f���5�)�,u�����b�����B��=���4�Ih!�aQ����"�Ob���$�2����ݺ����:^���K��WS�����ZK��b`j��N_�4�����8 ��$�/�H~.��z��%V� ��f
��°����HM�����Dأ[N�����1⥔o.��qB�w�vV�����V�3\�
N-�\�Bv�<���%h:���ۉ	�J���||�M�vKK���x���/O�>'����R��Gze�U�&�moYYc�xj���i��y�i�`6�N�,w���-C����{kc~�#�]Ϟ_�Z��գ����E�bo���l�g�N+t�kF�7�iy��VM�&���}�Ͻ�l�%Z�; ��P��y��R�z�D�ZMv
��`�3qP�w#�c�j�������A�Y_��Aw�q��}��Vnj��d޾},m٘#I���E�+�_)[VU��<���d�Df�G�`������i��Э�,��$ċ�M,"�^8�\==8�%�4�9CHr��3æ�I���`C�F�"AY2$l��L��ʢ+m)�nܫ�́m�g�Q�&9ݖGA�V�]��?��b[���k�Ɲ��Q���N�%l ǉ[�'l�ã�'3|���A�d����*ˠ��թY^�fS �2 ������J���a�vJ(�ke�zS��J�U�;s+�mL��=5���.4�Q ��F������zC�T��1�vW]M )|NHO�WT�Z��;�;xH��q�<q{\���6#%��y�ɣ�k��5�s�KQT���ל�d��PR�ů�oZ^��-��f��-����r��k�����}�٬ҝ����Ǭ+�ˢ�6PO�$��ߗV�~L�q�I�{�����q�}p\���~w�w�R��#`dw�x� ��Z�\q��]��~��T�������N�F�w�Y�8���1��*��`6�q+����ㄛ��'m0@ף�U�)�ϔe����nl���+'�ߜ!<.��%\<���_̙m>Ϫ��XY�7�^dm���S���J���i��I�}�8� �\7[�u�pש���ï4���\Y�<� ��ȥq��>K��;f8>Z����9cuf[/����1 ��Up���#��nh��֔w��e�Vm���
�P5F�>f�wq5Ր�T�vo�+Њd^�[�ݼ|�%��njd��8�0��Nq��'8!������ds�l��o�J&��|iK���i�-�=�O1&{Z���n����j���K�;Ïf��c��2���4̓�����Y��{���Ly��	���W7l�i����ەS�=)L�'��EE�,�y������CڂA���r�MPj�Y���e��3�`�W�䡳6{�^��w��5�m
/3�S	a�-��p�9�
zټx�l�=��}��)���al\��Y���(N����=}���̻,���eq4�`N� :�2�����]���k���b\�l���pg7���e_�G��vj';�S'ZTJ׌�������s�S�fh�C�ٲ&�0�}�D'�J��� 꿨����>��	��!`Qs�4����A���:�+ؐT����������Ț�:��V���`ؔYJ�t�"�����o\fn��f�P3��c��5ި`����'M�p���&�t^�[��**7%�^'=}ߙ��T��j*^.�s�|����Fٞs��-��5��{�;�=�9Տ����`<�r�Pn���:
6v_|��h�+��w����+��+��>�n�w��it�H!E�g`��t~[��+��}
m��a\L���	c5P.��`�����);��R�-����(i����i��CL?:|��{�.��I��?mŃH�җ��流��j�;�ݺ����ʁ��U����V� A�-^��� �!N�u�yG9��HO����6'��B��q���i��l��_��5к��)�ӏ�yN���w�;Z75�e׋wС�4��VׅM㭵q`Y����j�q�b q�U+4��u①���7[ -d��k��{��i��d�냩�03\6��_C�7o�����+A��G]��@�����rkH�	��o����_��y;%�{ x��|9 �<emv�˼2ǥ�t{E����o�����s�_��_=��������q���U`٨J 0��Il�g_Yj����_f�������+Z_��5�7����d���C���URR�3P�I{!mBlj
0�H�hk�	��=5/vk�	�:��j���u�(w�O*�S�Td�B�yh\7<�m��/�(ٜxyS���9���a��z' ���(����k��M�L�4l�sv̯~g^����b��?G`�itM}��J���ʸ�c�'�nz�.5�	�H������?ػ���	ʲ�%`
]o]�c� �C��kZ-f��0�f�L�aD����Ф(��0�2�YLA"G�h7  �R,��:�EΧ̢q�f�b�_�$E��OQ�C?�p���`��	���51�Ϫ��:�=�+j������O��o��]S�����?{G�����b�����͟!OT��I}<Bħ�c�B�K�9 ��j�m�0����f���� ��W �Ӹ#�i�`���'�p~~N�����ڱ�y�F��%�1߹{sº��ɦP�9�7G��	|��P4Bdn�*��<�@$5J)�e~z���^�����s����*�s�	ܯ�:�Ex���Yܮ��?�P(x('�㲦���̀�4{���\+�[��UT� d�t.���\d0ͭR|�*$��!��~��ݾM�����m�����wm�x���D�$��Y��4cnS1�U�kc�e��T3�(���3zR;U�%�H�ߝ���?h�ʔ�cd�$�,ȟ�(��²"J��Ӡ㱫�>�x��$�rs���ӓ�-���k�A�#�Ę�M;D%�$�V )A7�
ca�O�w�XC���t��(���,.��>�n�g�R����.���e,���MɽԆ, �#y��D���O>;'8o�[L�_�X�}���>&���n��{�鍩������s���ſ�,��?�����^��_��yHL�������=���S��Y�jg��Z;���hh{D!��<�z�L��}��ؚt������ew{n��XøO -�X��\&¿w��;@C}=J�pDR�J�2BD�2�DS��E���o�4<��̑yk >��Λ�Aj���-Bh��Fֆ��#<��rm�����E V^h�z���[���P�F������������>�<�$~RR�M��3E�= hF���d��:�Չ�0U�٢}f�$x�@OSbFc�7�l~Om2����e��,�È,�s�{����JP���Ca�8��X���I���LXmA�Q�� ����fR�NFi]��0h�N�_�$�"	�8q/�x:�>�� ?�(5~����T1����� 4�̬�,+Jm�H`&%��S�p�{��Ҏ�/X��#�9,�=��۲@��Hh�䖲io:�MۘHy� D�RC��y�p�l�	�ӈnH�)� �D�)o"vH��� fX�x�;���<���u��:�11m�i���G�.���ȝ3�F`��g�'�3��4��o%H�"���QfJ�������$����W��+��?��ۖ��җ�4�|�j�N������O`m�0k+rL�)������� Bc�1���m�t;��s]����u?m�#4\�C�s�j�64v##�WyW̃y�s���7�u���*�pӇG� ��BvFbg	H��}�?Y���jwZ���>��ϵD_%��z��ô��Z��ۼ>�@�(�IIU������4�����Q-���lǘ�J0�|f��J��0�4��9������dΙ�*<���\�(��zR#H��@)�{b1G&�����¿�Q��k�����f��M���F�9�X"9��0@����5��3z������&O��l�5`�Ϝcm����?���E��M_�p)�8̤b��Fض�:�\�ID>;��"%!�
����>��0��P40 �
=hX�ᷔY�q>05�:(�2��4v��
	�2����A�4K�N�*���δb"->R��S+�]�C;+c�h����Z����]�<O�k\�9t����~~�/Nٚf�JAa.�{U�x@��`o(�����!m�)fQk~�O����E��7�oֶ@w��Y�o��$|�?F�i0"�d���8�O<�� �&d>�`�Z��4���/�����Lq^�Ģ�^����l����V�����>i 'E�Ӛ�	WZ�-�����y|�mu> ���`>�����ہ`���և�����!��1�Nab,\\�q��l�b���|J[���%/ƔsH���\5��`��w�1_D��ַ�@Ƚ��>��O_�^X 0��u|&��{T̜�#)yw}}������'td>�ݞ��B���k`n���d1YL�+���c-��y2������%	�	�I����L2�ϖGk���b(a�y�+X�WGN���ҚMG��D^�_h'i&���Z]�F��d��Ջ؄����p^u[��K�G����elk�(}���������$�!�8s�[b����أ�_����0}+�efv&触�`.s���G#I�:�NP (ϟ�hG�fҁ�Ћ������b���[��Ƭ�A�J�ו�֚6�'�e{��\�����/���s忭�GNb��g}M�:���S0�\1/���<ȧ�d���� DL�kk�=��:�-ihA�"8H��B03ƕ�p]s@�-���������^T�z���=��;sR��5�jgл�;��O"ax<ڠs���g���4��v�q��?��BRqm0��l���˼;���g��f˚w�Gmѩ���Ƿ�Xs��a��^�\�w֥����ښ���P�S�Ľ9@�j�ޑ���Ɋ��BU~�T���w��R��b`�ˣ, MH�&sV���q �	��Κ�ͧf6��t�ޣ=ڡ:���6����L�f��8���f�^4`KI�ﰛ��6�Fj ��fI˚����-����̜�Y/x3KƲVkq&^�iS*M:�S����v�E�`�^tf�����fH�U�4�u7� u��bK#L�T�X�Ԛ��UdTe�}L�2f$٧I4#ot2���+�0�O2wL��6礓:����hp�_RŹ����_+/q�6#������L]��P���窞Ӛ�j�g�yY�!1����el
k_�|�$��t��fO�@Cd�S�ΦG��wc0�7�� ��ϘNc��=.�[�1�~-��1�1��T�a}�a:��,&[� Z@�}�
�4S��^�FкQ}�ͷ��;��t2��jE�fu���/̃]x=c��F�4�AX8�9�������R\�Юh���|G�# �e�h�n�Q��U*�i�?���2YCۍ�����0���rH�χ4`_�ܥ��U?�7�@���#��t�&�L��cP�x��@�zњY���B�VQ�x��R����|��<�Z}qԪ%�&@�5��Xm��s���~�Z�0p��g2�� ��X[+�����`"D�1Y�;�Z:7C�(�E��>VL��]:�>1i�Ұɭ4�%�� ��u�P�ז���mN;�)s�"^UX;|`n�$�����$�Xo*Ϗ4�h�Y�V�7c0'rY�ő�P^i�NA�4h��T�W��hoB��0��	T�9�bØf�N�L�ꪵ��bƬ�R��t�w̕5��S��F��eY,����'s�J��裏�>�ϴ�y��QI� �S���e1�d� ��[��*�S(%m�� #�0�.���f)~��!�s��C0G��&���|�@��>�H��9큿p��7 I?��{G�mO[�f;.���~4��_�W���׷-����!Ǭ�1�5��̿�_m�Z��,�s�������$�w�3�}���w`����L
8Ƀ;��_�@�>��Ve�9~��_=�nϊ��W���4��}����	1�!3/fH���<j`3s��m,ǹ���ӌ�d�`):'S)r�~�}n�̑�Y��`�vk���/��TU�qv&��<�6�4�Z`SK���o�r���&rk��b�A
�s������3��%sƚ���G$��I��Sd\���M�vPt+�YőϾ~�P =�� *u@Z�9�W(���G���S��&I���N����G��.�P�KE:vu���B��(��o�s�0�RD[�(���k���\�h�%RZIF�P��Z�y�J�ۂ�����X�Z�#R�g���N�_����\	���z��ԓO�|� �#~�~�Ĥ ��Z�=�\�e��1C�L�0"'�J�F*~ ��-�۲`��w�62����0?@���X)t���ǕFjNM�Mhk�VkF?�0����j� ��q�ﮘ��h���k�<p�|Ɠ���O�Z'�إ-L�m[p��ܩ9Б銶-8��݂�ϫ�xŚ��N���kQ< |M��0e9��wL_>(��/H%~T��Xc51� ��,|��,��hG�yS3�5$k�f�f�0 /�Zê��M����QL���M1�K��q�5U�g�U�5�Zk���s-�q�]?s����`0�	���y�C��B���js����~ZKh��7�O���i����] ���	�_FJ�{�h�بm*nC��-L���)��P�,)Y�!�MIXd��x�7;���y�Q` PTỎ�ů�G`��4f�Hd'JX�Xh'��PT�Qb=5�8>L��jt�:�.kz2���� "91�����)u�3�5,j���.
�cB$����Gh:�ޏ�c�k��.Db3`F�#��E�� @44���'�OL�
pk��`z6C;(�1@k�ӕCxNڳ&���qx�_͵�[P�h�mtН@v�}x7�3O�� �����-`h�ù}>������o�9�FYr�b�R9!-*Ӫ�?�v���\�AG�-􉠄�ڠm�Ks-g���Yb�3׺_�S�瞼,X�к������ՂG��C�Z��	I#vBp���Z��I"<��� �8m������3��R��q[r��+��l	��<P�H�Tl���5����ٙ��#Y��iU�8^M�'�@�g4p��z�|��r�9����� k 5�oW��M�i"��Y T���^�C��Z���A�D\�G�����2ɩ"qO�MO`B�תL��a��Ъ��y.��N�g�$W��;r��'��e��&4�b�$�0 �X�� )�.�8�b������*�F��*���^�ۦ�bR��Nu��{�fg	pO��#x� T{<�h~9����63�'��<�LEh��>�� /� �O�%!�/����f������q�P8Ƴq�7�����L�5�T��J{ �<�7׳��/6����bߒkP�iFiA������v���֮�Ͽ���z4����1?��?+km�DV�#7�{�Ú8s�zg�6��T4Q���)���t �����E ���;��Ќ������<�����.J�Z�㟑�ޤO��	�&��S2}�")�~}F��M��b8�_��y�D�v�!��M'����uȯ%j���RAs�p���O��ڞl �AO���Of��Ǖ>	�HƖ�*e�FN��r�U3�&q�Yj��3��d�
���zjͱ���!6�i�m�U��E��-Uh˄Z�2���ZXw��ÇZ}ù[�*Eye�#rsY{�-�L�-Q��A��EJ���vH㉛������MG�Gʂ5��a�~�^�o{-p����&��c��kӼ��H!�{-B��0�0Ճ$��1�w�E�4�EN'�1݃ńZLO�Ib��T�����C��s"9�����# Pu9[J|����Y��"�YgF��>
�6m�0'����O�Ƌ�2��p�6A{.���@_a�h���O�ڋi��ڽj��-g�8 d�f��@�����5p��@O��g͜yp^ۤF��� 9��Z���7>�� �7�+�V�y_kp��pe�x�Χ?� ��y�RS�wEm̈l�W�;���/�b@kR�Я�ʯܪ�[��g%ܩNWǧ��1����	SGt�0|�h�����T3k^M���^<֒j����1��d-Qk��1��� k0��
"JM*7d�X�c	����95æ3�e3%��9&@kH��T��vn��[k�Jktf��H�	�'R�e���l��Z�;"-�ac���أ�{��5qp2�~S�J�,���x��a]���+sYaZx*d=)�}�㭧�z:�
�?�½h)�*�F���'��W�������F ��#��VL�h������Zk��Tp,ݟ��[����jhl0�����8�,�:��㞻-�7���J��d�n�M��'�Fa��.�*Y=��-�;��N#�t������A36]:����s����azL ���M�E�P1����Χ�֎�d}X;���W��A���M�d,�~ߒ��|q�!�C�����ѡ���b�d�8���NnP�W^��T��[Ξ=�^����w �C�)t�q��!�1�k�E�Lk� �uPT�m�$͋�a_��Yy��YR�D���H�	{�@����Y�/'������ݩ�Q=�Au(6��jV�Ի���`ddj^��l�֔� m`���M,��P�:kFo�5^XUW;�~�[�f�[�p>�ɓ��%ȧ��H�LX�����3�y����%ǧ	ܖ�h��/��XJ��fa������Z��`�1�Aٿy~B�Y�D����h1�62T蚝��V(xMz��>�R]O<�n�>�c�[�/��F�U�V�&��Z�Q$!�	Q�E�����*U[hb�
���F@�H���"`Zi9�¿h�C�QdaE>�-�yi��E�q1~�fto1QF4k�r��dlī���QWU�/ޔ��YT�O bl���g��u�+�=c�=k	֦[ϕ���0n����J[	�H�$�S�xV~�$<���'��gx�����HD�я~B��N���oh��7<��¼,�䘤 �5�O��o��d=��Z�/	�fi����w"%�מ����g��`n �x��<�^��_�)�I�t��2Fی/�e�߬�e�L�����	o���l���w�H:j���$
� �1���c��Z��|h���v�ͤ�����������L��K��kO@�p��<�tyLe�>&����ZL���T~�q)�Z�M���c�oK������ki��Wk?>÷9�Ւ��<K��6Y-}bB��#]���bNŚ�@���Z�+\75���<�b�Q�� �S�!I<1��9ך�?����2���m�H�}�g���{N<�|֦�Z�����!�-j1I�r5	�,�! (�3vYG�<y�������XDj�P�����#�[p��ѭj��� �'���η�g������壘]�F�U�W 7*�Iijk~��j��֒�})%ʑ�9����X8hZ��j��A4�o�39'4cv�^��@����>D��/ZX�&�4�.#6v�8E����p���.��}��=Ο��
f�k-��{�=����!M fP���s��(�Ԡ��d�<�>m��O��Bcj-��0+�A�GD�'G� 3O��X�;ŧ��(��z���JhJ06��aL�~s̚���cv�K�3���c��|�A/�#���Yc�zh�}��N����
U�F���@_��a]����:������sԱ�]vk���,XAmM��f��ܦ�]��8 N+���">?����ݧ�� M�!��	�K�M0��L���w۩}�R3dem�k�r�52�b�ڢ�z�1��U�9KG�
m���˗�L��ȳ���g)*KpB:����fS뺀`EZ	�n�gˍ�C��γ�'�oj�aFjMB�Y�ɣ2kv:<��RKo�|��MR$�J��Ma��M!D>jW���>��O��x≢)L�Ok���Hu�]��S�f��F�}igum]�Q�f7s�b��i�b.]i���so��H���[}���n�Fx띷� ��1���Qņ���bbB�π�	6+2�Fu�y%��������D
�^Y��+�m+n�5X|�C�aL�b�c��oda�^U#� !� �o�G�� �
}�S�Z����$dq�#}B"G�=~�&��CJ�P������[��_S�A���	h9������$}9W�aNYG6oYj�@�Q��<��C+�fG��k��n�}V��>>�3@HR:�0_q�#A��u=4(��y`�h�PeΙ���3�vs�lg��s��fq��]kl��w��%������?i;_�h��y���&�7Z�3�ح�>��_lD��pW@�k��kǩ�"��g��O��wh��j0��j�,�@<@f�Y�6��y2�^$5x�}M�ki�f#3���d��ڠ�OV��s-ݲ�]��IE�ACp�( @�T[��/�w��ob�k��I����p/��yF?������n��> k���P���M[�<�kp�<�9����S�߭I�����w����z���_�S<��i~WT��Gc�Q&����~�L+�C�9�{�i�3�J½*�qn�uV�/\�i]RB��3礑)[&�-�U��!	1�W�C'ɜ(Еbj�d�Z�>z�q�� ����l�7��ZD�J��R[sY�F��wo	h>k�����gk�r3P�HEka)^�����3���o=�������׿�5i���a��*�`�\�:g�m�tޟ5>��^��9���wo��MmC�.�����[��i9��J��n�ɂ&A$Й+氎l��Ź�4q[�Юl�Z�0�X� UQ�#m"�sh�<��ti�5� x�K�'s76�J��kb��s���p� Gx�y�w4+t�)��_�]�2ӂǏ����6�St��>-ȷ�*s] ��׿>�b�lw���_�E��.�8��v�TnNg�T3N;=�a�8�����f��:�k�M�Ǌ�(&�Ҽh9ώ^k�&D о�$my߫�zJ�0�Svt��<گ�ۦ�4q��w�o(��'���<�鍚��ڝ�����쓁��ܧ��,}�m��W3����͒h�qs���:L&rSgu(,��f�3� ��?��H���`,�,��M�W����	�1��F`���EP��-��D�&�� >9J�]�i��*��Rk��ri'���8P���䤮g?��(�.M��K����]�(���+�k����4���`%�B��c��0M�@ �C�T��p_����0�ڗ\'*'M�O�F��L��MG���O>!M���1
b��7���8D����[��+Ƈ��o�% �:���� �����Z �F<���׊�?�9 4 *+���Ϝ�d�mٌ�(_�����NI�^#�K<�y6P��M9Ў~Thf ,so��4}��b��&\��l|���,B#.�M�/����E��������lU�m�ĸN}��{CϹm2��@��/yD ��
`�ϊ4{ZL�&M֨}ށ�N�q>-0i�}[M�\3`O�M��0��͢f
^l<x}�M{�e�ی���>�;�Wk�L*0��1ih��8@@ X$`G�E_{�4���h;|���܋/�V��%�wY���J�[k|ek3 ��,$XC�%�n~��vmM�&d��?��8�\�F�~n���c_�O~�*���4�{��!̒6�r/�1�m���[01�H("Ws�Ο9��7�x���?i��*��uJ��$-3?e�AMTh�H��?����T�ԎM�'|&A<M��_���|"�ah��4��M �4�e�����32�0�"Q���B	����)(e������#gT3 �-i[���q������ᨊ��q:{�� z&̥����@6�۬n�L�l��if�ߴ�����;�a�5H� �M��&���y?��3w{�ڲb�3��أ�a���)PC���3`A|��iZ0��#^�'����dy�p�nW���@���p�#GS�c�������Pd��&������Y3��	�A#|H�g:�<����wk��=��2�a*�������7�������Y�'���L��d�d<��F��X-7��f@�	��y�ݶ�_��� ����-�s���3,kmɚ��GK�YI&7���p=��G��];E�s�v���/>Ų[5{x%s���b���`гӠm-���O����M4S��ϷFl@���s�dLO��@nmý|סy�+���?�z���@���R) ��6o��Ǿx�!�����}���T�缪��.�{��?j���Ni���gH=������@��#�,�"�"%��`�v���f��%�\�)�S� �H!������~'�Hb?�2���tM elmD�����s��`��8F�A�X
N�<��N�t18�f'��o"f���ñ������'xAQ�n�	� aj�`2�e�dsi �m�4��J�\U����ޏ{o�����X͢W�.��#~c�m��w�ڵeM�ߘh���Z�o�m.^�@H�<��7�ޮ��5к��������G����Jt��[�L� ����m����3ǠIp���cN֧��su�O=���2���uN��BT;:usu�@��;��_�*����!LR(6��d�fF3ck >�`�>g-%xj��6��~����~�~�Φ�d��@��C��@B�!.�^S���[�^��d��'�P�T��v4�_��ECB�3�W�9y֘�I�m2|���j�r����TSB�5Aku���A?�%���73@K�䯱U�O~<�(U���Sf���y�1(��!;̏(�@���;k�i_�7^~5"�(���b^�8-*�h����}*�� ���G�
�؂�d�e6��,�x�u���#����`��&}a�c'�2���U^x�H����P�F��E��QLAZ�b��0������a����I�i�9Ӏd�P�L��U�{Y�KZ]�E��4�D;�[�^�]���4B����yh��b\X�c00[�j���n���H��=�m}b�a�h~hé}�VaL��Flq��ѵa��[��=k�<;mC+ܟsh��?��Ѷ�{�����(h�@@��N�ܟsy��p���W�9n`D��Z�w�	됾x�XP����1���V+/�?c�n�]<kC�<����#� ���.>��a���f�Q:t�f1:��Ԇvʻ�Ѓa���+_Tq�-y�n޽%��.k ��� �53s�Wm[���޵���I+�(��?�c݃�W�c=�m�h2~0�"m�lNKzH�# �H�D��H�>`��'�����g� ���	�@=.5p�Zo�?���L���&}7�c�[��1O���		 2���7:�5"m���!(�Dpuy]�	Ҹ��p&��������So�R-f�KH�����7!`��Z��Bqu&�&T#N�k=�
r@e���z���4m3�j�V��X��i����X�.�}D�f�o�q�vF)q��Ȉ m�4�py�%�8~�Z{� �|�}
���0S}�p��jL��J��Y�^�l==�+�����`< @�&�'&P��6�6A�iY��8�7 ������p�z`<�J�D��ԵS9��v�g,�'m��N�ʜZP��@O.g+�j��s<�@[���ϡ3����FjK佸���F@��׏;�'
ً���`�z�^�7��7��Oh�֑�׋�f�lέM�5�r~b�p�=Jn�������e=(�v��`ѹ��M3M����ɐa
�a�6�Z�� ۑ�=4�bj�*�ސ��U�3wgW��m��ύ{4Ͱ��֮��|�P�UG2̑0])�}R�0i�$�F�~%�&�hWfP�\E����EC��� � ��Ui ݯ>�\o������-�L)�<
Pح���mJ�5�6�Z���`��1��^Jy���t1)�����@��N�y��S�x�5��G�TC!���P|�a�%���K�]Ѯ����$A���E�|�b�ʙ�Z��@/�^n-*?O�&MO�k�'f�9�R��@sDe�x�)X�Wo@�c�^��d�CCJiX_�F��v0%��q�N j6i�p�4%&
ľ��2쌁:�~�y�������K�,]�3-Ѭ�EP�3�?6�F�ȜB̬�{{𿬄F�]!�;���;�1����aY��L9��CY� =����m��P`¡���G��dsݙ6k���������1F��������
`��e_ ��� �F�4@�qD���{F�a�\^�#����]{�)��@�U�(c��NL�}�bM@㗔��(��u�%R�P���[X���ߺ,_�E����2���)�Ck�5�{bV��.B����u�|ڌ��������B����	�%��� �ɵ�8`��(��|�^�y��`�����	G��
yDO�0j���Z�?
��"&] A2��K���|Y�j}0�3��B�~�
:dWC��J�ym�g�����_�ĵ�[t��JYH{wbj�a��r"zc�s�䞚�����6��-ש��^Z����)
ɋ�dC��ԋh�SK�����|��W��:B��mZx�Xck�M��󘵓zE�Q$@���P�_c�;dn:)���d̡��Z��g�T���X�S�,��/qFg��R�3*�tE��KZ�k؝X���M�bg$m������;0��m�:@�wLܚD]��_?��9�S�2�����c&if�(p0������i��󢾡���Y�Cv��. ��"��{�;B��&��x�)T���bvY��V >$x�R�#��\o���JF�����n0��\��tӴ(t���h�^c���v�-?�|�넵R��`�<0o �8ʓ���*�
���˵@������y�[�!��
H�R%�O;��@�������{g
����k�i�V�(��z��T�5��b�z�R�א���]�ɼܖC����g`yNL�N��i��;��έ�ޕ�q�͌EH-��5���E߻BM0�|R�`�#���dh�f)�Dk5���\L�Pp�SJpM���_O)���g����qr��z��4Uv��lu��l��b� B�c��Ss�⟚ OD�牷�iM�{����L"���'�-�S=��ǰu�A,�	fPk���1��������V���dlbs�G�^2���5Ss�K��F�쉉xz�`�
��+�D��%y=�@�m�e���1��ܣpPfM̢�ʚ����o��h��7�x�����4�E!�rK�]әk
0���JA�W_z�uB%ܦ��JuY���!�-Ѩ�]x���ƹ}G��i�߭�p�綆���]��q�/�E��L�~^�_R.���ADUh�X�4AI8$�_}C���(��}��U�e���p�,�����	J �	������NjAl'z��3�\C�M"|�k+�}D���m`���	�6B��ô�z����X��]IŁgV,��9c�`�*�Z`���i-��
��s�y̷�{*)��l��=��Bp[l�9���6�gDb�N0�APi�ߋ�vL����<���p]�j�.(��B�&�W�[�������X� �m�0O�6�f�(���?�������ȶ�m����!3L&�oTaaA2��k� ��Qk���$��ms`�!���0�Zk���c�۬��^�^�^�	���+���1M��;ZN�{�@KA���d0�8�)�\/�&�2�bHJ��v���R�h�����`A�vH;"��+�r2��7�8.�6{1�h�YP ��.�D��·�]�)@��K��� ��U�����̌
p�.�(���5��F�C�[@Z���N��:w�l�*� ġ�!8�ҋ	(j�&}:b�cԴ|xQs.�̭�\f9@L���QƿO{���u�LJ=�n�ٔD,���W^��q���otq&�j��c�`�2s�o]x�?bг&����f P7�jҍ��^���A�Â��P�����Z�	�N �����v�{o[e������hP~Ԝ8n�y�����]/~�nc���,��:}����hk�Ԯ��(`�Xl;&RA[��#*�m-�/�}��;�8^37��c�/�T��5h���.��1h�ֺ�J6W�B��fʹo!s�*����竒ղ@�|��n�D߶�F5Hk��Y}.���,���5�΍i�I���b7���m���:@�����K�ͦ�N�Yր��<f��
�$�+��4]ya�oynj�<3_��{q]�B^��`mþKl5�7z��ݔ�k�n�i-ԾC��C�뱵��8Ct�h��Kl����.�v����5��d~Ӻ�~����-)҄fl��.�2�6��X�3��{�&��̏������eU�� 3����#5�e�#�-���j?���sb�����S��X|�<\��I�H��z�*���05<3p˦s�����:�o�N��]���U4���|Џ����y1�0(��ڵ�� �f�N���zͻy��^wּ��};��\ۂÜabc����l���j�����rs`:Ԧ>kl� ��g0�BS���3:8�B��u�PΧOЫ���'|Qk������D}��8z�4���w�U`�!�Ռg�W[��6�xfzȒ I�}�i�ca_(�/�}6@�O�\8��;m ��/�vц�m�����N��X�Q����[,�s���a�c�$�ڄN���DWL
`hZh\Y����D��F��%X��Ru��*[ �}~z�ru������",;D%*�Ć��˻F����U2��gTU�$�Oej$�z������\�n���1 3�����J�$Ml���2����	�*$6�@�an+�Sk�֢&����l���[S��e�����ftQ�"I���O&�� ӑ)�J���.�L*�_��@r�z4�D��hb��9j�G��}_hϔ�"��N���5C�䖊nx�>���� $c�C��65P_P�����8�B^~%��KL湩oOk�P��P��@�q����C�;�\��tz/���>��:[(�[��^�3��:�>a�w��p����0h�%0�$���6�X{G�������Զ�Ys������2�z4 :�&�&����{�9�۸vzAk��q!�F0��a栎���4��3�X4op�Z�׹y+�o�.0����X��0nXU�|�Z���i��ڢ�|��dΘGƺ�<�H�^V?4���UV�@������Q�������j��%�o�i�]h:M���D�m���f�p�Y�oq��P��7�x�\��߬=�=K�N��5F��WǇ���v��)�~�!kD��&&���"�<�\A��lS&���ˎ������I��m��s�DAB	�v��, ρ?јM,2��jk�%���I�8��ԞR�έ��I�WR���J��̵.�6��sF@xE9� a��D���1GF�z2�ý�rP̊�5�!�$B������a�:R B{�(9��s��V9�<�^_��ZL��sXq�J܋I~�:���[xU�*R��p1ݠE Ѯi��U7tC$}XC@Q?���c8a �������G����_S[@�n���vB��<� �cr�c�1W��ܖM;�h.a� $�<c�V�P���NL,�?�-k��T��W���Y����\���w�k�6�Q_P�{>XoW$�b�'�4� �����_#7W7�{F��~��pd���[`���O|���3�so�v9n?��=��r��rZIIY׼�뽨y�}��n]���4HuS=�z�.�Yr33��[�gpY�p�@o"�J;5!���LM��̷|��Uks�I�`�l�kk�L�A���$�9���3.'O��ӔCvcҐ��X\ΈI)HL���&��� �f�hJБ�p=>{eP�X����h&b���hP�8r\�%F�ce�7�����y#wi��ok��Ly?�!��;�T��-�fg�	��4�K�BZ��&��_�Cp?��J
Ό۫Zx��C#N�oT��  �H%��|.���~��6Z�0@?� @��	���� �X��):@�`n�i���'�Ѓ1𷓫��3#������L�ulb�u���c�ph����S�+]�:�^���x��v}gna�*�Gs�B�<��&�#�A�w�C�D �1����3��)�[�?^̕�T�4M?kA�F�5����L��V;��u
~�u���v�!X/��g���n�/g#@��ZF�Sͩ��`R�!Z�o ��/�׼����Z4:(̀��\�|�M���Rq u�~�Ǭ��y���g߽F�Ĩѫz��*�����Q4�/k��1e2DG#�,�#99U�����2�L(̜��M��9�������� S� ��a�qn1�Z-7xl�����}�|���9�%LL&ذY\H,\cFI�\�]�#�4����y���v�a{����uk/ڬ����;�KM��(Q���VuVkISx�<s�0�JQX�O�ꕫ�K�W�73+sJ��@���P�6�H3v��֧v��ߒ��t���e����"h��N�%�x'�a�N�S���� D!a��(c�9�<_������v��E�ԇ��~�3�s*�����|���cŴ���T�#���Hn*�㰂n>�]�|�#:.���@S�!L؁7��~����'*+k��砍HO0�N�� �4>�=�5&g��\��B����_.�(a�6�q>o�ڭ��y1�d� ������-,XayP��2��¡C�$"m2f��긾c�܈5���$9]?8c�}���)�B�#T]�o�,:5/r�^����3B
y�<� |���q���.i��:gyhhdo@�b=����h�y�`�d�f�f�\����3���4���j2��[�w�?-�xpQ���vS����R�µaj�^�C�Ձ;S�3!L`�g)1���G:�ܣGg�@D�#� ��������m��'�1e{����<g;�K}��T�ԛ�g5R���#�;ۨ �H�P�4�4w^�͌KyT;�t�g�B���e��klf/^h-iq,K["4t]���LD�
��}1!�1ʠ��)��H�m%�G� (f0����q�Ӥ
{�-k���ni��L͟>��ᜐ>5�=��q�����ONjM<��S5Z�\�%壩�R�A1�
s?��.�t���	SL'�[�m%�v������60��q��z�ka�QCK�:�v���l�������P�<�*����ܗs`̜�]�,5籛R�v�� �6�\T�S��2��|�E���oP ��I��`O��?�7�aQ��\��x�/���+��.�>�����x.���ݫ
��;[�����Y[�wZSw�d����a�FS̯��Ui�;2�k��`Y���& 3�`m�#l����c-�q^=�	0�h����Z㱚�Rk��c;s�͓L�����M���v�$R&I"c�l@��a�R�d,)r=g������������n��1�=�L��e��:��L�1U!��7��2h�0fn0��8m��l�FH ���e�7����ȶH��K�uh`�j)�ߢJ&����_�,��1o!�2���U� ��蕉���Qy~�n 蹨�I�]"�46&� Ղ�1/��ǶD�0������[b�x*�ໞsyꩧ���c�wc���}���9���5l�M���D�J[��ynkx6{�����[�'k&�ラ�t�x����`��sCLw0d��h��t�/�r��Ia�. ي̩ۍ���i6�םӣ|x�5դy�,�ge�q�w!��LYk�K�оT�鹳b��በ���ODa��Q�vʌ^����!��?)�Z�/�3�p s��e On��E	��,�9"쪽���s��ҏk�P���=��#��S��hJ/[�G���� ���d�f�[�()J�6��)�y�jF�<V߷~���Ga���T��v�c��ؖ<M�L��:���̀��@!"�F��NB���up�1����5��F�c���}�D�>7���va�!�:z�~�Lm]s0�O��"�PfE���E%7���Mհ�ĺL�Ҵ0
�̏v�O͠��=�=s��l�km����"N��i����k�B3�盭��b�ek����␴��IbN����ђ����-�D?��az�y�*��H4��1�nk� T�Fjzu�
�Cd]��y֔+��"� ,�F�va���~[��sf�(�9����VH_ �C�û��n�W�&j^�s�*{I�mh�k�E1xf�0+�t~���N�>B��YX�0��LI�AK�Z�T��}0��	7��L�#m1?�
�7��Th*�nZ�r�u�l�+�X�.`�u. A\y��g\W�~Y�\7P�+�Z|D�F.�5*K�&�՚T�����Py����j�e=�݀3�': oeଙ}�^5�������x���g�@��os�&�`���02ẃL:*=�A�@h���@�dBb����s�s4A7K�	��P`��V\���q���D���TI_!pW������:��8��% I��̅Q	��h�����J$�3��'=�l�;�0�F}P�%�b���s�� ��^(��,u��5x� ��ҹϫ�,�casS?B��tM��/��hu���P�t`�>�o+�C�����qk��澦�zyn���}|�ϩ�4i��A6��oo-�q�X{�@d��\`�����\;G���hm���:�h��1������ (Z$ ��R�@@�f�kڽ�����n�Y璺ҕ���a��/j�}�zk�_�g��堢��=�s=O���Do�E>�1[Π��������'�0���2��5��e�����z�y���9�]�P7]Qjh�9/��M�l���A�'��0���f�n��Pj3���q���<G.�[���]�ۚ�	/�`�f�k�E�<��L���d@,6&I)�|#�P���i8l�q>�S;N^,^�<�%'k�Y��np�=�MfY;�q���x�깡��;�����o�"�;�<@��B׺�8	���ER�W `�Z?��ot]R��a<
}GX
I�x9'BTa��QJ�X4[A��eD'�nQ�J�-2�JMȤ���NI�XU��a����,.m�
a0P�����N�a�=휭�� m�_=&5����MS�'t��h��i�c��^��k��Q7�R�i�&��mׇ�0y�A�U�L��S��rR��{x-r-��z��ʺ#&ʺ�e�9�����A'jc!�p�<����� ���.�.���	.7B�1�0?Q4_�N\���y�ѭ����+���:dLi6�%�x:<�|��0�CӬ}� ���=�+-� �T!���Df�f
��"�[v���&]���]9׵H�gU�j�½�L5���[���K�e i���5'\{��Y�LܵI�@����"�����f�ݤI�_�Q�mKkp���o&�&�(��1x��0H����8�b�'�N���>��I�����^;�5�j&�d`͹K�'h��d�4�hY��w�� t������y�sh!e����x
,Pz�P�"�/A�����x4C����A�O$�e�e"K/[$0��AI�ЍMaT�g�wF�j;�b�N�-e�2���X�+*զ�����,�x�k�#��闝 ��"VY���-��4-"|��%���^�ל'ϟ鐾x\�
D7$k �k{5�������6C�!�q�~f3`�h�y��T�C��8�`ʸ�_Mz^a����;�D��z����+л��`��gt��;��^[�_�Ik��/K*��[Z/l��-੍��2N<kvNnƀz���G�y�ѝ��@��A0\����;����#�3/�Qc�8��&[�X�6?ҹ� ^}[@ȍ��@�j`��M*|'��ڭ泎/���*W��7��f���-�k���F����lJ`2] ��j��A@`p5R(�#$��	h ��ؼ� ���&/4�y�X�w����iz�w;�fF����S�lě�:�5�t\�V�p�xH� ���0�xk���Ht��SL��*��E3�FM�P�]��v�*c�@Ѯ�x�6���¤���iB2M?-�-�.`̢
�8�)�@
�t3�w�5:2������,i+꧓#բD�B���OȽJ)��2f�2��B#��6Mh�	��5�5q�פi��nmuy'���h	�����x&�`�l�d��)0F�%�Y3�?�]�%���h�M[���a�����hEW5a~훢��]!�O�O�}'c�v�����>�v	ܢ��צ�� �5Aŧ\��e���!]!i����q����/�����L<��ڸS(��桌��G_k}����F[6��λ��n�mƴk��\�p�X#���$n��~�	��'�-�-�s|�L�>w#7��Є�g���B��M�����<�����D���%2� 	���o4`�h�N�G:�Yl�&l�@�U#l>Sm�-��}� jF�'D9#fe��7{�(��sڂǈ�R�"�#H\G�Ԣ\!� C��y�6�fGZ=��� �P�cI�!�=K�Q�礼وv�`7����Y��=3d���"xF.,.���{��3��X<L�G4�w���}�|�q@��;��P\��Ƌ�C�Y�*q�L��/Sl�H�|���a���e���u̵��y�|wy/Ɔ�������j�=�7k��03�q�����r��8���`� #t�z�z"{1�"�گ�zv?��v�q;�X�p�����} ߫1�v�����F������m),f�d^.b����ڜ�ƴ5۟���>Ҿ�ZS�\v���?�������\�}�8 �Z�5?�cO��0�q.��k�XVDgW��v�vc�.�Af�J�>ǌ�6c��I�5B����I,�e��&��������kDG�����J�c�<U?��ƀ� ̰̌X����l�o��gs��`��ۮж��Iw@�M2����Ry&|wƦiF�6W��KI>'����:��~�ߗ����vnڎ�(�b���V����>�mnP�Lc����B&-8��.��	�&h�s&�����
f!����p3����8����G���P�&��K	^�ih �f0@�o���k�]�	�q��2����������7�������^{50� �QWf�t_xA �胖ؚkU�DD�0�B36K���n;V��?s��:På���Fp-8��O��d�`x0^'��Q[�bmq��S��~'kd0M�� N�����6���=R� ���=�2h�A'���ق�ץ�ٱ����<���F�Y�B�:�1��\?ټ(���(�W����[������/ i_-c�}�2�ј�|��Ƚݘ]�y�6��	_�v� .�;H�;V0�W��M�	�s�<����EKz�G����9���Fi��vx�&� � �K_��8�:�M	j��[�~b�:&�R�-������o���!�R�h�/�~*M"�T������a�@�e�"�ڬ���8O�������ٚJ��|3`�$�ǳdʂ5?�i�5׋��\vj����t|V9V�����E],��MS���������L��NJc[�<γg� Q�J�H����K��0�<@� ����/�����"�T�b��Ar��
�FA��[.�a홸��T|D�a�y��S�!�J3��[(%�r�f6�%�N�v�uw���6(U�}H�T�Ͻ(7�g�֩7BK�����~(?�|��!I��m�ti,��O�j}�+_VAn%f˔�̧>ݺ���W���;���N׼��C{/��n���S���	= ���l���,P!�X����5�!dZp��Y�@[w�?���X���o���+�`�b��;��fE۰��ƀ���b^%&�Z�;�w���P��?L�jT��,?m��e����a=C�!ي���+��DmG\J'���a]$oS~��+ECX#3q%�)bߺ�7x%>�7k���g�¿-I�f���W�I�\NG��������ET��<�M��{��6�To�?"e���,��D�Xg��� /θOɱ�M�"�v���@�߹��}�:���9ϋ0�0�����-O.�ͣL>& o��"tAi�Ñ�6�0���rd��~��̹���g{'��ۦ�D-���;�`X�\��W�G�B���I��A���hkmOZ߰�`���������!�Ԣ�� ٔ��i�,"�7e�]v�Ǵ�=X�<o���G���ͱ���+MpA�{���ø�<gs����<����Ǔ2m�ȝ��g���|%�{q_��8���yi0γ�/���$�g�����^��nε�ݹ��s-��7��r�#�����5�q5k�1�1�wf�X+hk�%!�2���7αV�}XO�5t���庘�(�`а��{�1�Q<��G蚞zͯ���O{�>��c�v7���ō:��!�펵��
H���_���XC�"��*@nSś������|'d!rtpP��ьT��H�A��`=�S	Ē��y�7cm�i�����![Y��e�ߚ�>�5GKzS�w�WW ��+"���Us���B2��8���MP�RT"�Z��>,!X�K0��cm���ϭ�"4Ķ�Ӊr�	���El�}��e���&�F(�{L�����F��R�"9Vm��Y�|�D�z�`;�q�z7�F=nmZ���u��� �1�_,Ҿ�$4\=�EvLW��ێ���=p��/S�J��E�OϢ�{+VhU�����x���Z���Zc��3R�d/`,H�o)7Q��=�����w�c;�� nS/����l�'XȲ����C�昪1�(c�\�WƧ�悅L�<< ��L��i�����0�ҫI;4飁����\Z�y�dm@�Q��d=p��1Vh����?�	�d-p��/�6A[h}���9��J��@ca�n֠��õ0g��jگA�{A�]��dڡ�XE����iN�<.� ���M�CU)kb*��������#�,a� �(�M�%�c��rX)��[ �06&/���ߡ'��H�"����|+��>��B������AN�
��̚l��6���nOZ-�z�y��]ɍ*�<�+����e�&%�b:��.)FE�CC�Z���0s��jǀn`��Z3�r�ہ^�ԭ%�7�+"xqYBe!{�b�q2�#���l.r^�KQ'�{���� ����gMSt������Q\��b�~5��7ŠnS��;�[�[u	o�l͈�7Fa�nބm������4m�g��	b���`2�����x�E#C�oH{�*�R�EW���e1, ��O��sSR�h��AҔ|�bvC��> 6&F�QJ����LH:w@�5�'e޸�i��(*�F�9L��&>���a����}���P���	��^��k�kӾr�;+~s蔷��HX��<k_��g��{3��`����:�9��`��A1$�I~��q]R������-��+�C�8��֚IDF��뙺)��T
���:|���,Ft�~�a� e@�
1���-a�6򵹒���/5-x�8Y�#�����W�A��oGD�Ud��0��M���j��	D��Έ�^]��F� ���i���'����{�v4�w齤"��i��[�%J/x��$�ggq�7�*� ����ok������q;d,��}k��vT��y��ce`�۶6��-���`������j%��7������l	�z�K���a�u�k	��"��z�='aY&Գ�����L�6�Ik")��/�;�Z#�� ����%�JpY!hF�䀴�	:6�,*�sX`B����1��Y8:XW5�����`@{�M�'+W�/ߢ���=�5@N+~a	�U���5���q7Mp�"t�I�_
h����JT���o�8_�R~��
���f[�f�`"w`��'f5�w0�x���y=7;-�����2�k�H�wY;X�~y�)1�"	�b�yN����HA�F�rMV��@�� £�(X��jM�-~Cg��y���vy���D����Z��w�	p�-6�f���3s�����e�M���,-$����M���
��@`}k�-Ѭ��Ix9Z�ѣG"q����p8�B�4(i��b����sJ��_�za�-�S�(}t?-t�5F��w=�:w]|qI��L��]���u�'Vj@��u��zҢG h����L��\{���l?fm�4�zl���&����k��{�Q�Q�>|7(=�|2�0?F���X]*�Ѣ  o$%��*�eY�\����A4_�g9�Dcᦹ��{�����A^Qe~�Z#@)�@�e ,"��l]��tF~�5I����R]C�\��ܚ�bY�ڄ�E v� )�Ԋ�Q�7����2�y"u� c�ܒ�b'��qu�>}c�`���s�m8��y�;��-�nop�mi�f&k��� �Zf�Y08����#%�f�)*i40t(�A�?���EQ�ݬ��S��gZP�M�����rh	�f|�s%Y�ޢz��y6���\�3.���1�ў�\�Ʃ�}���q� O0\݇��O�1�vA�1��{�l<�醱f��󺱠�|S���A��ˀ��8<���ra>�9�og~Ms�lڒS��ZXo�z��+�-��{4GӳE��!�S������2$у��IX�uA3��ĺt�v�Q��M�܏>��5̹�w��sa3�-��*�tC��΀P7XU'�ި'֋�0�(�	�	��#?L��՛�� a�����Oyxv�;�Sk��MfP�F	�0�ׄkƝ�p-nG�5�4��z1��@�<&F����'�!�q�0c�ߙ�&�C@ b*vn��O�P~���5Jύ��sה��o�������M�Z�7w銴Ĺ5y�uP��a-̔KH��י�?�@��Ne��s�VP W��sʢ�|�ho�f��L;�-1_֑~����zh������\��� ����gP_I����J�\I�c|��6��HМR}&�p��s��o~�ݸ=��h����R��^�ב�p�;}���`^ku���Q���+��l�bKڣ�w��	��r~����8�L�c���'��y��.`�=m1�va�5oqԫׇהk(��5N�xs�M}��,cM����҆�� ^ϳ�Q󥚇۴k��V +[�J�V��̡1��r�^�Z,.ʊ���=��5���A��?�����'��`��ޙ���_�X
�����t�u^;��ӹ�B_��ܲ!���W�P���/��z�,kRt��T/8OH0uI0"����>U�7|F��&���؟I�@��4HD"�"�d��()E��CE��x"Sh��ifs0M����mR�6�k���O7�q�Q��|ܠ�Oh�D�!�P�	b�E4)�A���0h��E`^��dn�{��~x�v8���N먼N(�f��!Д��@��%ʚF�vy>���Z �T��e%�_�9�S8�eiy�A�=5ϲQ��(RL*l�DN� )��#b�h��Bl�TT��[��V]ga���\��Q�,�>�	݆��<Q���I������`���C�ø���ڋ� X����ͱ�͘�-}&�>RJ�͋Y�\l
�&��A�`*}U����{_h�l�Da����}Y+���!{]��6I�:��xf ��~�V�*'��~>�����@ke6IL��e�5k�>����s퍓�@���dM�����5�O@�#?]��Ec�^����9���{��ks�c��#h�CP�L���1k���kw��[{����{̎a��z�����=��k��J�ٗpdX��{�{X	��!��!s��v� 5��W粖�+�0�ܛ�!Ȧp�ж�@�q�h�|_���� �6H�5�?9�H�ڰY�g6 �Jb��^�^%�s7�|��Q+B36K��ٓ�.2I�D�W���9� ;Tk��	3Q� ��[̍b�n4)D��Ij�Y�H3H�H��aǬ��A#&TmfRg2u"=#h��vz��`f(5��y,qZ�dB-��)s��P��5��!|S��q;�+����Ñ~H�������LliD�%�
�D��
���J�HF�v
d���`��88�L�����x�� Ϣՙ����CD��<)S��L+8�1��i�yo*��쉒kɻI%�^�Yd�f������ ����p[�d�h�*( �u!ٳG�~��+��A30 �)g�Dr(��E��`z��sĸ�^�Zmc#f��o�|��3���:�6a���bFS�Bͬ@I;̤o�:��:ov��Y�E�;� C��ǩ��2�=�=��U��zJ�ɛ9ͨ����f��K-�Z�Q��hB薙�:@�o�(B-m�r�ɢ���Jx���e6�a��Ƶ'�-��&8�!�z�8����[ �q�NCr��5�`�ŢE�[D#땚�a�yy����4�4��ւ�G�p	.!@���vS.X��t��9�2�p�W�ѫ��e��	J��$����t�X�����ۜ	�]11]�\.�����/\��W��㭛�F[�!
又�yS�b�~��Փ.h�{��#6bFZ�T�9�G[E�q����aM�Z]`�D㳝�����)�Y?��m��A�ё�� f �ŧI����[����:|�cVj
m�$F�0���-�рm'�#�\�.�25�T`T6�%P���M����'�~:�QK�6�ٯa�� �Bh��YT�y�#�����V�y��:}�vf���U	k˹�`�'4.@*7�=(3'�9��,�2L�zزPO��SS�`X45�vh�����=F.��2GaV �ڦE�vJ�e�Hn��VH�r�ϑ`����� +[<�mr.��m^M��#��(GE�`���1`~|O�m�If1LMh�9Y$���xA~��j�tt<��U�agL���L�	�Į������_Q龳�Z��_�Juj��Ř�ѕ�I^��-��+e�`$�� ����?��7^Fd"c�)~P�6�4��ը1�	��i����b�o��iM�ȸ�+�9z�p1�"�]�=_m����)(`L�y�xn��w�w[?�яb]�x@�(��m9�����7�21O[�]P:k7v]�������hn]�T���k�`<5e�ͽ�3X�`��?�1�o��2�.k҆%D�pS��9?Y��z/�'?'�Z�o�qU>��K��i�]�Ugu�W^��((6��=!_Nk��؆J��~R)8K7 k��kUk��k��,) ���y<�����ߡ�5�͵��=����e����O�` � *�ѻ��X��n��Z4��($1RLr��M�H!���f���w�	,����/���s�I����M3T'h��#L��mf2���j�C<&�l�/�1����d� �D8����AZ�7��N����'��˦��(0�n��1"�x��:�Nͽ~���׎�d�9�.�p	��s��5� �5M�_�T�!K��S�/�徆���	��y^�+�؂��"�ey�}>=]�� x=�́)��N�>�B0�<���x衇��bB�l�\�Z�(ں5�M�'ZnFw�g��� �{���� ����ß�@h�.	�A�y+W��\�7����k�ǹ<'�fX��ַC��,�9��Ϲ��ַ���x��K�ߋ>s�&Z̶|��𓕊J��Zx7�־~���x2V'O��2|�k�g�u�B�%���8}�M��]��fgq�Z��*r�u��i�'��P�1>�$H�z�څ���J���>M �T$�T���G�x���+�~.Ɲ�i R�7�ظ�����M�P�z�K��۶1��.��6��Lj�(����oƋ��tβ����F�Ȫޡz��$̤~|�R�ý�1Q�j 7j�9(3"���ŽT��{��|�����p���-�+,��2���k/��f��\BD	�����Z;t
�wi�0�γ��!
��u\�q>��＞���!�-S:��vL��BK���k����β��<�>��,<�����a��,����VL��i"�S��1��%���r�o�{M�ܯ���|lN���Yl���W�B�08��O������a��m��\q_u�yy��潢5X��|�h�&�>����)��!�����gNk�]��8��C�� ,�Ņ�adG�s�kh������Ĺ�> tЪsi��+2�߇�Č�q�:�M8�y��۴����@p
-?��y�N�k��"�a����Zd<�Q��r_�7� hm���S�aL�&�x����Tr�/,�[sJ���_au�}�N�-�o��> hЯ�N�o��q���إ��=v(�y�7h�\G2>�r,�++���r�W�;�0J��N )��h�v�s�
A���T��C�#o���w@�>�-�D:TT��c[�hM���(� b��������v��xq[��:O��t�I����O�ɫ>nfE����@�g�M6�|�{�%�}�����&
K���z�3�`��J($=�����@�x#Ĺ
�z���ɡ�\�صT�w2]��^�h��ւյ�t�5��YJ�}tnSj�
3��f��[03s��D[ж�C;f��={���L�jk����@��>8���U�ɳy��СÇ"���8��&6���,����8�&9 �f9��`�����#8��-�6a��ǀem�	���~^�̞���.���8�2��/�]����@`�_�Z�5GL&/H��k���	6�8�d�4���1���@S��'���Lښ����<;���Vm.Q��E�+U������7/5m�=v�5�2C���e>��\9�:z�X�- ��s?j�� F n��ڣ�c�����5[Yk��8?����̛�Ж������<9�O�R�ڦ��icU�]���,�j9�N�1X�h��^���BF�Uu��sp�a��j�}�	4�73�N3���tJg�FkH�	��2��"�(��v���	�m�|��ġ��w�^�����?Nъ-�[C�x��"IH~���T,$�l�b�Y�6Q{X;��ɸ}�7��
�%��f?k�7jL�A-��Tq�$�m���٬�&H[��U7Ӗ��<7�ônʾ$-�bl�2�6Ǉ�6���=l�
Sn�xm-�\d��;ґ��]��$~d�����C��|��N�"���rKFQ2ߖ�#���� ����3���<�ʦMΡO�p�nN��qq����7�;tL�y�%�%c
@Z$"���:xv�#mYx���2��`�y1�3��+�0����<����X8��vpc�	>��C@b`0S��xs>�#�����Ĥ�6ĽL�~ ��id��Z��V�}��i�:ztP�ב�9�m�j���[_��WNo��t���O�>������aF��4oG�`� I�{�I{�.r��#a='�+��Vl�k8�~i]��ߨ�����O�g�5��z��|oJ��¯%fL,��ښ�r��wjj�3B�{�9;n�����lSH'�%g3Kvf$�gF���^f��o�u	3��IN�����}Wڴ��nL��Y�0��D҆�\���rFu"�Ŀ�"�Y/0�&�2�QNɚ�M���`xQ�m�i���v}��$8?�g����(��C��m�!�����Y��SS5��+,�dXx�am)ٮ�5�%q��O33>�«����J�I1T�]�DĚ��Ѥ^7LL�?����_Gdt�ӓ`6��9Շ�0i@��aҀ���'����) �j0�&/!�_������`�=�p܃>@�T�A+fm3/�܇15�4-G���m�3���t_4ĚGմi^�Ɯ澵X��@?��϶>��ϗ�P~���Y8���7�U ��~�'����?R��	�2� ��ς��'#pk��וi�֎�/�W�N��2�����d�駟
s�<���?��(&O�#���ebr,v�����@������W�\U�r,�;Le�Eխ�p����|h�yE��D���S㻤1����?�+�f[�$�C��1i/ƚ	�bV4���X��f�^ه�rT�M&�Z+�3����%wK�/3E��������.�Zbf�b�m��w'b���&���q�-�y�0�6q�x�h @�^�d��qD��v06�jcs�}2lY�"H�q�ͼt{��
8o?s續�l�9�vi�W����6����ś;�eL�����AKm?a�`��0J+H�6���oMf���w��-��Y��}�"D#�PԜ���
�p��A���Y/R��Pt��>@��ǎ�1��܋k��@�������}�re�M���l%r���]�y�O�e�� }tr5� �^О����7�,#��[DY�\򆮱�Xç-�l�&��ɳ9z���в�L��r�i�� ȧ'ѻ�<�H�D1�R�(_kw�/�`:8$wg�W;K2�^͞5�vP_��WC o�6yv��\R�N��-$����H)�<��\G���bjJB��:F�x"}��~��h�N�^x�y%У��E�/����J��.�����{��HEb�x�'����3/���m�����.�"������m�P��it�@��WF.�\S����i}W|P��5B>��Dꇉ�����Lܵ)�r��a$�_�9��I�!�e���픀ݎ�Ϋ��̸yy�>����6{�7�a����} �a��2W�#�ɢ���ʂ��Р��̜���թ��$��������/����?�\[d^-�'�u���j�!@Y 1A�����6��[���<3�&��?�V\^u����`���9�����۬�cJ$i����f*`d���"LM��lU����s:0�Qz�;F�|	<r����/���[���҈��͝�9u��d#�!�a�>�"��;��5��)Y���d0��62�|�	����wT�������UkS<}���u�]��X��/������gN�8�?�a���oo���"_z�'�K	�̸�OfViS+����=�ݵB��ܽv��҂�����{

Y�4�5-D�r��R�T�����
k�u�]h�w����ﴞ�ǡ%b&��_�� ��y\}F��.tn�K���	�j�m�eK��4>��<�]d�^���ت�cF@��-�x�m�MPCe���ڮ���\,�2AU�Н_A��k#���ESKY���^�y5X�֙�d_ ��������y"�bDuG����_��ݕB�������c�d����D�!["��F�vP`��<�JfP�ҡ��^!�B�O)��e-Fr�lZr*1��� �킦����kZ�S9� FY+r6z���Sܾ/�1��3r4���,�ﭳ�E˽kڭ�r���ͤ=�]a0"W��B�A�9�N��z�?�Ĝ�����0׀ߥ+����-R%�z�L����;[;i 0;Z���hZ���=�5Rh
��6sz'w���� o'I�G�1����7�,�c�F��>55 ���GQq�&њOA2�X���<x,�n�a- �>Bp�N�u���ZK���A?��#��Ťʳ0>�͘4�{�'֨	Ɠ T(����/ ��ƛ�k����}�N�z}9�Ǽ�.YCMv���[Y0������;y~Y��{GQ�(wٯt����HW�n��]n���⵳���zJ�#e��D�ڝE<켢Mϟ�@&�[ȃ�4�홏�'9�7�2��#�M� c	-1����9��}W����zM���WLV�뉨��#���Ñ�uUL�V�-��[M�t����f�f�^ 6axR�@����=��i�>���Z ���g��a 0�)����̻3�k;���,�f�zL,Q�|j-����p���o��`?��G;��~�Ew�~�?�~C���	���[i�1�s�P�Ia�����:~	Q��Ot���t��sl�D �	�:����F�ܶ�h|��M��[�1K)z�4�����ִ���KP-��Ǵ��j��́�D��&��q��,
jC�_��υ��3��o��k�B+�kв	.+�l���V�����瞋ka�h@.���yڮw�w������Sk�-}�A���N���Ï�@  ®�J_��s�<�NiC�!�aȾ�ڢdA;�DU",jݦ��f�] @鿌;%�����q�A��N�t,�5ċ~c�E{����� ����ж#��Y�`��\{���b�R\�[���8�k,y()o��F���Yh�*�MA��Z��	��M���G��/�$
$P�-� \����#!P��v&ȴ�r��M�74n!�uG����s��������@��ۋzo��7����`X�#�L����k01���v$����e0f@I�P�����5g�"gE�Ou�p؇M�R�
�?�$����#UPKScٵ9�"̚ض#R�M�)����Y����w��]�����_����з�� �A�5� K�"�B��������~m���	�Ϙ�)+��dҹv��bJ��b�� ���G&6%X�TH"�2J�KB��{l��8T�f���R'�I6O]oNM�6�Z����������=_\Ӭy�&��0%A�~K�D(�f� 5Gr3���}��}�� xh�D2"h@6yրa�#4�h-
� i3-�DI8�/.�E�8��q�VNS�>v���j�Y�SL��+�u���55�*CC�e����5�zC��;���� ���ǏF//��k_�Z�W�W�|�Y��^~6��0�⇳���g:�po��g��o��<����h@���&X�|;�r���?A3������=�J�T�XX��>̩�3�6W{n,S�_h�4Χ-,~�s����[�s��3�5�J�������E5��E_X=h^�H�5�d����J���u(��}Q�#� �ɓ���~;�L�2���3�,u��S�	@�E��.��үZ;��{���y��v��	�0� ��VbM��F{�	��f��ѡN�f,�������z!��1s�\��b��1����3�n���yYDY�2�Ú�N��g�b�����ٱ3V[��*���5Qk@���Z�5�z����
;BY҆���$�6]5̷5�m
\��i�L�O�ҩ@��"�a��i1_N�ɠ�cX��~�%��͓ʢ! "<�������u��x�q�3k���0$�ƎfiA�>c2��xf��:�u��J?�tay�-�1��������^�8ǴnA�sR�U��mF�#J�?��1ީ�)�����w�^�<��w�c���� ���<R�+�s�[��:���T
kq?~�?�uI�I�׏v�&��E&@e����j�F*Mn�{Xy���sw�_�|� 0y��5��@��cn͚��Z�k����x����� )zY=\���\#,�
m�a�QY��B��əq����"q�^̜k�`E�M�0��H,f ���Hj����F�)M$���,�5#MH*�����Mzډq���\۔`�p��2��"7���y����b��1���H?��d�x24s���c��68X�(�p=@��5�}�k:Ul�-�n�\��2hd(�ى�6A�>�V��|��j�sS�h�W<Wh��]�~�V��L�`�(�:����M�Aδ\[K�+b~�/�yu��t,89Ap�p7�����Zq���/�1�`�}z�i�ch�.� �����c� 6� l���e>�� �uR~����l&��о���$����|� �sm^��z�- ��d��6��#�0?~,R���Ỏ���ߑĞ_�=��k~i�o���|��aSy�Η�y��k�`H/uQ�<8��R8pz)�����W4^��A����4jZ�w����.T��mG�o$m��8�\6��������+nV���E���]�����1�.�����w�7m�������`�lȪ�ѽ�����kٓ�*&��H�����ӏLD�oi�����VH�%�i�	�iMS_�Q�{7L�M/�5��k&���!:���~����}��n��v�uHUF2�y���^y���¶H�N��/6�l�������{񥬱�|MK����>Zr6�qo�f,��ل̯!9�:L��f�B�t���8�n�St�Z��35�"�K��Uk�1��d��-�x}p>�+��iF�z�����J�^I@���}BCx-�~��s���9	�VK�q Bӻ�bL��L~�) ��,3pm" �iU^�<��c�E�K#�zA���1������#yP�k��������u<��Da�x��٧�'Z6�7��?�	,Hd�n��+�kmӰV[��nK�y������00�h~�s%��y=��_����L}Y'x�뎾:B.��@�Ʒl���:`m0d�xT����`\͏ۊQh�i�M�f�jh���M���S۵h�A̓`@�
QV�Yt�FX5��W���NM\���8<A��r[[˾18΃���R��9
�e6ۥ�L��M*9���	v5�u��֔�D������~7�x�H�J�w���G�H!8�Dh}�.�ݺW��H����0�Hkh���0U9���s:�Ό�#�:�}k�f�Mn)�y5�wy�Hv��Վ���}� {����a�b�!T��`�Ȱ��oHP���*E�3��S���#�m�J�hl���dQ�4������͜mʴF��p��۴��s�?�d�w`Hxy��#ɚ9rZ�����AN��s���h�P4��2��Y�%�C��h��m�#G��3������K���힨�F���&1o1f�` #�;t�6H�+��u!�e,L����;�	��5<�߻lXh�W���/�ql�ЮM���e,H`����f�kഒ��3
��`�9[�[����f0�,S?����\���P$����$��.*
���>%�~����i"�)��>��־;|3�Y�?<#ߡI������-��g���w�-ͧ��G˽�gd՟ k;9��P�D'�o�^�F�TEu*���7gb��l���ҍ��f�5�"]m��R�Z��e�\y�/�D��6:L�p��4CZ����ꚹ� �ݜ���`�EX����\�K-�X�a�3~�N�ӅXlN��m���WW�Þ�iL=@���х�3�.ԯz�?�Dw��Rn�H�`o���-H$��R���\A?�|��E{��)���Tk.�:�T���f\���p������=����q.kH\k1Я׌M�h$�Kps r�
�3�w�>p�m���$e%��ͼS^��	]��o��K�G�Dұ~@0 �f� ��8Fێ�6pZ����w[A�y��da�����n-X�!�Fl�y��־����/B�+|0��3��#�%q���TP-h@�C�-А�k���e��h��e+�Js�G����I��h�mm'�햇t��F;ǜW��k[�H���<���D+'c�2*ݰ�}c\цme0�0f�ƹ��Ϳ8��@�[��9]�_�4�q�1�:����@�a�`����5	�����5H���g���_L8�k�7[bB�©O0���f�M&f���l6���.�V3(�m�-�]���>����	����ہ�މ��~�܏Zj���ńc���Ⱥ�W��.-�~h���LҜ5E擱g�(���
́}u53r�* W���Bn
'��o 
�d�+��̹٧:���ۂΓ�#��_�ϟ�,M������v��ɤ)�Z?k�x�k�9U�yF����>��2?���$��M3�hXC.��<~h?|B.�E?\�P�I�2W�~�&��BgN��`]�q9#����s�����5F� <�Ǯ�ս6�g�Ral
�������is%��gځ���>����?�@@k�7{�����`5�3V�B��s\\��^ŋ�5���?��Mo��t'�R������w�n��-�쯳�eSߣG1��H
b��-F���rD�)�cM�6�;�ƙ�X@��=�m`�Rא�7wÀ�����<�~��y]$��Y��7g�/5�R��ENg����q-XZ�RZYt-��:�6	:Q�fV`��s��M�&�Q��h1�6��F�M �3Xm�Ji(��M|;�YZ��[�k! ��Y�(�מ����۩y��<^���Y�H.i`�O~�9g0��Z�$g!ʏ��HC�@�AEd������׆4L�iR�͊%SLJ B��"�O�Q���&'E�T� {0���3�'���2k�+Ax��pU>jM%t�+{P�}P�PBʷ(e�J.�����U֜#x�m������[c�ft@&�_{0����k�c[>��o�gvN���T� �*����$�v�����Q�^_�C�W��Qm�C�Å�i��Օ����О5.ǣ"Z�ڔ���z���р\�ˡ�M֬M�d�8k�W�rQ}�
G��+x0r�d�^�l�la�͛�O:Ҡ��U&5�)�C�1_F �ހ�zI\W"��^P�ƚ�W��n��u����C>�rg�Dɳ�J�����1[(<�M�,Bcb9�B�1���{�ΩĢ��	mg�|��bK��|2f�л��ZS��=j��B�#k�5Z�����'ۗl�	�����,1���xAV���ӡyp�>�>XC� aK�k�KwgF[ﺦQu��23�)[2�%��Q��{fA��۩"
�$u�����r<�C&l/�#����g�6^��a�����,ՙ�v��(,.K|�&��*�`��������V���ց���~����q�H�c:2H����֜�Z��kK�6�E=آ��쩍xAaN�s�8p��s�8��	Zs�T�%�W�)�!��#������L�PXɣf��6�]8���Xz�@H`
������k�ր7�L�k6vܓ���j�ݳ�z� t�f�J0Y	Gk�K3�N�DfF��T�!�nB���}q0�M�6w��:�cS7�}_�3Z�v�b	���>����޹�51��#hF�ԉ�܋�t�V��lK��!��`dH�.	F�����F�a�9�
���'�Ú���j)0;������P}8�{LI�$��C�w	.�)�>�i�<"���Ü��*B��t��\I
����e���?�NP����ͥ��q�x��SO=���ǟ�0�k�E@�c,[����d�V��
:.~�X�I3�DO�3�8�?�y�xz�ynA�������y'�)�>̠=Z�h���a`�Wh�y��#�i��J�31)D�mQ�9Y�4˭� ���t	��H8m��U�����cL�����3�"ϷV�����wRȳ�[Rҵ� `�<�A��t^�4DL�k��w0���3U���b�ЬZc?���Eñ�`��X��f��S65�6��rJ�U�Z �O ��ך�ǣi�{'&��ɝۉ�cه�v+@{k��^6�p2+��6*6[� cCC�iM�O1�tӉ�4��j�on�9�Iz�<�?�<Y��s� "�ɷ����=��>}����,�g���*���VLi�G�I�Z"�p}=}�9v)����b���_���w�G��n��͝\��6�R3�$5V�V|C=�oA<�5A��L��:`&��ӥ�*��0�ܗ�0%�M��;�� Da�Lebna�hM0{al� D�aW�TY�F��m�Is:������3Ё�*����|��bq8,%�=g._m���jߞ��]8$�h��M�} ��
 "�AcB����1ƒ�w$0[�����9�Aߗ��S|��"�:���R俉�`I8�
2ܣm�b��B�m�`1��$d���f-���\`]����0��8 h���`X���6A���X[;��ٽ�vV�|�\#~�V��n�;�ﲂgxV
m��WX���f?54�9���m3*t���F� � R���r���dV��V7�)�J��u�Q��!Ȫ���
����H�al���Peu�b�Z�����U >�KX��^0�0`�wD��vB�������D 2�0
·x8����f�]_�Q�(2��>�ը��9I���ْ�'Xկ�f��	��6ǸSl:��F��n �]c�o���n�'DF���౯ȦRL����E9-��98ұ�r̄�/KKTQb��G�`[�*ø�5l�S.$�SӴ�c��:�=b��ssW��6s'bÒIt��-��5��Ƞۤ�Z�j���,$jSeI�H�/�2�R�ۆh0�G�_���b�o�����\��g�}6�]2�\8d��}h��t
X�6�����A/��a:0��s96;;��WQz:�# �ҥ�a�P1gqn��of�HP�Q��bՀ!��_�<�z��Zo�
�4���\�M�P^�
���4��)4v4��7/��"�<�2���3��>-P��U�"��'��㠣�5�O=�t��'�j�wϽ�i	鬡�`�/��^ao�>C�H�v�	��9�f��KX\�>}"D�)I��|̓=���q������ט��y����T�ET�5c���S	?;C�o��;[�>0w����P����[�Rٱ����
�O�KxX��:��"Z>����P��W�c�� �����~CBH�8Ý��t�2���,�82�mw�h��l���Ae��n!LF�$8�I��7d�LT�t��`�Ln�kc�y6H���	��bLQ^�y�6�w����W�_PKt�Z-y��e�sQ���3�B�Yė$��&�5U\w@>C>GUd��A����*{�QZ~�+����4����WF��U)=���)[ǂ>���Hk=�-`�R���JK�d�"� ���4d�ǁ	�Y�Q�a1@��w�_��]3����LԦ�x�̡E뱶��LN$t�3��I� �>4iMG���9� �|���O��.,�Xo���k�߼�	�]X7h��G��9�4��tD����~���/ǉv�Z ���C�ե��.+a~L%ÅA-6u�W��}���v^"rX6`��� �2�p�t�z���o�X�7���� ��ڔ�<^��H�K�A
�٧|�����t��DO��O�N]��Z�N�b��N|zo\�sv�.}w:`XP>v��KV�	 ���.�Z��[���`�%�8��!w���:��=�[;8�ڗ_yS��!�ܵY�kwB�PI����dX�~�qxB�Y!y1@y��B�p�z@����>�'Yo�O�i0��8�&/l���xQx�Y�,^3F���>�q��XkQ�i��3��g �u����۷B���C����6�4�5�h��ӟM���_��kAd�����k���;M��mG�v��m�|�3�%d1,y�ik$���e�2$��E�~��9�+��ET3�c����W��2g����=@H_�?���(�i��֌�@���uL"q#w'�ä��]�aR���h7B��j��˂�����\��,;4���*�ۚK�%A#�/c�;8ϯ}y��&�y��N,qܡ�.K�T��K�1��!|e��2�e�L'�A$��/�u��L��Q-H � l�!��Q�<Llk+Ҿ{|�
�@�bƅ�2Uʑ�!��Z��WLa���s2gI7Q��dSG�� '*�]�) ��3��"Ļ= �֥�K��F�R����Oy���mY螶(�5�Lj�����������
�����/�é-�\�n���Qb��ޏ��.���5�df,�zfne� �eCm�8 ����]���6�1`L.k�"O��8��sH�	�p��� `�,�]���$�m�=)���F�mT��c0`�s2�a�3L�)Ѷ�#Y��6�>`,q֦�Z��n�jP�-q���?��!t���E�Q���z��/�f��4�s9r44��I�7;rð1�LH�?��OC��.J{-������@	sXӤ��?��G{$X����үdp�H��ܲյt��a(��zVjv싦XR�/��H}I���	 �7��F8XG�#X!��	��@��<Xc�'�t*8%I�c�J�Bj�Z�Ae�x�F��@��tb�u������q��qg�E� �������>��H��$� ��I�����N���j��u�v#����X +�Qo
5���-(%�J+ߟ�%=�Vi_�3��(���(�u���I� �S=*-z\��N��.�!���{���O}����U�%E������h��bg�Aq��'Qce\���Ф��"P�-��n���:��C�� �������Z��G���������,@���^l�O~鵞��^��$ hI!���oEg:�j���]�C\����hX1w���FP�v�=�l� ���`�� ���aV����o���;�����F�{Y:�z&��"���*���<�5�}W-�YC��8q�vk�l�t����&� ��v=	�Z�?w;���y�����7f�<~��
�?�ݽu�L��fT�M)��*m`&�I����Ά��mX�	�����N	�HW|
D`�*/h`�?Iii��TW�T��l�����_g>]�{�Qf���#X5��:@���nt$�l�ea�y����n�XeY��Z������;��u]8��2"y	�pP�5�f?|�n��g@a:fD�]�s��f�u���k���K"����a-�ã�F<�	�30􉹍�_G`]D6S�Ro��zѯyůJ��̽~�q�A.,�!�������;�)��L�=���޺{�������O=���"U��!Ea�,�5�9���a�`N|��x���(3��!��]�|��s�?�_����,T�E܉Fw�{MGX�w]���!�I���R'hW��m�Lh�C .�m��TlF�8��EDÛ����o����!4�=��I���ca������c@�a�d)�a�5(5�ЎV��lKwN��l�8�Q[[����{YZ]#߱�|.�a|\>��䵸ؓ��,-+'F~��c1P2g�ȸz���5����F�����oy���y�|�B�f��I-:s�0�y;J��Ŏ��c�����O�d$o qR�>7K?�e���# �]�ӷ������w$yV�[�$ 3��W���L�0������2�ʰ!_/�����������KH�,<��f��k-�Y�:n���P�3G�c���
������	i7f�5�����y�/qj�)�ee�$X`�DS��`��Vf\�|;�қs;6�o�j�ͬv��$f�N.J�D�`I�߁)Y�$�����u%��	 h��SP*��M��W��d<+ڪ�i���Z�0�O�����bh�?�s?�v? ~��ьm( �:��i�pr��+��b�w�r�5�x8z��٧�g����{��(�4�w�j0ދUb'Z�����y~7�A��������N��%c��3v��&Q����w���CЮSt���h���{�b^W#���җ��QO�^2	"�0R��wLSP2f�u
i�/´!B ,����*V�\�q0�Q��;�����0�y � )�h�"�H�|�w�"
;R&��S����ELj��M��~$D��@�� ���jB�3\�؍&�&���2�d��cM o"���s3�����뎏����sg��ۧN����� H�@K�|�F��GsAaϧ�������!�%�=��)� ��Q�4p&���.dߌ��h�'�|���jA��9k�<�5^`f��VTl�Q��p��Sj�kN�. ^��Ƿ��+��}"������h��2�=`��6 `IX�zGҗm��S����۴��Tʸ�2�q��9��OG��0� %��m��̮^U��s����pcȔ�}�=�����/hw�7^E�E�ߤ��> �m�uQ��.
�U�^�o�d�����׿�%m���h�.`���9K���lZwŔ��b_���П�N�(�W^}M �R>w�yW�G|�φY4�!s9aĢ7�뎈���Q�`��iwh �2�*��a�֞�f1�q���Ka)c��f�vc�Lh���ü�ۤ�k�wD�mεoۦ�uSY@��0K�C5�ۇX�R d�WyN�g}0&��`yº���j���n����M���Gg���Iy��4�� ��E�v�s ��0kE��rQf�ۓ�&U����R���mɐ�@ r���	��8D�	���$��/B�)���$Dk�M�7C�{��U	��[�n�fӖ�G������Τ�9cg��*��"���J�o�!A$C�a�gC�'��c̹D5:9�U�!~�>�~8�	f��Y^��� ���44��D������m�Hrv�6�h�ʌb?��֋� �e���Ƕ��b�<�,���na~5gij�j���_���"��_m0,@�+ �V�B`��3zف3���z2m�s�g�������	qn.�J`6����&g�0�ZfoG��� I�T�!��ԩ7c<Oj�|p�9�
R�A3\�'�C2mcV�t9(0I��oha�ϰ�r渘Z�РC�����ZG��"Ax�ܶ`����7�<�KX0>��϶~��^���D��_����:}ǅG鯘����w|vxW*��؉��ҵ�
�8���?3/��k�W��5-�wE�o;����-4�j�NK�y9[5e_���k����2��3x���(�St%���:D��%��}�X �na�;�p��YxEN.&K�9A�f�Y�9������дً6���	#�y\]�~#�mX���g�C�9׌Ҧ4��wOL
�I�R������1x�v�ܻ��rZ۬WI�������+	���1��ܟ�x�,fR�S�Z#�G��\����9`!�u�%.�̽M6��KrW���5�l겏��k�=ΥM��X&��^���L�UG�l�e���� �&M9����6u��pU�S�9G���#�Ûc� �H�p�+���:�S��2ߘ�i�B�������rTiz�ܑ���2����2k%��bzG��
������Y�V3��V�m�#jY�� ��^��F� lv�x�g�l�X�h�)@[!�C�ˋ����<��l�hjJ׾B�F�,
�A�-�'�3jG�iH�{@�8�N�-9ɰ�VRA�H����94��W��grN
��m�Szr�2��ż��W�Qb��@�� ��!	%kgac�ghw1��	����M=~+REަ��o�ҟ�Dh´����d�1X�^��#R��)4%�����G�&�����8-Q�v���1�T�@�	�fR!�G���&m�b���Sjb���������$yC�H�T�f%��\a�h���&�0�0{j�t�Y"�D���S�ssSR�Ə�lV�_���o�2%��V���>��Z4���<5
���2U�À:��Zx֖�p[a)>�~2Ϭbīi%0�X#��9�AǕ�Pϟ�͠���;(��8��qޖM����^������+�g�2
0����ܹFf�	�I�Z��������]I�$p�4���Ks��&���� ͤ�6�y��$v�GI�xS@ȳ߬��?�p�B�~�6�����`Wݦ����������� ��=\-�-U�]-����F���L6������X������3�;|!�1t�v-|y+9���H�y�`J[�^;�F��gڷ��7�p{��N3A�%쐃��� _&Sc�����E3?O\Hb�΅h-M�y�ҽkQ:�������
1��63������!��^5���n��P8���� �a=�G�4W��h��ˈ
�b�en`Rq��a��8�� P�C�@����bȲhTIs����AY̾3-�ڡ�\K�K�F̝3�8�>��՚��׋8�7*����a�]{iXP۪%�s�5P�ϵ���^3��N:E�6׼��55�|��gf>А��9�k��������p��ƘoA 	�;��۫���p��L�Q1�4���ʨ�J!�=��
�Qj��&Ջ�PM��烇��D���]XصF�Z��g_ә3oE?x��֣�=� ��h�^�d8��hE+�}�3xσA�k�s�O��us�j^c~P�F�ݱ-�o�O�[�7��v@�uT��@hm�($�g��g���ײ#�����I\C�������OvM���mA�lM7�Vs��ѩ�[�n�ir�B��es�%�|؎y������w;NF��'H��F�7k��o�7�L��gS�3�zAzq�w�v��E�9�נ�H��G��1��c�Il>��n �ZIm~��x���w��� b 	0��� G4A��M���M]���W_��Ι�FT))	|Y�W����a�;@ias�i:�*	v�T0bq�Z�5Hx�=�� Îo/ǂ`�*��2_�4��	�A���Y�k&��,������Yo2aәMx>��}?�2����
/�Ǽ0F����k�5p�~�C��Ϛ�M�.��ܱ�``h������R�BN�Av
�+@F�z��K�����%��CC�[�Ϯ���N��!�����`
%:���1�>%��g>� A���ӟ���Y `��gY��n���p�fka� � ���^W���2��(砧*�t;�������xL�����B*�:�@��D ��γ����7]ٚc�Zb�LzSt;����@�βӜ&MA��&{Q����nJ[��n�<K�U5e�L�6-0�����T��j�b&Qk��զ3�3a~��Cڰ�x�v��kt�/<��M<�"��Wh�$�����N����WK�<�i�~�����Z3���Rm��0�~ 5k=f�3o3�=�����B���l����x��ީ��-��G�7�e�r{(��c�T��xV���i�11�+��&+/3r#P!�=�4mF��t�i�������K3�i��$wk�n��צk��9���Ęe���L�O�;t�2{�p�?���m¤ ����1ެ�+:���)��6Um���E�T�����4<�d־Ү�B�Mi^S܃>:���i6]Dz�ʦ����Ԧ�$�C��t�{z};��¨�Z d��*(S�czs�q��MS��^�{[�4��&��yӆi`7���]6��n�1]��ga�َ-�E�ʕ�*�Q~c�mFf\����A3�+,=%jC�ݒ��ƚF5�kjtF؎�%L3��Z���k��3%HB�I2����"�Yž�(�U|�5���+25{�	3k~��0)���'}aq���o{�����hI�h5�z\�"*2���;B��s=`��4���B������,��( s��0���A�#�F���5�x����F0̡ ࠂt��[3���Xb[�N^�%j d�m��ϫ^��ۋ_;��m�Vb�:ƴL�����M��1,�#�Sr
�2�LZS^���g�i�A c��B��=w��po ��{��,f���FN� �����s�=��#��]a����	c���z�Z���w[WU�{IU�&'�Z���b��SzeW����DioN
�~�D̮j��N@���
-k�B��N��_��2�������
A@O<�#*�MzO�/��9�<j!�s�'������^Ӟ���Iu��v�z70�^k��Y��������p�&�tmm���$>��S��yN*+^���=�K�\�|��T�XO�B�̍�Q1�fO�v�S-�4��3�&@�	�%�<j[��	�N[0�a>���tn�D#Mx���މ�5��K䴞��;�k�ǌ����{�!��}��wMK���K���7���j�M�d'�����^	��I�D��!�C-L���ʹ�H��wmǚ9�!��xe梤E1C^(Ӥy �*��-�H����T��C��4��UY� �n��(�q(h"}��70JPU��UT�۫^75#�A��S)  :���X�.AWWG�vߚI6�����&�5$�:��%o�P3lÄ��s�fo� <Yw $ccc`rG]B��a��d[��ك"��\�Kg���J�a+U"eƂ`cA��;2�n��r@!m�𤶍�w^�/+�8��-W�b�nMﵵ���c��dm��8�en��>�c�'��:аIOM���s�.� �����x���lj��y�5]��yr^�Tс�М���\�k�Z3�7mB[X$l,K[���=4wƷc��nH�z��I�M��F�[�z��Ơ��k�t�_KΖ�o��l�$�ݒ����B��2��l�<K=��m��g���A7i�̇8k�Ϧ��7簨a�	�&���ejb�^ �f��p�^�����My�悴��`�y!��*��� r�����f!���0"M�X�?)���/�>3�[���;\Y���R���-���TL�l\���\���E[AQ�hB��m �oK5�C*�
6�f8I�e��2b/7<,�g�M3�,��3��c�"̀�M�m+������sp�����6@I3h��30o̗���J�TJ[��s=�}�sJ��W��R���O^�I���|��Լ�+�?x.�v: ��4����򂿗��M�W�Š!���NBu_�	���E��Y��������;��c�{ｧ���|�I��H�h��U%�0�ds׎v��X^V�N��T��a�mFu?m=	:a�t�$=�؅V,��s��7����Ľn��{s]�}��B�Z���ܘ[�j����!Hg�-cd�y7�c��~8���o�5�%L�:��"�e�F�L��W뉾>��R�V�-4CA��~�Vt�~�	1�v��a"�XJ����5��gw��Dk	΄Q%�L��F4�FZ����h�̕��F��޽�Sk��� ����RQ����$��`T$�J	��N�ܮQ�8<|{h#�.e�o�/�Ӫb3wU;:,�҄��a^���t�]�6��?�����Ϣ33���7h$���Y�-�5
"����$U�3��2�!A����
[�q�7k
�gS��4^��<M@������� =V�n?�b󢅚؄Y�y���h�D��}�{�h�ܫ2�&�� ��D�N�O�:���ވL����ȶ]	P��2���2]y�2�0�Q�p�	PyP ��ONjs��3��~]�1[,��?�@��+j�i=W\}��i�����m�r'�6�&X^�ۅ���L�kdm����m���y�"�X�~�4m�K�E���  �s6x:2��=4�=8�k �"u@���1�y��5�K�� �`�d�����[�nǶ��]����d$�M�g��d��~3Ú)&�L�v�&��W>m6�P��y���W��˱mޫ�	/"�k�I��H��W���C��f��K�|P�a���X ���Y��H��,���2�ù�WTfI�z�g�����ⵉ�����ܤ�䮉َ����Q����x���>�c�� �
���kKܦ?{=���L�� O�7�l35�0����)���o�=�A�.�����,��j!�y�>ޏ� �sb\�����nQT�"���`����+�/�`���*�Я�x�H==Y^ͻ��s�1o*M�?�񏷾��/F1m�7�K��糩	Y#��ڪ- ��ե��ozvr��Dn7 ���s��Tu$��Ě~�;vZ�M!{�=׎i������OцM���q�`i�����c�4��v��y�i9�"\�*/[�j!ü�{q�	jݯ�����\�=�vBu�0�p�ns�v]����Z�ܹf*5�01�0��k�����a��{Ky�F,m�i�ܿ0MJ���%6M>�=m������4G�	�;�֍=�s����q?+Ǒ�!vvQ��h�d�͟OL�����n��~�_�t�&E!�&s�(�uu����>��Ef3��!c�1�3Qd=5�4�S�}�wt�*�	1nÀ���AS1�Y��(���p�^�����m�C�ƌ�<�`�9�h�'>y17��}�qW�H��l�@a� �WU���|�/�<�H�����~���Q�)�T���^4�Ui��+��y��e��r�b(0p�*�^[l�6�[P401�a��ӧ�}�sQA�4�,�H]�L��ڪ��:�s}k����؂��p�0�N�����0���1I��}�5���N4B�i��kü��b��^2��cPW��k�O�F��:k�;G���[��JD����@#TW�f:��B=�J�Ǿ���u���X l2�d�X��a;h��o��C�n!�m��ܚ1�@�,G�qnGs� ��}�S����f�<�w���9�����j 4q���� %F���!8�
���7���)�w�}1�.���?{��e�u��n�2
9`&EJ��VK�(u�m{��=�l��;���{� #@ܿ��j�)�A�A ��}�9׻�:�N�N
 �����^k�ޙ`Ƨ�ȧ�L��>�X���b跃��I��=$��UE��׹c��vƛ���{���@�~�dj��p/E��k��t��A��)�,��}!cfce�5
]#� |g�{2���`JLh��-� �8ƃ�e=�&���j�kM�e�ݝ���M0�0(�ﴙ5E}Ψ�z�j��c�$�N�:�U��iD ������R�q��<]�Q5*�}�?��<<�̳�MK�HV�w'y�ym<c�gP���j��J�]&�xt��l��g-�	!׬�e�z��il��j��՜���c�<�0���B������P�؟�J����uge�[�uC�����B��+�3�Mrs
�q/��!��n~�m�� ��q���������d9݇t| ��Pj�l��f~�"K����cA�8�Bpn�mg�5�Em�M�"[�Nמ����ZlLC����uX�����X��f �w��k��Xf�5ܜ�0�T'@��A������$G��� ~4�3g�6O>�t[
,x"8�,s;k��h�<so_�3Ӊ�+�1,P��F0K���sM*�r�L�A-f�^�	��6��_?���m"Q
8�m��ɜ�ڀ�b��#�t9���2���
t�߶fX��g�����3̡��`�p�B��;�}'�C�� ?myTMw��e�,�I3�s4p&@mB�M�F�	�Z{QY�j�ɗ���(�M򸙳�9��}o�`��O��~>g�ws����>l��[[A�|��/Ћ�ϰ�3߹�����d���_�y����ЌQ���{�|�����Z���}�����9Ful�1>��x�ӄ���04���<P�7���uP��︤��3V����8�S)�"�qv��Ҝ�)u���*˄����N��O��z��Hw�7a8���oo�`k��dmG[5�	�5��C����e��a����� �0�6@�t/�?�	���,�}��
N���di��	�T rk�@r04�'ޓ�f�'�P�9�LǃE5�]S���)�<fZ�ǘI9`�����/�%amc,Sa�J�m�,+Af��b����kL``�e���$$���V\h!��>0r��$���M������qs]��}Y�e.\	ȩV���c-T�:���r`�,�w��fi�6)�->B��eERt��S�ȉ�����k�yK��.�3Qzd2�����Q��0�K/}������Y7���yY)�:{�u�v��o���]-�~�t����5g%�k��qvLi�BZu`U��K���a��B�oH����336�Q$B�ma�w�� AH@��ֺ��Iiк��}������l�)Sof����%Ḋ�p�,kTAH��F�G�[���)0�1$i���ʹ�21L�m�����1.��o8�sk���A0��Ӌ߹w�R����R�7���{]�G��Zs���2��I]��С��Ec�$"��a���:����'�mNz����p��ӧ�oR4�e"J�+[Yymt��=iy�/�}0�NŨiē�<
�>Ê+�m�Ř:k���0�q'�&��q�k�0q���^{��l� �Bc\ ~R���o����L�&c�}5��{�y�΂�y���`l��h-DYÂ���8
���b'��j<KKYkrM�{����&c#0c��3�x��!����?���@�C�� �)�rg�(���ux~m��<7Vrk4��p=�>oWD��c	8<!v���H*]".�����=�_��Ih�$�ؚ��r�٬��Io��~��nE�	k-�B#��4h�"ʛ������%f`C?��� $
a8J���w�1�Z��s�LD&�<1��7K�m_�c(��X��
���f���^탺�h��u}}G[H�F��l�Ga�����=�B b�to�L�N_*�}����-	��!��oߚk�~j1�?~4� ?9�@vW�]i�]���%�qY�C�	���F�5=}D��.����Pe0�\�\�,��{��^so!�B4�[=O)x�gd��ts�fxn�l����G�h�����g���\�f��s�΍>0�S�&��v�!H|<���QyVG�:�(��u7z�I�I)>�����tAr�$5d%(IIɼ�,�/�q;g	���U��0�	b@�A�A.e��x-�����Y��V�S��3#D5�����`%?J߉Js��];��N)��(���i�]w��/;v��1�D�v]K�ViV�wEt��k�7?�����"���\��KJyz��kRt��i%�.(����lו�L{\�����zmS�~W���h�"���u�%�xC�/�⩵C���e�&�[�����2���{�Mb�)��VI�1I�0.Z��Q͜VC��{-3�	,���"j��+hL�#�����n456�uQ�ذ��s   IDATV�	�0�9h�@�`���m/c2D�ZE�y�E!��4��[�K�̴h���-�o�ae?���x����3�X��(Dp�:2.!G���2���gt��W����m�  �!�:���ϟh�]x����'���o�Oa:�l�F*�uh\e�HY(��+�yb"�U��>���k�@J�ڊΟ�Ծc���;Q�����|_8��;i�q>�`�)5vmE��ڵ벌?�ϫ�:���ЩiAf09�k��>??ז�JKs��9���E�p?���A	��e���߾�4�Y���%��M	��Rf��*�g�POA��n��5%��X�z�y�%M��27k����P��?�>E�kv7�L����;���o��'�o���כ��?&�&*�h����A>��(g��z��"{�6X}Z���<V�x�n�a�]���9#ރ"�_M~Q[�<#���W[�2��S�"�I�.��t0�>�S�j�+,��GYɾ�/������<6˛��4���:�q��������G?����;Fn
�̪��B�����QW�E��.,k�h��hk�gu�<�c8��	�ta����]����9�'�4� �����vA����b��`+z،.��Ԭ�y�hgcZ$ZO�\!�ml�֬�0'<OM5���hI$��������!XC���2t}�N %<r�Z��(� �����d�}x'a�:�&��3��Ƌ��@�H��6��`��:��	���7��V�Z��+8cA�H�ۀ���E%ޔQ+%ϼX%1W��>��$�_�u7t�	���O�*��������<���|�����o�%�r+'&�3�$z�rtM�[�n�ҁr�ɋ���6�;���2��x���7ߌ W���#�q�M٦i���`�p!H E�ڮ��}�(�i����J%�Z�)�|"(y�Y��g?�y<'�����v�y�d3��t��ͦ{�Am�����=�6/%�R�g-�P����������ncJ�c�b���AQP����g�{�О\���X�Y��aR|�X�'9�}s��pOD����
)|�|�7o7Ӣ����\�� _0�����h�ƾL=1��(f���9���߁�d�.�a���6�Թ���A��7$�6 (�����Z�dޏz��>�n͜�Y*bB�����>2AY;33�ҋ�6+L˾�����N��چFj�/#+z���ю-�zNؒ��td�Ж��1�����?���Q�-z����c��h�*�`�I!d֫���'�5�*$�#��6���5�[?C- ��5���l�u�s�JB��Pr��j���
l5�(�;a^��x?��"lg���y���Z�ks_�Yp-�(�>�97̊kp\�~t\�R�O������Y�}����e���*�3�%�?�2J�#�Q���2�Zg��k%����B9-�Bc�]b�V�|���Fi�M���MN��[�Н��{U�+�����0����^����_�4$�wM�Ç�o�@z�i��]��T�b�9zs=P�����z�; ��K�x�qc�9k���Fi�8Γ��)a8&���B��ht7�h����	A��Op�Q�M+�S���6q�x^X`6�M�ݷ39>���p�t�&�@�s32o Otp���~�zD��NC�$0��k�>V�y�񮠂>#X�g���x6�^X2�}���M����-@�f2|o7����S�ҷh�T3����6�.n��x6[�	�f*B��f"���J$3/���i0_��DYH����q�%s�y�W8a|FG		�0�i��
8��|�"�"L90�����g�t�u��\L�
@��^ ��9@Xc�"��c���+}M�%���A�����|� {�̯�
�!lZ�C��0D���qp^���
u�g_����I=�zXN����.��t�u��k���
 )-�	]W�G�c�S�������&���C�����B����Z�>���:���c���a�3�C�v��8N�������Ǎd����P���{~a��d�8
�L�՜
Tٷ��dFXo*�^��~CAh�7���3��>����W$n��=��s�����C颞{�f���%�0�h�h����4p�1��gN��0P�"ѥl$`���?�M�z�@��¬���8���a��R[��=q<�֖V�oYc��Y��@ 9�0m�&b���d,u� �y]��Z�*&��+�1�yw������<׎�s�s��IC���	�Ss�}��sL�$D�H�Q�':� ��Z��xM�����m�E+Q ���(Q����DRO�pf%x?���S}�}?�4ѷ
s�RVJ��T��`1rT��sU�T�0���>C�aї�_a�)`��X�t?	$����c��>\�'ֈx�%����?eeҊ?��K�F+��3��(�F[�Qn$��bN9qD3c�w���y�.�R��D�����L����]=ĺ�^Z������/@��'�b�
˫��3tc�HO�o4�M(�Z�����}}š��+�6��$��"[�d6��!�� �i�7l^ke$���-q8L9������DL���X0X0p6
��7ڪ�>#�GWrӜ<IjŹ晧��/���'|�nX�0U�w�W�Noob���טX2��V�LG5}��I�̍�.�9���l��8����=	� ��}�hjJ�f�27<UV��w�}/J��9�H���0��1d��S0�=�9�K��)����B֜8 $,���Eh.)L��[���������A{X�C�?��?j+�ؿַ��:���y���^�����-=C}���=��F�j�aaXW����}4���q��ҢL>���>�r`���֛`&�w�/B�,!x��歷�􈟵��Q1�e��x�{1��!{�b���`hҹ��Tϵ�^����~]��㄄��}C�>��Q�&	�@��I�G`=�s�VT_�0��SX�؆��Z֌�c��Qo4_��d}r����ps�c�n$yM�g�͝����7�ÜǇ}�>�����cM`�l�i�Q��T�+������5f%� �h�D��������N*�ub/V�O�FXwӄi�� ��2$�F��RŏUk���CK�#�m&J��g�#�gL��%�ds�u\��"��02B��8�V�+�DA�"/�Y�9z+�%�K1�(�vXG%T>Q��r��ul��b�K�칣
�����|^zVK@Z�W����E�웴۱Vn_�����1�V��`%�d��~�m�5�I:���X�>��GFgх�A|!	��Ie���7��m�K�H���k����<�k�I޴�{H��a�}I�#:����4o��h2����q�Ʈ<c%4k��^-y�d7h�?�P7���m���;i����t�0,�yq[�x�J�a,L�L��uI�:@��0���	���+7G��B��%��VO] �z�b*c��y@S�H]�f��ֈ��c7�ue��@��M�yrt`xL��hvW?�p�[O����#����}���.ah����U-P����k �(��~��Q��ЦI
��;��knI��2��cE��'�p&�$�]�9B�}��i)�6fNp�Z���*,awMXwW`����&���B	
b�>�,��7�C�H	H+q�Z�w��i���Nǚ�_jW�8O�����)@������9@�{_���ۧ�q8 ���5�de�>�ZX����&���?�B&h�\��G���T��.!�n�'�\�|�I��.w疚7�H���e�JW#�Җ�]v��Īԛ���e}�钖#����@�vEؗͺ�+��D���1@wz�-�m�&X�P7�G8����d�l�{bKD�d3����E����ak�I������p�V��X�̴�;�@�r��g'T�2^�OB��^[�aMTP7�s��a��yK��d� x�{�	=:+Ax4�������r|�;��@G,"�:F���\��p����N�ɠ��J�-G~:h`ll6-$�;a0�Z�1V,X#.��8`BƏB��#�hU�ʡ�=r������x�9��=7��F��X�� F�KWw��o9�{&�,�.��tOx�hߦ�T5R��^���B��2:�zP9i�P�jC�S����*u)�q�P�����e����Qj�2��[�O�����E:����J�W��u�NBRH5�(��,�Hg[��\���4���5�;c$GmND N�؇����ۂ����Cpz���B6��y{Yڑ�et3�d�� ��yS�P���;���0-�|<����K�}!M��b�8	-�3V_�p����y0S�s3�$��U^>�Wn�L�G@fk�Z�5���e�n:���|{���y�(3���1>H�l����8jAX�Xx[f9��4O+�cR�ȸ�`֚c���:�<D�����׌�ߖ?��sW�@��_�@�:07|'�%���$�� *?[�$� �*7�ތ~}�����|�kแ��;s�T[}%��%<K���ϕ`���t���g~r}��2A��L��E�>�ǽ��H=F���Cc��$�����Q�@�F��=�>���<���'�L�����������E��B��z�[C�V0=w�"U���Q{�W5*f^gz��(|����Z�Q�������y��<�h?�8P4����h#�+/�hP��H�I8Z�����O.	����o�P����w����E')@X���<%�4�:�tl(�(��DElZ�%�Vf�N��"|�?�������xv�q4���s���Y��W���9v$A���������Z�5���LD}b����ER�E��m�?0K:e�A�l>߰�#���j?b��h]��R�'��q�od3��柶2��R5���=��Uw`2���7�ܢ�Dm�տ�����Z~�"±־�؊��%|�X��|v����'�zz����0iv�H�[�9�6L���}.2���4���6PJ���¥B�#������Y���	Bx�LbB|}/����:l�P(��\�;�ѩ��&���*US8�E��k 8[塜뮯�1^��8��!�
�.��u:�uy/G���87������v��'�s�fͻ���#je��#-�&��/�����ּÿ۰�y����-��+|8ۡ��ܹ���4Щ���>#p�ם;wJ
Λ
�zW��;���'\�xYwE�PA4[t�gV�G������Z��/$B�s����]�g�<��=�J4�=�!:�;���F�[�b�����b�Lq�E�/��y�0�W��2ZԋXo�c��gض�"lf��@&�zSڜ�:X_�RZY�4�qm��oX�-wU8<�z\5O;]����5⃺�>}-݂���r�`4�����](_�B ᇣaS�Z�wn4/.?/��K��� @~��K�.�g@��M�Wy�6Kɸ�^Q@A����,V�Z�d+�/��Ǳ ��f)S� ��������;w6*��;�Yw�@�s?�R3l��s<��l:��H��B��@F
��L� �&������wm����L�@��؋�!A��6�A�a,XB�+DVL#��M��~�/kz�8�F�P�	��z�{n"�D����e+xQ�����'3��Ъ�ԥ����H]@��R�+��~���~��o��ܾ��*G�R0.��q�E�Ƹ
(|^
>� 㴱��m�:���k������ ������*R�5�C�q=\P�",�tm�Ԟ;%�drsdU���ڍc3��Ќ�����/�;�u���F�3�Bm[�AѼ�]n׶Ff߄}G�c�YD����~�7!�E��]���<��a��M���[�,��:5d@��{�z�j(n�Ƽ�����a�V͸jd�>��8�04`1�ҷ��Z�4��[����А�mX;n�4��_��NDˑ����{� 8k,�?��X�ّG��t����X�ڣ;V�����0��ҽ�C0 ����㏵����"��(]tRh^�n��x���ˋqp�cx.,1����pN���W	�=��a}�������Z X���6V��EA�|��/_���v��o�6��u�J+E��֡3�<i���~1�֖�g�P��1 x��qy�w�,ײRd��~o+}��e�Ѻ�yn��Ҕo,��%��jt���E�(�ߛo��T�_4��?R�7#�V�b���a�U_2�/����|���)f-�6�ҿ��şQ���3�}|��>�4�g��`�ߎ^��0�5Qh�݊h`I�L�(7�X!�k2��R�2i���5�Z��3H�n�l�ن�w;��_��{�w=�O��=���>�bY@���X@�s9sm�����e�⸃�"l�h�����{��rE��5j���gkv���'��o�z��	ښ�j��?�(�3�I��0w��d�`T�?��Gl�(,��`�Ԫ$'���a
DV�:u2�n2��=k������:�{b�ѾB�I+��'���Y��-@tc%���4Nh�]3�R}#�����eK�,���R�\��	S�GE�C�q/G�^V�I��?�"26|�0I	2��RQ���@�^;3�V	�t#�UƦ�"��٢\�`7c~�W"H�ri�/�\״��h-Xq��c7>��.��t�M�9g�܂)}�]Ҹy_�����3[���l%ִ͸lxdq��a��7��2X��Y�j�mi��֛o7��������#"A�U�(R�x#��3���n�r,c"6մ��fL,�p71H������� ����� �n���ސ.��b$��[h����@F��"ΕHvÞs�������޷�	�D��,�C�]~Ƀ�"���Z}M8{a�!h0�{�B�v�d���5^o��B�Ｘ�j���h�X>��+�:���㾇[%u���q���p�^��Q>v'k��|7Z��ة*��! �0������iVvPr�	���c��-�X#,$��ٲ6��|T�E��U�K��}�fH}��g����0��g��d�L��!H�w?��C�s+�#2�������} |(�dN�A�
�c�q\�KPϕ��42�MJ����¢�	�eJ"@��Ҙ)��|G�)
�ߤ[�`E���X��a������^�~ϵ�q��Ѱ��Wú����׉�_[����W��<�W�MT�A�.L�koYV#-�~��?i^��w����J��T��M����4 �(>\�օ��=�'�@���Xvb����p�K�:�t
�Q8>sC�cIa[�ƨ�{��ȂP�tM�~�NM~¨�0 G�9��B̃ ćqMÖ�|Q�� ���6Z��+G0����O�5mq��-_���z��J�0K�a�ͣp���4ð�`�Ì����60�퉓G�T�B� p��������=~C�hk��������h,���P�
�t&am9r�-@a��6,5ޮ�A�d-x^�B�s�?��i��AW�`�8>�J�o����eU�������((m�g�D�|T����˾�x~*�4L$i�>��w�O��x[��nF���'�5��ۼ�~����p��Z@�ʙ�A<V��R�����k�᠟� Pzm���@@��N�D�`�#ͬ��D9����������y�-�E�_,Kq&�RLE�����%�����xN>w#���S����M4)9�Gumr��/ Ul�S�A�	�mBۆ��Bຮ"�EJ�"M�0t��yK��������,E��z��f_g L��˝�����	�^����P��x3������5sb!y��P*� ;�$�X�2zOU3E�Oj���ZkM�-�:�#�l'Kq����j��`x
z�
��iݎ��lH��4H����)��1�Qx���V���U���������U��W3_!�����j��'����{_�p^� f ʬ�ł����&��0����cU�Q�!�i��Mu�	�E}ՐM�
;��>1�Sd�H	=g�`�F�32�@��oKܬ������d���̿��p�ޝf|L_ZI3ϴ�a>S�}�����$IS�|�-T��2O�J#�{��抂d�A��� D���o�nQ�j��?�v���/�:(rB%�H�����
��\�c>uԲc/�eh��AL�u�:�	��`��̂��B�{|�,��[ت6�&D����(�1L�H��w��}�m��}H��Zk��u��$j6q.��V�����X��C{*A��s��b'�`m�iٺ�"��
=�I����p�q�M�m��{x^@en��h��SiM�?�Ɓ<ɥC ���Qa�T��Jɂݧ��R�A���N4�o�-�#{&� �_Ҋ��IDc[R|�=j��_�0s��'$�O�\�qV�,Xuu`�5��7ӱ2�Q �� d�MϏ�7�+�R�%�^P-�,�����	��HR|��L�O��F�%��;���	_���]=���ݾ��K��ϰr]S�ò��_~Z�V\�'����$�y~]�?�� m����ORA�o��v t�@���
c.Qp��`|@���_��j���Ri�Y�����*�4�#G�B��E��=Ý�C�'��̱�QB6�N�m�N���Х[�q>|Ա'�4m�����h�ϴ�^�?X��1�k��-��b���}h���,fB�3�)��N�LD�y������?5����Ѳ�\"�](3��i�;��!�៉Z�"JE�>�ɫN\�����Ax3%!Q�/�jl�`3L`%Ě����O�a�{Z��	�s�9�W2�,?��&�����ÍM�����ȡa�O�J���R�i�6J`��)�ȶ]:8�0��I�{_���ȧ�+7c�@+KI��q=z��z�)�-:�W��iާO���-��]����2Sa���Z?ψ֍E��K�
p֙3���t��4�7��ի�i�/Gb���.�D�"]t��9< ��y���bdl) �?��O�� ����R$�W?�A�=.��t�h����L�DL��=�?������&{�.��H�gU�9����m�HhG��Pe���Z���Y'G73�Tn�Iаy� ��MO��A&�o(0��2 �G��[XX�� o�%+^���ܙA����-��P[��zt�W�K���M
?�>:�eAmڝ5�Pe�t
�eV��0V�晳����P�
ˈW
ǈ��Q|A�����9p4����s��꺶#Z^�y{N�`F���m� Z�M'7��B������ �:���9��}a-,����?N�A6A�y>�jE�Y��)L�B06I�ԇFZe:��)�2�+���� ��!���Ekp?�9ĩ:��k�W[[�h���Zh�ô�lK�t�f���j*0lwb�rAh�wQa���O�7���L�c-�e���8���}�R0�l�[�.)j.)�|4���X�#\��C0��D�:�'Q�0Q�k��v?a�ǎ�u���� �z����3�'t�.�ݾq�s ��0y�*2���7�2��Pn��۽Q�����~h2�ɵ�E��<� �o�9RlXW�k?�"*儙�+[�&��P�x�iH.P(Jɴ�OFقhP����>h��۝�I3^`V0b0�O�Sx�s}�3�Jgѥ��{���f����B��͵��K&o�k�ƆE�1
ɼuC��Ҁ6PJE?6XF���XqӒ)�!�ޤ0W�g�9�Qg6u��z�d�`��[����!H���]<��O��P"��wKc^|��a�g�o��ٯ0��K�[�����MW�|����\�rUT�&��ƻ���J-u
P1��B1�@/0\60�e�|XO���`ܿ0�آ�zet�Q�y�28(���L.�!	E�s�h��3��hΏ}8�X��P"�>'�;Of��j�W�i�ܵ$��Bѳ�ʕk!�]�֮�4��%n�k2�P>��)�����Rd>��鞼{9	�DK������gK�A
��
W�W�>

T2$��n�O��0�3ʖ���J�X�(�5�U�wE�n���#Yd�]p�hvM<�"�|��|�AsMJ�!��A���bΊ�K�K���J�JX��(�F��$_*ty����B-Dj��E�C�sH��Ф���G��@$R��}�K�[�x� �@V5��"�%���9�?V�j�si�w�6����F���,���c�!�a�U���[C��Z,��Y���na2@��$S�|�׈9�=1�3��}��x�O���|�|�͑��y)r !�@H�֓~��� d�0d���R�V�nE���.?�Ʌ5�E#���%tԀ:�0��W�p� O����QqE�XX\h�TK�.�>�<��;V �x.�i���0�,����
d�?�8훲��H�aA0M���ȵIy����B�������u�*���E�@P���r�k�' �����Q+>���|��Tj��^<�c��Q���7���>����׊�/�.������䔊߮���_�-H��*�t��������?Pk='��K������g6�]m��3)>}�B+��Q�p��	�DA!MH?��s!�R�~��T�Y`��#6a�i|w���:��c���p�.�2
me�X>w��ƽ���h1g�4*M����X�LfֿLah��P ����������`���²�x�"�(��0���fP�x�Z`�
]���hR�=t�x�1��rSt�®f_mY�10��W��y�_��Z1'3n��Jgz��ܛ�Y	�{�C;��΂K��-��mFX�t���>��7ba��?��q�e���xR(�[	� N��i?��͛��:]�0
�?��q���D�"�-X����8/\8/�t"�4��ߡ407˺���X�����O!X���������Is|<_X�	A�̩x�wK{�ch������p>��>�G��Mk����Tzr��w4�-��_���*4+��X���r$����"C�R�����O�w�{W�g�mh�=���s�,h��pi�8��A�	�ʛk��"�O~�����1(F<Ct�P��}��3�,�@ ��÷�gg\F �/F��3���{�ֳ�%�H?XA�0�����Ӝ� �3�N�����1!3x�Z+�{ky�l,@G%��C.fB��+�����-���Kzs�31�N�(!��~B��C�E�17#J�p��c��;5,ؿ֣  d�P��.�<���e�F6�uy46�-r�͛�%�����C	!&n$��4SC
��0.]3�a�f`�n��- �47w7!����ꀓXb�<
-4�	���q.;�W<Ӵ�c�e�Vd
^�BA[�~F��X2�ønk�)�pt�w!c]�=Y���j�Z���w	�{���`�^����*�m�c���E���V�MGX���:�3J�m #�y'T��;l�Z���4���*��V���5�E��Kj���y������ϛ��O��F�I�[�3���m#%�u�k/���\Gq�(��R��em�X�2���t�R�X  �tº&m�ެEi�s{ޜ��/��r-R�
<��=��g�s�m�<r���*(��fS��0�#B��f���O���-f�Mo&�e�;&x���}ԃ�jˁ˛�r�w�W2��g��M�;s��)3�8��j�R����aM=��Z!=�����=w��I��z�a[ID���5P�,�lQ�{�O�#h"�`EM���s����&�G��-Z�El���A_��@H��x�Q��,\_
{���'d�u1J����n�)���$�ʕ�\�y]�@��+�^P�����rOPkׁbs�B ���d^�����b��|��c���t��e�uC��| 'ǘ"w��X�܉ϸ;Ž��BX<z�)����X<N��R���XE�\SAH����8�cF��G�3�8�?)��
�B�Z�ųMkݧe�<q.� ��~�������s�'9����蹬Ym�8�*�!#����Y~�vf7���!�Q�!-o�X��YK�$�،��'�|JѾ�I�:�@@�˲
�4@o�t!�J�'�A��,A ����q����:�GdV{���6����^�@&�O�L���� �����ӎ;h`�1?��j!X�܌�L�/4jK���B����e�\��3�u��A+~63rkֵ@x�_�h�|oh4BG��Ճ��F�{�v�pXsw~�m'Sr���=���|\X�ƨZ4!���2�0]���|-���ΛQ	-��3J1 �į|B��E�:DK��f����o��@�u�6,ˌ����+��k��%4� a��t�{`^ӕ�d��@�%!�g�3-Љ�E@N ���V��iCͱ'�'�\�N�:
2S�M�I�F�v�Z|�a���#*����+,JMq���W乞Ӆ1r]���{\��,:EM�5xEAK頋�mA��[��Ψ���B��/� �uA�(QكP	-�*!%�q�/���5�y�Nt��7Q&�3����æ�e=�x��%-AH�K|�'O����̛u���ȅM�ƅ����Z]�K�4j#��gSu��^�՞�E��&��O�9�d"��݂���9v~:4��v�[&L�?�É
a,5lҷ�W��Q���"�{��(�92Mb̪&����k�`=��r�RC53�?l�p'�to�f��[Ǝ���_ӟ+n�F����T2�\j��׶9�8��`�eM(�E�Ƣc VO��������P��XD����@�:ϝ=ל9u6r�B��4��� O�C��/�Ej�aWC�7n\�>�-2$��ńx�0@�K6F����
)ٓ�Q�Y3,hk��dX�z��{S�O'��ƀ�¨Nb���3���h�r\_�����N���~y�T�r���H�+]�)���3/�������ϕ�sB%�&p�P��_��]�tʗ	3m6��4)�\��Fʖ�hb��4�%�"�ȨTX�z[&Z����nc�5��}��ԩ�\�鼎�@�N "�_k��(5̍]m�*���o��!�"�J�AcvQX������λ����-DY�z�W����
y.>â�E�&���a��f�������k�KYQ�Q���k����?�K�M�F����Ʃ���j+�/L���" �$�����0��$��˶�9j7y8�A��~�g�}&��k�ﱣ)B���y��*��o���}�ӏ�2/ˇe{%4���L��2U1-+���sɀ�͒�XX���1/�H���$ĩ��"����ʒ�c����g��L��(�f���9#C������F��1���e�S��I&K�5��!��o]��R��~T�*K�oѰ�k��)��M#V<�����P�NZb�,k�wu��T_��޴b�^��t�����j��U������g�J9v�T�ܗ�7Ͻ�@�e�XR!>����Г���\E`�O^�%:�T�@X��"A�(�$x#sɳsMp7f��Uk�~y�G?� Q��`���H���>�;����G�d�#��Yk�GXB������GA��7 @�8���B.�#
���}��Pc��)����x0ܶ�j��H2��R}b�5�������3��9�&	S�0	6���2�sh;r�^��wq~~����Y�O!�%�眤?Ɍ6��*D�X��:VL�~�_����{
�_T�*�u�G�������S��-����V4���o��V�g��p�1�����R����iCh>���f@c��a�f,�C̋�/��cї/�چY�+��`)�����sj����nC�ʺ�R����%��(a���f]x1O��W�蒆��J��{�B���BZ�:�k�8�v�B�V<���]�|��B�q  �vgl�C������zC�8�G�G����C�4!�2ki�we���A�E��� �î�`��8R�bI����k�4�@a��a%<b��>C��6v�z:���Jt�e൅>��Vp���R]�<�"�"�` �b�4�k�9�<FD��i5B%�ιw��o��qX�Y�j���D ~�+/E/F�)N�2-ǳ��-��ߙ�|N'h�߆�b�e3wr,Ur�*�4q���(�]�=\����|�6�������� �e��-	>|b����)�c_�9eͩX��ָ��D1r��
�!V_��>��(Y
T��>���x�?X���p�>��o�;h��Q��$�DRx���̃&}��p,B`U~K�Z�D�! Nk��<,�+���dR&�Z�5�{s��~'�7-��a�.����d^֠��pá}X�w���0ȡ3`��m
��t��}��ב��)���6�)�&�ߏ�%�2(Z��56"������րS����?\a�G�aK,�2W}2��C�#ٺ��
�9?w;)f�D2\���{�3��ȵRx/�z�,��qE	菹��cF�JWmaz��qC�P�ך�?x����~U~��Ei�_�Ӊ�Lm�E`���6���w���V�����p���u��EX;zy�L!ݶ��a�kAg!�tJ�?���B[��a��!��Q���C���+z��z���<���z.��1P��+����﵅���;�y��P?O�i=?�~fC~n�s�p�Z����x�{77��Ҽ�s� $V|�� �Y��3��������O��� �dO>�ԂS�N7/���v���^m�\8�kso�#yygX�駗#�+��8��Q���	w.^�X��ۡ�Ü`T�D��my���Փ�?���Ҽ�x<ϕ�B��7��.�P2��$c���--�w��w��z,;�W+�r_C�XR���sl�Y�q��!~���ܼy;���2��o�n>x�C����'!�1PbFbf�G�lАP�V�pE\�1��q8�=�w��2��qRH� �BS�5��;�����W��ՀF�.���|ף��X��Ы�71F[���I�Mw���|��PDHu�[�"`'&��sB.?y;�I�9�E�z�`��6G�}�[�� ]�i_`�7W�V'1j�}���9�17=��^F��c�� ��,�ڰF#t�	tad����^]"z��sH��OE�p(<yfur�ap����T�a�Ee��!��a1�w�������(
a���� մ��PZ��£�F^l����V7�2I$v��0Ѷ*��L4�����}��E���[�@[����b�������)����]��P0+����BX�kQa��	���J�)���?�nȁ�=mJ~�Y��k�o2��-�z��+��%�+^�g~C�\��)ǹ>������ʃ�)���
���מ�'�̺���h^%����������.!�-���xA��_�9�����nP�������Y� �~�+����\
�Ⱥ���t��d�L�b�i!�6s��aH�p����s�]Ž,���*�S��1`(�1������̍�X$@���>�ѠeJ�=Q�:�Y�J�O�t�6B�#,_s��/�m�4�s�u��e�ϕ�BO��6cG��r��^-��@ڷ�Ь��SZ3,�U�!aT���ǌj�:Ȋ����V�c�A�:�g2&����me�ֱ=v��{���� o!눜p/L���P��6?{�ƕ2�>>׵�����Q�a_�=	B��"�Ш#Ey@��̶6c���T[7��^C�z�/褾 �o�Q�;���Vd_�yΆ=f}l�[�`~A԰�ۖ�;���[_M��3e��jh�.[����*&�?�T�މڟ�DC�q�:��5\0?����9��dث����*K���e�;�˴�M#I�S� ]�p-�2��K�F9���R��.3jWF:hi0P_g�����on��U����?Q�d...�%N�!R*f�15����"�< [�,м�y��U[k|���c0�F2��nkm�FS�P�A�*FE)�p��5���TH�2ZFfXh:4R=J#"F���Ah�3��E�g[�><A���]�Bmꭵo�����}�x �QK�P� �'r���Q-��R��[%���Z{��cj���c��̛8������X����6�^�������6����{���{��|P�|/����׶V:��5b��Ia���Ǳ�F���f\Eڅ��q� �ݗ���Jr���87��3;%�)���@9ii>�	h����3�����g�4��_�+�?��7D�b�8H�g�OK��u��3�/����)�_�
QeU̟g��r
��P;�|5�U���t��A���.�|m��"tQ��QӀ�O�4�g����E�����w�\BB:�/nL�#gpBB�Z�$�s�AJ��{^�������skD��&�>�Bg�J1�WѤ���������1�S�ق��ި�k���|'�dxACДsPM�K�PC��'+a��:���r���I^��,�L8��k��&T4�:����rS$��m��(�>a����Ѧp��vcx�l�ZB�c5A��{�<զ�S�Am��."`�N���M@���6KW� "Zt�q��a���l��2�5vf������5��wv!@ ������SZ�;ڕ�5�n�:�Κ�0ah�i玖P0�"�'j��a ��@W�@S�t���{�Z�2xRMk�`���gY�$|�)�WB�Q��B(4+ҜP �+�;�4����߷9�<�I��h��(���F�a�#�z���L֕M�B^b|L
�����@�f�Bf�5_�g�Z�z�kE��S�m���ߣ�{s\��f�-㬨�B,�-˔eZB~G	�h�7�*,&
��)����M�D�BI���1�kC�R�˴Gb�;�E�4�l���VI	����szD=�.�I�p�׿��H��X��@��35X32�4b��&������(�����������Z�u=Цb�	qI�Z��Gh�����d��f*��xFc_{T���q�o�V�Mӥ?x3�`<��p,�I�����Pk��	��}�{�A&�s�σ�ÿz��)��k.�@3 3RcwF��"�O/e�����#ړ�Q�=�p(���C�	��D�4��(�M26{����o�&�믿���W�����}�q=�<�ACjQ7ꆦ�`F�g3�e�Ϲ���gZ�<����D(���<��(+:��U������,���^�Q�5�឴�ִ�Ⱥ���<�V�MB�'���y������'-������T�H�O!nE��cAX#�K/�
/hۑ�<S�+�u�5���8������j���J��2+��$�}��l�!ք�J b�N�y�~2�5���ٜ���f�^�{����LrJ_;��j³Fm&W[r��X� ���Y�%ړf��+!�>:��zD.�	�}U�{D�bo�Pf���F��5bӖ;��q�i���H����hVp�� 
J*��~W�}<t�f0H���v�����:�p�L"c�B�ft�����gHQ)�V�_ܟ�&��<K���;�?�D��"���Byt��������<�q$ڕ�&�tCQ(}�2Q80R�j\�2yi����Pka��nx��a��A�dJ�h|8�R��zڂC�!�0�O]�B��C��b|�Z��xǏp-C�� ���ϳ����5���朳gA("^���%y1&ӹMƈ��-5�i筓r=���Q�-aK͚��:[t��p�M~ϓ	x���������?j�$�xԞm��o�rG`���J�ٺr��2\�G(H����{���a����4�B��o`��)�����|�+��
ߜ��3�,�3�,��E0�I2C^�rgۦ|q�%���(���zi�&�6��(:���^��0����{B0�%���(p����p)c4  �z�%H:�68�{�9+A0�V�B�
��*�Zi���LV�M(.��4P��A2��AW�ЬcHL[歆D9�{9��4U�t$�7����z�=Gټ�1�Xk̜&~��\��Ac�9t�kh��X�Ո�B�{�(����n���CY�F�c�` �	�cp��(����/��nB�N��~�T&��~ R��m@�z��~��Qo9��+V�F�zܙ��1z���?w���әwX/B�P �����q��I� �/^��oQc��f'�;�0��B�Qmm��%�����ྙ2c� <��dz�|c�3���[�I�Ȩ��+�X�X��nʕ-���)[��	�Q���9���p!%��������&&6΢�tw���6r�>d'�gq��)�GK;�z]Z�1�a�I�T���RRl�{�1v2g2r�+~2f>�{��q�����];��kG�d���C͋��Q+�}�3ܔEy���(��̞���� �K
�YfS ����-CF���t�p�8̶&��<��>ǌ��l& GĚ)�skY���Y�b�<X�o�����A\��X�=�k&�E�,�`fc�(!��3jx�V�L�C·V�[��9	٭��V@x�րHaR\!��(�U?`0�V��9X�^�2�?��R�c�����ߑ���� '2��K�M? �N��=�p��`�q�������G?#Q�F���D�M2D�2��pOˡ��n�1�1��oӒv����b�
�d��	�e*�|��q��oh�A��I���-�\j��Qp�1sMD��{~��*�<��ז�a���ٞ�p�I���.��`���3K}@?�sDj��5��I���ӷ�IM� 4�n�ף���PiZ�����������`︓��>����g����������,��A#��(���(�ƞ��������`�:����Pb����ϼM�X)B��K��:��`����������ˡ�V����-�௭5\������3��kE�7-�~�^)w��FD��g� %�Ք��w�^�R��L3HR�Z+禙ֿ�2y���\�1P���ܻHR�a��@P�|��E �Ҵr��X�k���b�kT�����6̋\��������P޲6�-m�9$�}��n'�&����]�[���c+�Q������E��!�ܐfZ���9S��2�o�3L��H&��Rc����M�sx��<��jor3���K&�T��E�)�(�Tru�=�G0�)��~%��o��?aV6���!	ږ$�ð}���N$�(Q�@]����,��y�'���5h��`��	?�$,_�s�׌�;�H�1w��A8�E������ie���vX�k��V��)
���T֩���\+���{�ր7TJ�_^u�LMǶ`���g�'f�C�?�+ �)J%"_���a���[��?�}4�կ�
��=��r��+�wN��{GϽ.���o�h��r�6����n�FW����Xc&����8hh�r�M�6�� [�N0�����`�r�a��Z��|:8���Ѳ���?�����#hˑ���`,�瀅_� DOՌ$��9K�Ů��hs�����>ǎ�+1Թ:eF�0�_*1���Ƞj�}d&4����l4�3��;�Mw����v�ח��>���~Ѷk�7aìR��2��c�4���?m<��
��t��}6֔�P�W�3��s�S��K�M��06�G@:��Z��-��D��7��8F6�vO�/}���P���]A�)���I�R�dȏ�p*���nǘ>��_������!TY��TSX3fGsj���XW�۟5��{�!1�S�������շ\����Q~�nis�s�I1>H��H�����?oB
@��4s���Y���d�A���Z������;Ǹ�y\�9��|���Ӧ5J�;�/�'�L��o����g�����|�����D����H��	��"P��q�h��W�k����[����wj���ņ�t&�)[b\�I��%�I���)�HV2?t(KH������L����0�>s�s�ě��XH�bf�$$4/,��I��8 d����m����sqZ�+4-*�dx�����]���w޾�� ��c0�4�_�;?�&7eǼ|�ݯT1��Ǻ�{���a����έ��wc�>*R[��W��/B���3��p+��gC[�mZB�O�^\XXl�M,<:J Kaf�ۉ�i���~���aO�og*��o"��0��?�㸆n�ɥ�J�]��ܝ��}��Gt=h�����C�h��h��2���B'���� ��T2Q��O�jA起 �x�h<Ă���Wz��x)���%Z
���7I�e�D/@<k��Eȅ��.�')�C��Y���;$�
}~g��~� |u)<X���?��̙ӥ��z��K?���F
�ɂ$$��ڠ4����d�L��M�Ջ�����l21�C�q���E��^�ܗ�GH$�J�N�>5�ׄC��xYΩ��f���1-�H����c�ɥ�24�N H�=G�X�`�;1�L31^Ϲ���Ȱ�S�7�^�/���G<тd+,.�Wo�����kmq����Z��؝��9�Ok�~��)F����g�����	>3m�b��ZLy�Q�Kmnv߱*7)3R��LZ�J��u���ܾ��v��1(����O�3��7�ٟ���C�N�o��J��Z�^KA�E�oޤI����ٸƖa�5H7���w���W���Ҟ���Uj�̨ӽ�u�>￵[�]�{�Q{mͣ�����X���+ױ������ܐ�B[��Z��°�H����h:~t�k�� ��A��� ��m���f���6߲�ʚ���]\\����J-���h
3�EBK2�&�ql��\A�y#�o^\��5�{4,KN������>���@�Zd��l�яeJ�X����ft�����ሷ�>�$frM{�f�^}bf�핑�z���g��o��%�#���][K���-���O-�ڡ�1���bS�p�0匾~�݄���A!<����9�c���6.8��Z0�����3����20��2����f+��:�&|��'�b�?ya%��[�^����4�P<�0(`T���L�I�*���(�IaF0�;w�vO:%πF�Xo���O�W�W�aT�p���z�y���~"�І�g���FΡ����g��\1,f��ʉl-��a����f/�R+7���tP+F5�A�	W�o����ʒ�V������ä�/�Y�1���Lkm��!	5�	����*,B��)�R���MA�:>�Q3g���-�=)�Sq'�W��Vࡥ��ۿm����-��a%Z�ٚ3�O-�*��8r$Ӏ|_g� �Չ�����]���y����k*`f^8��C�=q8�6��(�@3�:*��[�	�fL�� G%��&�<RM�5[C2�UB�P9Itm�pg�/[C������5l���r��|v�������ݿ�0�h�`��F.0�k���F��\�O5ӭ���*�LP�n�cK�f�Q�T��`A:�.|<Z?��֨C�3Y?�I�;����J� 6��F�
;K0:��9��P*p)�a/���*��{,ߩQ<�����>�!@9���s�O�R�8�	ҹq#�(K*!�5�Eq�h�D0RR>
��>ۯ�/5��t���<�/w�7G�.F��;� �>�~����ӂ�sC�L���NAH��5|��*��(�c|/Bs2}�\�����Z	�!� �o��=t}[s@�(=�'�t�X���� #��4��N��f��j��X��~2�:����i����7t��,阇+�`+Z�y��"=�Ö6!�\�N&� �T�����Nj�	*u䘓BMT�)a�k�L,5|X3C5�:{�&L�����&�v�(kI&��!���M8��~fCI���۬-Cn�A�����W�{	�>c���Z����
X,3�0��15-���a���X��5��4]�t�!��Ҋ�Ӗϱ���-8+�
,�@lI/�&�߈���Ar��U��f�����q��� �B��q�,�j?N2n�����	��'%��8�8����R���B@������vα�!�A��Z1���0�������
moZ����}�|�}�T+8�q�<!Ƈ⭵k����b� "�QAG���w�Cl�T���m��"��G�E�?'���<�z��0�*TX���T���PJ$������Ck(F ��Sgx��!+;�%�f���J��CF8��?Q�P�8���.��=�8�=�����G�G��L!"�~A�m�H`����/��G�F�}pnM��4��D[�l�A��$kuE&'0Ѥz,Ly6w�	�9j��A��ݯa�|ؑ�8������J���31Z݋Ŷ�h�p�#1a�� ���i\>ƛ��x���K�i9aiW3=9����J�[�.��`6��.�#��!�k���k@f�C���'���y�ܙ�n���LTM���?��?5���/E�������tBv���ǱRhAQ+����W[{���)��~g�/�V-����
}�Q�t�0B�I�E�Uɩ��}�!�����lD��a#[zV\�x��;������4��@-ÙL�*�o�t	֝u%�E���@3����RК�%���t��ǹ����,�>x>s
���������N�:�+XF7�]��㤌�P���@<Dn(`?����`gxB)Kx��YGmJ?	�4'q�VwP$0ױVo"71٪Km
� +�F�_@�o'�*[ϠQ:�󚂵hn.?dr0c�_e���`����n�i�l*�C����zY�چ^�ր�,P�Ǘ�`Z�(�(�u���q�D3�P>?�Ҍ�X�m#CX��g��5��By�N*}�ԩq�/~�u��UD��/�<A�a����wD��+�P����?wC|�a�h'd�������U�{YX�Q�{	ҚB��!���4Ҳ�@�AC� �ʝL�2����X�:w�RLB,F���EX�%��W"�13���^r�O����I��W�p-�u'�#Q�L��u�u>i�賡\q}d�$�<H�,�v���!`w-?u�-:O�z�@��ڷ ��%n5
�J��N?H1�doS�����V��3k�<[��M£�Eh��o�EL�O���O��:�Z����#f���	�a4;G$v��&��ź�:� �G8�QY�A�[.}y�V?��Y�i,�+V��q�̓����B��4J�A�H�4P&cÿC�7�)�7(B/�Oe5�	�Z#P���4�k&���\aF��m� ��b��#Ϭ����q��F���9�����bQ[��J��u�0�cL��,��t�U�H��ץ|����(8�[v�z�P���X<�e3��U�Q�9)���Qr|�?'���+������oLB�n@߶޸�-7+aV�~�?k����@��p��[��#�쵘�]�Vo����D��׾�&hCob��+�H��J@�(p�xe����Dڰn�Zb���&�
�j1:'?0�j�B�6���B{��8��TF���(���΢1� �M7�f����L��Prr.�Y'�R�7�U4�{��(�6,E����:��t�ޗ�;��*J��v�~���ڒp-әE�]��6��4�0F�$�W0K�M4g�_-¤`H��
�C�-�/]!
��8�ܜr��Ν;!�t�Τ��ƱZ(F䣊� ���y�x86��a�����[_֏~���|�%Α0��X8���Hz�� �-��b��y���+'��&�������8��8:+�i2]z.Ϙ�0�f�;��2+1�)�
�IH;��;��U�0�HOL$����BN�D��#Ѩ�sQB&�yu^(��Z�;!����E���/����������g5��a��[&���ּ�Y�W��-:Z�ψ�M1��W離st?�p�h��Dpp�R=ӽ��r�d��!���eK�iҝbR�"f ��.o7Li$&x0���9�db��J1��Y�d�_W�q����.�v4@��9��{o���w������=E�~n9��AX?x2H|��(����ؚ������r@2T���@Q�	��5M/Lm��VA	j����M[Iu>,4����O��ΜE
l��孴�A)��
I��_��̱f����g�g�9�X�|d��+9�zظ��{T�ü�/��t���So����}��4�S�+[��s_��S,j���-Q�����J%c�i	O�KB%'�V`�?�j*+�|��8$�9�8}����k:��M%Ej)d�"E�H�_|!�d���{Z`9����]U��W&�ӝ"���sj^�Ϩ\TR���yeR��� ���t?�pQ ��@L������I�Yn�~�P�Qj-4Ly����zoH����P��y�;�c�<@h��Pa�;� 3�6h:����c�PWn҃�����@�H�8���G��ҷ��E��n����"�<:2�c�@�n�f�<{���'��;��q�G3,G�9���`ӱ��!;3dG��X���R����>
��uI���)�%Q����;��6�c�k��C��,�������>6i �j��S���|Y��K���$#�ӧ�����poqٰN���#�k��u����_�T���˿� �A�Cya�l���?�C౶\˱��X0�xT7�f���� R�m��m��}N�Df���_A��C���p~%�2��MI��V�}�<��S�0&��2I\�U'�,�XF���9�8�eDř�%�BC"�
a�(��g�i��f����������h8� g`���)f5(����_��-�>����L�QƄO���7"��S0#W��>rG�q	�4��<�8|fw���?k�5LXOY-(��/��P�+��	�x���?�9sM_��{]��P����/��8��=�u��T[��p�AkM<���"�|O�qx`#*�h��L�'�6Q����L����:чL�0��Ws�[�"t�|��?��
&��R&���S(��׵��O^n���Lיo/���p���Y�Tϵ�;�^�y�/uF�E��lh +z���;M-�W��<xO����:$��C8�|� �5��M𠎯���p6v �@�H:��X����XjMѰF��a��׃z�?\���@m����fR���Au�������T��;�缊���'�ʜ8q2�`.(b�7$t�۩܏=Z���Qކ�mQ2��։�ޯDG�v������r>�d�P���c�5���I��[��,��썚�{�=׵��� �`���u�cv�>��������_�NAxH���#|�AS�!�lCP4�@gH�}k�B0Q����bߘ�-��wJ���y�iY��Qy�?H��`	��\a��6��5vp �r:�猟�u,`X�cxހ�3*4��e�s
GA�6uμhgߝ'���,B��������f���fT\2�,��96k�b�&e:2Ț��jM)�)�_}mm��T�#�݄OmZ��Yx�h�>`s) y^4(���}2%�{����m��M�AjA�Ӝm?&��~�˶�����c���V��q������a�>��S[nQ����V�9E&5�dYi�v;0W�[϶J!T�\e����_�<�E@�0�w�-�`2�!g�K�X��nm���ma%�y�??�B�U[�V�<�����3N�|�`6cI&���V�ǚv���nk]��Ӿ�צ�[j����c�r�
E8a�,M3^���Ňk!E-�14�
���N�)�2�<����k���/˱(Y�D�p=[�!�T���Ϋ��w����e��9�����@�-C[BC��9'�G�o񇛧E�~�� ���o�T,B��H�eI�[�|�Wy���݈f��������/�e^�Z�<ۻԖM� K6��'��N�e���5����Qp�aVkޣ2�کkmM�Ee����w�8�ڹ�^Zd�d�V�MI���,��x����?�$w�}Af��^t�K�R!�p�	;��:}4f��J�e}� 	���w���A!�����]w��F��BЩ�@\�ۮ
ð�@�=��v/冱�<�8���?0B"9&���B����c�}��vD��bE�9����sڪ�L}��:���N�ܦ`mϚ��;�8�#� +)@̗�f�x)����5}�>�7����y8��߬G��Z_�2u*�J��_�u�ǐ�L�=1 V�xfӧ��g�-��{;��c��!^�y��v��i4��Q]�q����-9Q�[�G�ɭ�0ҫ����hι3Dʄ�Aԋg��(}�Q��([b?���քц��x�Hд���Χ��\��=�PS��n�����Bu����1�g�f��	�h�~"�<����t��~Ą>ͼ�}2�d����ۃ��B��=<%�pКC�������k��e�5苽��5C[��l��=�s��(��f�1�c��+ظ@�y�����b}�a��+���W������&Z��ݍ��B��׾�Z���B�_�7�kk��^�v���	�/a���<�{��%^Ĵ.S��tW�J������E�Ro��ȼʲ�y�4��9W������;�%���0�۪5��n�b`�IX����i>�1��H�+g��n��G�'R/�m�8"�I�6e����[���5�x�ﶉ��t|�T��gAJ�*۔tI�5�d�7c�	g�b��)�fp�������.�w�=����f ��m\֟��1��޺9�����jߟ�7��Q�*�]��	���!���PK$J���|���:�s�q�
+oљ@/E��Z��Ο(������aH�V����֌!���f���R��N|V�˾u����h�ؑ�����J1��7'�:-�sD.�YJ��%�!�Ww���O(�P�p���?�Ih;��@��A!�oiy!�aF� �6Z�}v��,��o|K����Ru2J���,e�3]G�X]%a!�:rZ��^l���=���cJ�$���07�1߂�We�^׹_H���	��j-�P��ڮ_���b���
�ꝾE4X*�Є��S��Z��_"��Ebc�+�hgf��(&6�ag;�\_��{�l��ںe�x;9�q�(�F��M(^x_��|WkD�p�iC�*��YrD�#��w���7�vM:}T�j&�����a£?�a��;�N7����Q3���y��V�w����՗���f�t��sw$�����#�
+O�We�;�n����M?4�������1�~&G���f�g����}6����ڷ�>"\A��q��f��-L�%�<����y��Q[��_�jf�ܶkT��5|`
@���c����9��j��o���8B&e��ҍ���\�v�R�w��>!2�I�%��XW42v���+eD���-��;���~���?�S�|;�o�=:{L�K�T���Ѓ�xV�����Х�z�O0-�䟙K��̣��I����P1$\���Ѩ*��$�3��V��a�L��#�%��-��!!(K#�u(A"0�h9��l4�*G�:���Vjaς���f�F�	%��m��Q���t�� �!�MS3����lm6}�U�0��u�~��5k�h����t����Ie&S�J�|X�%j����]R�Q��-$b�G~���~���c��M-d��*��SLNgI��,�Z`����^�gM�����m�mXٴ%��<��E��ac2[?_ݺ�r}��ꋅ�Q���Z1��s��:��s�m(�$��i�[�wV�B�)HK38V���ĺ T�;V ��(�BA�(E���JD��8Ou0�p��&-ѡ�@Q2�	�q�C3̑}���b_�\X�+ɝ8z�w~~x$�
��1��>�Z�:ӝ��G�rwI�5=��u���P��Z��a�$�tɰf�$;�.�]�E�cGtRH1	�B��X[q�<Y4�f�fDJ�=W���{�C��v}f���,,-���dP�[Y�<�r#�J4���{�S����z�R3ܝ���qAEH(
O�vǥ���f0)��f��!�
Ahv��A��e 4
A�(�HD3]�-��K�J�k��ɇ�X�L�I���\��w/�\S����,��k�1�������:.�[C�j���],�\GO°뼹���܊F��S�I^I����emנ��Q�&�E�s\m�.��J�=�UkԊ��?�{G0��`XJ:fq�����o|CI�?��z)�ߡ)����Ns�<��;���c0���2?��S�H$��ݡ�Q�\�9����w�:nU�~1>B���PBa���j��9�I���"ړ�j4o"?��x3��G�Ң%��g�ģ�y�2"-� �7� �Ţ���"�C�7Jm)���A3�::��ж��"�f�̒������3���#���V6̜W�Rj&�u��Ž0LYI�&sͰ)8�RU� ���T
�C3��A4k�)CS��`~�c������nڥ��0�^��gڍm%쾞��(I!����� a������m��b����:�;�u��ׂp@�)�>>?� �Pl�}q{�Y'~�9�v�v*Y\�\��-�Ч��k��Kt*ϗ�|.�l��O�����_���a�n�ct�+~ּ��aD��5�g�c�6/u��sN�g�[�Ь�-ꌊ�U|߽c|{%X/fO�9~]�p��%�L��"AU\�P_޼��>eUŁI�1���s3�J���r!�����a��'k��>��̰��s� D;�Sȁ�B�~�g�Y�nkBB���"�
��eMl�k�1��W�Ȉ�z��W�I�Xr��q�W�����=�+��L�A�#("iv)f(�5��+ZZ��UD��A&(oH{^n�^���됟X�0�S�N��ֺ���-�º����S3�ִe!V[;������g�і�������}!�댲�?���J9��@�����7?��Oc~��$�+��:�����e�j!���.�e
T��.�����QX=|�Yc6Z.�}�hy&Ӄ$@�r�X�0NJ
����	Di������Gp��+!�ʌ	��߼�(_�cP�0�`�f�~�@�L~������y1�
˲��\7Џ�	*�Qp;�S��k߂P���ɻ%ƾ�$�n:��#G�����:8��(0�HG`L�?��hT��,��Fa&{���^���z�!\Ɏd��%�xf�a�x�l5lR�V�;Ǜ�mMZ��c���*�]3�>sʍW����(o����6��q�e]���E�5��R-0�Z�A����|��������(�Q��g�Xɤec�`�0$��s�8(�<��C������=�����	�怗Z�2����3��L�{����{�k���ӘG��Z�L��K+�oõ�;�F�}�w����'���an4�eNϜ>��2��kZ��[�[ ���\ga�,�<J��tQ�;�`�R��D��P�2��|�<�{�n�Wp}�y�4�E ~���n^x�Pء#,A�?ׅu�ik���F#��9z��3�`�E�@����L���m�]F5��g`��AS^���W�(�ݷ $JG���6׺�^y�,�J����b��v(6��bx@o��� i5!N]DL�1�A�e��1<��2~�Q�?�0D9��_��k���&E��,�53?����=u�<���xB\5����z~�к����?\���b�Y��O���͏;� "@ݿ�L�8Cp`ap�X��H�t�<�:8d�+w�P����b �L��ua|X8�-~:�@`� ������ׅ!�g�k:�-:ϋ���"�36����3��+���o��Q/^�����ﶾ9�O�	/��&ֿ��ه)��L(s�F����j�3S�����ޮ���x��?��[���n��!A ��1���N����|��g�/��Ŝ���擟V�	�4�bn�8oz4M�(�m�%y��绯�یq߂PLwS�ϼ��aY
)�P�)�uf�8���0�)jSW��kt^�Cl�0�c�?�L����"���I�}�2����&cB�E�� ���U[���ٕx�q���ґU&V�:f��u��\j�F���[RÆ1�v�=�H�u	�Z z��u��'3�AJa�0�[@��t�<�3,B�Hz�:�IaΫ�D�eoB�a���_J���0;��Zh�4�A��V�l�|�a�ȧ>��a#������������������`<�(�Y�a4,i��\$�{�GuFA�'���$<+��t��b,�@�Z���<�����G	H,X"��)�μ��7����o�x�@':G�2.��8�:��9���O����r�-��|�#�-Eh\�ںƶ �������굡������r曠E�H�E���g�ߴ�	���w0�=��W�^Ms���`�7��gaѰh,8Z5ߡ5B\(g��9�5�.�������ԐWv�V�UUМ��ש�M
�Ax���2���3��] ��]H}�"c+ߖ~��"�(�TTVG�l����#�i;(����0��.E-�3�A��	�����2��e�B��tг�)�b�����_w�t!䜑�~����2/X��\�z-�>+�.��2y�k�+���@rti��'csd�aǦ��(��̆�}�+���a�ĭRq���U`�ݹy���$B����f�s@��܇�eކ�����Y�a��M[��mZpZrm7v�4�ȅ�"-�p�9�9F����Gx_��%5�Y8��(h�Ǐ����~|L���mi����Ex-���:V+4X��	���Q�N�NF���ra��0�A�ZD_a��L-����6���+�:( �BP�3 ��{�Ǚ L�5l��8�	�x��c��qp��=sc-���u��a����B�z�Р��s�=st^>���4gD�3�D�i�<����c�K�y3��ۢ:li�ohh�LQ�����ޥ(2#�Q��������(��������6�ːof6�}l0D[�뚏|'����s�Q�e���'&Ĝ�XB� f��* 	SN��yY�޳����5�?�0�°rD+�� aj���mL6W?�4��~��V�Bǟ]��ӟ��&��~=���|��~pO�=/�睚��|��C
�Zҹ��7�Pt���>�N��>ﯧ�iH�o��#Ƽ��s>vX�35��ŧ�ˇ:==�O������5��as�|[j3����G��Yp����<u& Ω�#1�! x���_��Ȕ����K���),1���lKA���˱o�9ӍR�x�8��g ?�z�uK0I
g��xW
x̭�V	�_��ך���Vk���e�d��3���gϜU����g��
z�0>y�T<M|�=��];~4Sq���4뚓Y��Y$�oݼ�1���2l�TFb���,�G��֡��pƄd�a,Z������}C���r��L��$�C��(���f�L���`�S��C��d��q�� �]\B�#ªth6igB>Uk�����V�[@�QA:Z��{�'��gԛ���}xԁ,@�7Ƥ/���c�[f�X����Z0!�x;��8A��H*�y䓡��̜��G/�����F�X�:(tI��r�J@/	�D �[8�e*=�#��?��j~س�Z|\�{{Qج9_��(*�0�J������B�
�B��@wԅd��_H�K6��j3w�x���駛�b�f�@T��J�L���k3>1h��w�x1�.��n�l���?YH?i�+��=�uT����кw@�(c����@�w�� �pAa�(k��ڬ׮}�|*�q���,�Ϟq("���9O˞RgikMd7��h ��$F��L�Z����"7Pe�O�q�B�\0�XЈ�B���z�e��P�Y�o}�[����>~A�$YS~������TƱ��<p�5�s�gX�Z+��<תPA��1x0��Xdd,��VD��I����y�����̭]G��	�{n�>kz�w��!&�pG�Ac��4��٨g�ƀp�G�$"��j�Ͷ��4[c��43h`�L��5\�Efl���Ќ��AbJ���`�v⚁ٿcK��50���,:���l��!,;�me�9��>���`n��6�A4hJX�=�ؑ�RT�H=b�aq����rSl�� � ���隦`�L�VD����7���Z ִaa�����N�?����e]��m��q<7i�ኘ��L�8�1��?K8�6�aI�6b�Q���n������|l���~��� �S��ݐ�P�C� ��TJJ������T�^�7n��㗿�e� `xa��b?1o�$��B�0��֦��c�b+R�I��+T�2�0����¨�Y�A�
�<-�8�?�A�L�f3��3E-�u����׹��sK�/x~G�_�؝�J43� ������;�Y�:���Я�0t��G;�/N*�d����wW�XaB2D{>4)B��*�MvU���dZ �h4� ���;H2g�����!�*e���A��f����:�6;�/���_AF�>�O[C��3c3��Lo���9���8ΐ�\���d f|��k��EC��5ׂ��Q�7��<&F9�"x�Lc�A%��[�A�N�)psK"�U�%� ��4��'uL^P�v@V%_ʾe3�����S7��"��uȒY|)0,-VX��������L%��F0A��{Y�@8^n��gk85�.�=H;���.��QM<��-��:?�[�Z$V1���݄`�[�����8�eC�H�Ih/ �@]�}���"qqG�2V����Z֡N0��(�|!8��_� N��BlTj!�i�2.~�緸�sJspb�By����K�(�%]�xsUV�s���6����Μf�s�����a>d��s��pꎟ����\î�r],B�q�(#X�{���_N��L���t0��	L�.�W�)��$�C�].��&P�8�.���Z�A�n_\o��Pc��ޫ���5���A�f�bqj������O��Onh���A2�γ3��SK�E�������8�9�
���Jg���o�S��
�!��,��y��l���gj�I��AC�uXޚO�Qҁ"�0��yq�|�����!@B���d�A7��06�!��2=��Ձ�Ah�޹r0-G4��:Rz��:p�Y'� #8+��#&)�s�����1����L�A�׽�_�d��:|��IX�)��EZR"~�����7ߌ���SOl���o��A>�;C�p��a�vъ����Z(ڲ��`%�s�0�s�
,��� ��o������ל��B�h������@���ߖg�HJh��:�e�"�"�?��^8�y��w�.��.�SL8�96���>V4���1ƾ8��E�V�&�o1�Q�$[f@�DK9B(�e��%Ϊ���[�u<�f!h�U R�p>; � ��gհL|aU�j��mO���	֖���q��#�j±�cF�w��}��5`?2��}�yJ�~��A�\���'��Џ�r����_D�	1.a�0D��{CS��K	�g.s����2���vzt�i���?�b�*���`B_����aZ�C�U�J�V�>��?w&�9�²��ʗ%8z^k���Vk��̕c8��`�"1�I�dZXf�~N3�6��gl:\[��sS� L�s&�Pl-k!���|!�������P�����%0��?�q�����F�
9�����Z#���c��n�'��������a�®^��)�W��0��}橨�5����{`I�&p?���EV!��2�|�q�BCi|2����:[�wU�*�[q7�ưt}9��+u���Z��n����)�Fu��.�%s]���2��1	r�g�-2J��b'ܓ�yr-�
s(���hOf#���a�p�m��O������e�pЁ�)o3C���S�o�� %�8|�_y����XK��M�����7gΝ\���ʗ �p��>e��}/ߣ��v��?|��� �z��B-�~}�ߦ����������=�I�����` �b���P�.]�$�LN���aUJ(���2��Bek���"���>t\�m���f�?�-A�7hF_?��W��YM����j���^&�-+^���yii��D�#�|�͏~�����E��G�%&o�����|�u������ˈ���D�HPM�5���e��
�i����z����*�����5H�|���d�a��cL�2�1m�s+I���p�$㳏E��y	c2�E*�����i�9� 쯡-Q߃���k,K:���5 2�7�XW�'����t����[�L��Lׇm"��o����c�Ô�?f^hW��*��lq@���w2x
~��K ����_�b��"ay痙T�l�[���>k��5�[�4�Ղ��-D��C+��B������a�Ƥ�!���N��ĩ�b��n�R�J�Wl���bƺ�c������� �����t���fD��a�H(Dׁ�&�Hh���g��۷o��ų�ȸ�#�|"�2J��9��y�0:��2��wZ
�����SUD֨#	�T�st*�s����Fm9��򝭝̧�v��/������ݯE	O������C皏������5?��?4?�я#H���y�N�%���P\�4ʟ�"�C����!�ф�!�o*e�:e�k�e+Ж�y��'E�|��?)e� y��q�o�
�04�
%�H�xxFh^��u(�k�sBl�yÚ
Zb!l�v8�7���p��1�Kd�Z�;`��4�/�_� Ԃ��G`���599-P��6!�*�F#�C����g�NTjӸ5�	���)�s/�\�`���Y��X�i%�+;Bu7���3�����OmM�eQ[�w��ʺ��f��=�Gt(��$�>!�(�kZ'��_��^Tu|��G��|�YǠ�+�D�be�Z��`L���nS���1��g�ePb�WeAX[`)(�ve�uK@�ψy�_���)<| ��+3M����SO� �&d��5�_��9ʙs�I�{�^�O�!�Y+�I�)p2��=��5�D�@�~p��S���O��A���#�~ȗe���u� %��_6?��h^{����06���m���@�'���D�Ya+��L���=&AŸ
�V2c(p!�hn֙7���k!hK3��.�o�z�X�?����JI~\A0����b�~tGxu��ȅ�A�x��b�	�ɇl]����ފ�*:.��:��e�b!N�ApB;��.���c��<�ϡ9�s,���ޘ�_l��&mS��|Y���������CIz�m\T\uv�9<�rc3�yZ��7&T�XZbt�*�D�EE��=Ӣ2�T��X�|B�Ou��VLIX��N�C��bi���RD@��CW�!��C��Z�7������ڭ��>�l��ڟ�e�m���0@ D�}M5�|�(�e&�f��ec��z�y����ׯ_Sq��(�=-f���������f�ȍ(76O�]��f��R�v?����Y�m+x7	�0-�zL�}�V��D?�1��%\&j�H������XY���O��t3��^LGU��e!�y[1����|u�P!�Ӳr�1���C#0,|�K`5��>r'��wJ�;�9���`Aؒ#�cZI厢�:s_η�"��֑��ٸ*�,-9�q��Wӗ�i�sh:�X[\��{��������I�����aX�0c;�ϖ �3W<s�2���y��
�O���*<@��P&�MQ�}���X�q���
|�t3@�`8�� g�KM��>cR$����ۄ�#(��nw\ρb2K�\Za�I! ��ʷR�F���a3�H��\�l��it^���1�i9*��=��#�+�WrAWe���������w!��i�	V��:a�Rr�� ̰��%Tp9C/c���z!#���Ȥ�hh��P��O������Z�)D0�ʉtFB��*Q9���
j�Y�2����k��|��0����k��w����ֱ��3#���Ԏ �m���Ϯl���_�:B�f����J��t��FD���ީ�D��8R,|8�%���Q�lƍ��2y�s�&���a�p�U��$�x�c1#�<��0���z�XA�<��z��1���9Y�>������d2�B�ACD����h�$��l��"�s�s~G��z�����˖�#��U2�U��r����&��fA_G}^��A2��B���[�a�DٶR��{�Νϵ�>���<A,[$.�m���۩&܇��\'�[ى�/E�� y� ���G�V k��Y����RU���%��\#�ł�ևuG�MJ F�������<},�4�QI��>�aԉ���sF�s᲏<�j;��k�b�g|-�xK�=q|�枟�Y�'[���q�>���ͅ��~,CmX��'��<���s
坚��fKL�2;�h�ų�����Q�*b�QN)�"'�eY�3�"�"��l�(Ueò
^��xp~����W�F�����ڃT�MV�Y}F�kʹp�NmA�y�1@<J&J�&��.��ף2B�7��M0�c��O�FU�*�Vmc�"�_�<�ٳ�e8��[��4Z�*^�	{"�����/#�����#��sN�����Q�]4�.��
1���/�j+P��
���βL8bPx�4my��B2Q9&��9����nݺ�|���$�*zA���ޝ��͛����}ʵ���Bs�~���,&�(N�F8�����m��@�2�"K�Mk!���sz�R�/.f���9/;^�'s�p���e�՜x�W6By@ɓ��W�A�'������W�n>��������j����=�+HE�|�ܴR���A�N�@�L�ɼ;+�N���Fʋ`܀0���~�J����/�eѦ��c�9����m�w.�h����3��B��R���X���AS��ǵ�Ch��
�8u�1[b��}ʵuli�n��Ej��y�~���M�߲�Y����>�|i�Z�U-t�s	�>5X&������bD��afJ��R=�,��6�Mބ���j�*'�f¢�����`�&.=��g�@E��)�|����%�EDd�â	�4J�����wP�y�,��yfd�WQ�R[�xcX�a����`@ԂD�R�����H�As?*���w���f�<w�`|�n�;rCh����פ�&/��H�e%�O���d��� �U`��^�X�}k������ڲ���1�+�g�j�!�=Xq���;�)%���kj=�����@���*@��/�k�o4o)7����@]��3?��s?�>���B#�st�U,)���?ψ^m� H?��rVfq�z���'4�e|p���$|��O�+��_��eꐔ�+�`$��s�W�b�W#�:�� �ʾcN,����c�4��x�F�=Z]ž�LZVQ��k>
TB�����#B��3E�p��W^y%:H�P>A���?9���%�ˠut�(�)�ӆ��<���)��a��F�A�Q�8�1��5���"�~g" ��0���X+�|�5P�ce-x~�u|������/����X"���B��VX^U`4�z�	�fE� ���٣�EY�k�����QM��ŀń�$'���eQ��~~[��6Ф,
O�W��1E#M�
W���Uk(����Po�zS�g�	uP�����iFXlL�c��<��~f�>���-or����Q�� 6-���W^��SO=Dt���]��즤��U��˂����,�%i^&�O�>���� ��( �	egT���]�QJ��@z���&`w{o����i����ߛtL;�LC�V��w����sWi��J̅^�cc7�aa)��1"�l06`RF��)���>�h�Q��H�L;���7c`��İЛ�(㵵��gW�\C����뤐�~�C�o�H�r��.ê�۝�=63V���3or��(J�uX;����K`	~4�4����:r�aU��{2>#I}2�S��k�](�q��z���ֱ6��r^��1�����*O�P�$���i�Ӟ�pb����VC��k���X�~�5[�.�9<�!N֋�yN��+d�Z�X���>7�L@���sxn'ߛ�=����ׄ.Dj�޷5�zܗ�P� %|_a��<9܀��h��+�Ҁ���|�����;*Gqm,E�F+	�M�J�m��4)�R��qiZ�}ic��~g��~�Zs��g����'/<�\x�BTI��$3&�("
&\�ö�`i��~�ѕ��Y���~X{}=o:[�|�|e� M�J9!��h�Y��jX�������A]��r�򉗛�\�φ0�91
À�7B���`���>E{wjF���A_���AYw���Q��Ip��t��e.kE�L��)�O5|j�N�e����n+�6�#`D��2�0���}��'すY [3�ٙ�2.[��{����HS��#P�����P��Gr����T���-X���8���矋�t�Cg��˛�ʇc:CL8��$�����g�^�mm��=�� ��z�њVIѱ��c_��J�{i��N�	���%	+�%h>X�1��$���bBH=����w��C�I�`m��B���P&7�eoE`�c����A=���y�]���B�{a��?�.Y�`A�{0V�¢��P�]2϶����O�����s��#F�[��Ms�uopofk	<�Q�\�l1EK�8��ֆf&\p��L"��U�T�ب͌�ƑC��5X���IK<5ݜ;#��fs����51���o4w�4ssͳO=�\8w!�خ�r²���Y�6��R�!�����"Ga�;c�QC�5l��ެ���,�rX�Ǖ�	�q�J�{�\�7'��~��P(Ä��&	��T�;���ӯ)�7�����6;8�fX3L�ф~?s�r�nB�����!�֩M�g5�eJ���̐j#�rk����\�0Ϟ�{w1�-4��9�!��h��4����������,�����5J@w�h�$fL�`Z`}`|���cT�1�c,�-)��ַ��V.(��>�:I���k�}���=�vb���ҥOS�?�7Vϋ˃E|B��Z����uu���&ڤ�� �icJ�</�����?��x6�=ٿ�v�d�gu>@� �@���JK�ï�2����{��ӝR���2>�_6���J2A��+9:�u� ����V�ܟо=�.��4�sp����4��:�^�>k��A�#H����z�9�M]CD޸!�I��A�u"63\��S=�poiw��� T	��7/ZUO��-�ʂWcc˪�#b����͙���n��M��+ך+��6�}��(>�y�����l��b��J-�kl���������Zê�k.Ѹ�`C���"��Q�(�$U����b$�2��l6«��/�\+0�|r�Ӱ�ܾs;�6#�s�DyQ�e0�`^X�-��lՖ�Û�w�aB��~�`��a���E[�hu*a]�� d���d/YA#kJ��d��F}_,%�I��0G[V���.3ͼ���܋%���0>�?�f��!=�V
�4�y��r/+ �˂�{c��B�0w,�����Q��js刐6��Fݮ��xR[u��P~��'4dG���T;a\�ʶRx&[�FB�c�w��8�tmu&P�F�ޥ�ϒ���|����ךo��!�8��a��o�����?�<��~U�|_Q�X�@,0,�;R��e����lm�71{|6 Rs�:q���q��	�H�����pj�U,17̅�7�.�K@_�-���4�K+����G���2��q9��}'�����A�5�yAd�Z�w��/�V͘T�X���$sp�L�iy�%X�`�i"�M�,�U5�]ݔ5��ה��ghA���m-�F3ɓ�J&�M4O�>ќ��ĩc�;o��\��Y,����5Ǐ�Qh�����ƺ���/+�C�}f�v|CL9B&��u�&4[΅����U8�s�}���/���@����%AAh�l��0L��W����ژ�F3M��r�ΖW�(�YoV>�h�����ߡ�ֿ7��d���eBϙPZF9�0 �鶼�hBs�F�RI� ,�}�}SXe�~>`��ӧOŵ�aN��E�z6k��Sr�"�^�$Bk��}�h�/�� )�)d����������7>/��P���'y��:#��~+�����|｛��e��:a/��gwdj�:���V���sj�s,��%�of&�[=�$�~�����֨��VPK�V��h��ͯ#ʟ=���%̏���ʹ���?�Q���׾���_��ݼ�ʫ�sRd�A����>���'��Y�#��=�]A��Ȋ�)�,���*E ���(���ϲbX3֕��(%	Q&/�w+�b�xN�n���-P�%H�0�c��:��2��'k��=�����%�PX�T���p	I����Q�k���<.9 G��#�ؐ���2o�Q2M'j��e�-�꡷��B�$�S��ͦ�=6���J�[���ڭ�>���MN���O����������e1p1ASލ�&O�(roUT�9�3�HЯ,¾�p�Ɱ����o5}�V Ᶎ�j��a�Æ BA��t�Umb*�G��]�Ԇ��.VyL�ү���S�&6Ձ�Fs��K͇�M}~5����&dH>q�ds�	���8��j�����o�׺ �ڿ���Z��&8�JٻU굺�����l��dN*}l�T��=�Y������m[�x)R�9�%RFxd�a�=����Bp6�u��}UD@f�G���"�ׅS��E��B�6ɔafD��TS}�Q^Q'z��r�uz�-C�E��Ĳ��q���)�
����:������J9s0�:󑨵���\����
w\�|E��G��n�2��𛇅*]���| Px��Հ��Q�Y6���W��tl�0G�fb��Vg_��a�V��f87,��D	 =#��ls�"`%�Af�*��%�~RJ�UY�|�Q�����	���}���_�5����yA�/��X<�aYk?\�⤥�Ck�˓�W�-�5�o���������K��a�5:���� �Ϯ�3@f:�5���`"������&^�!n'�¾`��f�zӽX{����Sv0:ѣ~��^U:c��w!׼/A� 4 ���<���zN�Ϥ���ǐ�_�O�"��?dr�x(佴��@�*�Rã��#M-�9R�|PuaUZ̼[6�Y��tlZ��3�b6���?i��_�އ�	���<y����)�]�l��H�ǆ� �Q3���v���u�c��1ʂ��aA8�,
�����_)�bl���U�N��[br@����~�ig�(��\~]�q��z)�ν�wp�7��37T��L�L4��0�T��ك��]%��v��w���w����3T��`�L�H��o������ R�0��2E #?��͌��[�M���@�qY`�S����"�OP���W6rĨ}�Q
L��>j��8��}�\mX�B&ǜ���b���V��A������!^��`�|ϱ��U��9�J9#:QL�f��Ӿ�L���fĶ����9�M9�@�:���V�.~@[����_h^��Wd	~�y��g����K���������%ݘ�o��7�BP($
���^���I����G2O���y���o[��'��њ������^(ż"'0"�Y�6IeNѥQa*+�$����o��Xw'J^�����7�
�Z�Qt�k�g<��6|�D�~�>��."��MJDƙ�"3	�v�7�q��5�'���(X���s��/��|2kE��T���*���,����y��V4,%���T��ӏ����,���ܭ�X�N̒,���(�]���2v0	��Q|����K88��ܝs{� x'Q�:/�� #�>*b �\�OC&��ِD��5��⎓k$f8#���ǟhf�/bSMͪ�NI�`���#ɾl��n!"Gۍ����y��u!f�<Y��z��	C3�Niپ�5�ﴊ-d�:B;��Rk�Oa ���:A@P�DA�IF�t�<B�^7��A់��uK�Q�Y��ב#�����Z�0�H�%?�9�`T�	{e<L˚>�2�H�B�h6|P$S�ݫ���	U7J�9��0�?������ȅ�)�pV�ଌ�aCt�O~�V@ 7>��SB?�>��6�Ώ��ܼ�KPV��w��~wP��Q8���6a9�����&ׅ x�+�NZ��Bh�K�|�+/�0���sf.f��_�|���O��y$�3��CP+? �m.v�89���D�j�	J��f5/�����\�kk� 𰈅{���"��NQ���3Ј5�s�i��ᝓZs*%����D������o�OEIs��}ڦu���S�1(/�a��0[���dʋ�`sUk��[�D�jpm���ډ���\��Fege�Ɛ�Xk�)���Z�\�$��I�v3ƛg�M={A]�!�<U/�!�~V��������S/.1�U	�AcG7�<N�y���e��ߌ��Q��c�w���h'����;!$�BW-1� ���wi��V В �ȵ�z<J��q_G#����n+���?h��~�M��|�O��ϓO���)�:��r-�U��3��&��R�J�a>#�N�� uo��\9@�7��$ե��&cå0��̊'���q�1�B��ek7x'���H �!�����I:¦	?Ͳb�>�����d`L��J�����`�#9����v�έ@N
�l�`�cb��d)/�ƢR���8`�胡Ol'8S�阂��G�O�er��.Bw)|����w4��
��"��4��-1g���B�'��^�3�>����T`��	�'�T�O�πO���W_}5��Xx��l9;��j%���vm����r�貼�����e>$5}�<3�I��/����c���O
��U��q�(�-���kWC�c� �":T(O���('�h�l(�c��!Ĵ�?!`����BV�Q.�FwW�@k1�:>
¤$���{C脒%h�H~Y� q.fA~���Wk/>/�,�̮rg�:ax��+%��!��΂󩸔
WE�?즾���64r?����Q�l�����ʔY��lVqI˯Ȕ�̃5�	m߅R!6��!���/a&A8>���sǛsO�
�	a�G��"�^�&�#���gxA2˧~�ͼ4��W�5�^S��^�����ia�W>��|�ns���� ;sB�%�h��U������,�7B������G%Ӣ5��{��}�{�0��a ��CDS�#+����a�l�hh$<����_Qp�yE��D���kQ�����%�^�9X�L a�fDk_��<#?�W��ES�-O2��fҷ�����I׶Rd��cli����}��y��ڵ[��c�g񦽗 tpA
+C��B%N��P��s��K�z	,�}	��x�s�\V)i�Rg��p�?��$���a�0����ҧ���|�]���/Z}�������L���f%*�,	FVc.\y�B�;��λ�M8��e�7�E������?.�N��
�	�G�X���ַ�)��Bܓ�r��Mȡo�p:"�gNKJ�#�OLҴiZ���7�s9��o����sTѳ��D�J6��Uҹ��3!|lYF��ޮc���a��n����~�E����qsT�R�jP\0�ml�E�uG�$;�����F�>C�q\�ů��n'�����JB���O<_�ffW߻�Z��O���\lh��S�/O�ϻ/AX� ���
[�L�5��p��r��
2�K�hR#ː�����M�MD:{T��3�s������Rs��ÔN#������S� �s��1�|~�Fs��Ϛ�ڬ'��i����E�o4o��fs��'Q������&9�U�t�/X���Ӵe��4@W8���ª�|�����,���t%��Lc�\���Ki:`R�P�`D�⣹%���>T���B���������ꑒ*�y����%A4�.|J��;�nʼ-J;��h˔<P6㴿*��Aߘ��pƇ暚�N��I�u�
ƨ��t\�2֚���h�rsN =8ξ�N(�>s�5z�f��������/�1�`�R�v(������0&��I��-KH���K�!�/D���M�a��:�UT!o"a����|��LW$���e)�UX���r{#�LUM�	��wIڷ�3�fQ�&\(�9��b�ޔ2w}M�����N��w�j��}����A)nJ�K�V`��\ϩ̍�_�1��mD�F�;5.�S�k"�2P�TJPX7�" k˸�Dp�<zJ��Y�AWR��%P��Q:ye��zC  ��.l@ma����0�
�W0���U~&&UoxV��|Q�@{��x��$NF�t�3Q�&:��X�p�c��y�x��/�Z��>!y��t�#[[eAsZM�^�/2 !�����)����|1[��q��תD�(3����-²��4 �!Q<�Q��w���\5S��4
�Q���q�͂M(��`�����exg�f� V�%�赇oC�?��ܛڨk�:]V����x�����Qj��J���L�ڂZ�% M���,Hi�����#'h;D�`,	�ȫ�	\<�zjK�n�&���d��^ޅ����Zc�g^ցhf+ˊ�_Mׅ��lh��}Y��-m�_����~���2��.j�X��?x���/^S���a����'H�EPV&��	I����vI�!1jش'��a�.�]�eH�,h^̀��O��W�*�f�8�|����|ݷ
kn����4Ο�~-��]�-��?�I�n-���BΖ&�K
���r����dP�fT�I_���a&��Ƶބ�3�0@���3��Dor��=�iX���`Z�𸇫� �#���Cb���oF����FP�L�"��)����1EN���5�=|���`����%��8"F�Y��c�!�`�T��,���a�]/^���K�K�(�&���j-a����K��'�������!�B/�X�[��ɘ�{�c��cٝP (�-�C9��p�4��O|��\C�	�9�9[Ҏ�e�8-��>�Z�%`�q�B?��9�ČּE.�,����>�S���q�ծ��������3�����&9.|�K�?��́3�	t,l.���Dq����<�!R[ֆ�@.��e��v�}[�̪� $�g�Z��r0��>�0�Y9�&'��z옢ێ�W���%/�N3��@���IBN�ss3
���Įnͩ.��77�}禺G߹�l,�� dEw��5o���؀82)X`L!ñ�%O�g�$�om"r�z���Zu&/�ï��>L�y��c���涵����荀H�{���7���{7�� >��>W',�gdY��f�/��Ba��]�TЅ��;sb��H����bn0 �Ӯ���Ф����3Bj���S,a[>�&��,�[���a�ݮ>B0������7M
*��E��?^�}�\ ��J`�P[���}�35*#�,pc��]vƁ�B���B y�2��D���ݸ��\�{ eF>h�'��,W21<�XL�8�����E��)��[��)X��qŸO�f~���z��M�A>YM�@��JB��N @��q~D�*��y�������� (W*%2��)9�j,�)B(>�ܳ!$<_<?�e�Wo��%(�=E�j�f$*����S�K!�SJ� ���g�A���'�Y�� ���D� ����!����/���ؗ(�\a��1>K�=�WT
��jv�`}�	^�8)����y��|"�QZ���9��h���V,��J ь����w��a�;	�TE��+s혐P|cSf�Z��F W�K-h�:�D#����GFbRx�U�A�`��AP�	G�@���т�hc� ��/bF&�������\l�9E2L��Ui�`ߛ��I�YV%���xry���C�|�rs�������g�F/DZDݸv����OB�9{�L��I�;��sh��6�'p�!�ɫr�E�q��Q8��lc�V0���玟��#"t^�M96"���s���U����5利P��+�����`ӰY��$߯~�e1���P�Ts���ֽ#��	8�$~
j$��R����������A�l4�r��Ƥ�r� �F�	��#X��j�AP�]��;
���I�}x~tKsP�a�є�tB�`���can���L?�+"� 	o�Q�*�M%E�kXk�������3����X N]�3�a���I���/X�@�Z?�0�̑��s�rPx��dQ֫+C�auHh��Ǹ��\0s[F]Ԃ���H��h�����a��
� �V��ua��"cB�u�_��D�4�JA`�O<ﳲNS�E ������/�{�L���$E+�b��.R�'|�,
���$�!�/��g6�NK��ͻ�9%�F�P��~en@j}���^9�@��r������gesqYl�,��:7bJ����w�54V�N��\�\_r��-F�(D�(�ǁ�2��Ҋu�i��U�3?O4��f������8@����?�u96�O`��f���}[�Ԫ�K"x��'�y��5@ ҎIKF'fyH��A�`�Qk�	�A�!nɢ[��`Q���cL��!���u�.�$ۭ����YU��l��7vx�����ҷ�����L��70�
4����O�LDM�}'[tZ��B '���
A��2�A[(��kU�⚉dZr����N���͜R�D����5�÷�D�a�+�b�Z�9��0p���3��$a$$�o�)7�`-�
@ 'TҎk��w$H7d�����������\������9J���r�����B�}(���(���H��s�����]X��y��U~@�f`�����[���y�w�\��JA_�!z2�%�&�QQ9)�i�M�'�?/����D$?�`fg��&�7�G���c�=��[GU���I	E���GP����S'�aAj��&[#0_[���D�&��s��j�&����c=�c&����n2̾eN�tAF���EJAy|��T8Ⲕ8�>���#2������Ν=�<�l�!"\N�(}DbJ�ɒa�c�����="��\ s5%"��Xw>S|����M��9r�� zI��S�7�=�����8r�Y;.���hL�(<1{�٘V�I	��9	y�,�E\����>��Qv��,���V{��"��w�V��#[x��m���R�2��,A�1B2a�DO�aȖ�!R��r��{���O����_`hZ 2�GC���F����|j��a�b4�bR���Xt�!��Z��Ow&b���"F,>�9!(�cg�?X^V���@�D�RN�̀ղ�|B�!��Ǐ�l�+(fS����c3Ǜ7~�F��'�?���
@k�GȰJ��U�W^���0
�ZCcye퐍���|Ox6D�)Ĝ�&�0K\M����B!p����/��h����ν�.
z�5�a�"\:�:���	�� �0�ߧ��r4'���:��Dʃ��8�I{Hj]��ڶ���������3�8ˠՖk�jA1s
\6��+\+��c}`���{����s�`�I�g��%�X�E���?�5�~&U�r^��w�;q�Z?�&�"�D|���^EP�1�b�ya���%��������8�U��Y�����x�Ƣ|��r,��躌�b��(��Qk���=�q�K�T��������.
F%���O`�,��K�ԾHH2�ñ�;W���^�w���紅�L��F�P�����0�ct�O�c�?9�)t2�5��.m�F�=	��|�F��c����T���[kg8ׂ?P�Ka~To���m��`y���?����q�]�7�&�j��½�m|�aЂ-uho�0o������g�8T���G�N�Q��D2�4��f7f#Xc|Zf��QMɇxS�mG�H���A7we�-O꿠PEs͞�D��i�����%�:���t_n^��k�l/�/:1(��,�J��M:�$`�~װ;�W�Ӵ&����)��(TLq_4q )8&�ﲉ�3|���}E�E���D8�Oh���a��Ȧ��EE�^��rC�CG+��(JH�P��b�����Vd�e$�o?Q�7���R_�A�
?H����dDc*���ϐ����f�@�0�*�k3f�g��-SΆQC����(2��u2�$ːY����W�@��dzγ%Ǳ���8���L�gln�ʘP�t�J��?!�J��q��Sn�iE@"0l�:�0�S.��X����Ẽ>����޺cv
����+
�SjW4(�AJn޺{	t	�tEq�@�C�"YkT�"ց9�mcz�� ��#��C*̭�#sQJ��B�_M� aBJ��Dq&ի5#6e��.�Ng�j�>��?f�4W�J���T�+���,��r�T�,�c��\�h
_c���4?��V�:�
���>8��cm\����Z뚃e�|4,B=(X��h�E���-���=D_@`��l��l|�εb�ɛ�2����٫��Tѡ.�tG̝��Y��+����AQ����fe��LQ�^!�'��+�Ⰲo�>~6��/]�����LD��5I�o�� �zV�=��G�e��	��A@V8��t��+�͞�tɍtP����{���󂨳,��_y�Ղ�~j�	[�k�� W�hA1	�>\+|DҤS1o��E��Z�D�,p�Vېu��'�#vb'(�|���c�ъ$d��s���К<��6`	�Z�Z9����
S����w�[V@Xw#��w1j\�o�fXU]r�T�?k�t��5��;.�ɓ
��p}��c,���.���xĽl�"�bІ�	!�}ӧw;|���P��J�7�AA�΢���u���x\?*�觻-p=��s~%���p�ť���`���ӿ��F���<��J���G�J���rA��2�6�G���08�r���))���.E�^��b��ǇF�^'$0k-�����◌�%���K:�@���p�ڄY��Y�:�Wq ���kz�@9e�j^�b��)>c=�*��u�5]?���sK�v�!P���aOW1���<!�(rg:p�`Pi]@!Dg�K�P��"�X���)7Nv�=PjI���
H�M��6���b��O]g�z�B&t��>�.K����5Ͼ�\��[僧�%U]y2�&Ѱ(���u`SFR��o`R��Y	�W��T���(�_�F�f�-����9��B#���2�zSr�����I�R��l���#�@5��� ������	fѺ���:�&qF���w��6w�4)��54}\�6H��K;	����c���my&oZk����mQ��F�y	_YY`��[�N�ؑ�]q������j���V�	f�E�UJ��E�>K�#���`m	�3�wi����?J��*b}�k�V�&�!܈�$�F@J�h������n֟{p-��
q�A�iK�qrV�gbl(Lϳ�"�i�qew�����ي�H�dC�(�=�s/������6�̜�:L�3�%��FԳm���#�1�%�G���S��;}�5�Z������� p�W[�Y�.����ew��D. �9H��O?�\@zh��-�ƀ`56�Ҵ��0��YI�@���H���`�"��@טּBkZ��BI���d3s�WV|bOV<�������$�Mi7�V8za��<p��Sl�>[��4z��=6�}B�0�9���Z�i�#S��zr��-<�*� !/���H�\����|
��$�����n(F>�cGU~M��1��I�_�`�����&���
�Q�*Y��H���d����2lg��^xF��è��Gr��1gT�������3�
��Z����&��9��x?K�����ČkFǔ���o;�"��W��f
f�1l���O��7�FFj��L�E��W>>�X뫪�A�Lj��cD�p�PI��3�`=�ع����_��B�A(C�n��X�}�)�&�C�d�gބL;d�7�~7��m�Qv���{3]��+�z�J��*���9@���O3��X ���&
����֗�qm֕���Y7`q[f
f�FX?�%�΂���R/+*�ErI��+����%��;�����A����γ�T�`�fO�*<��� ���2���bIE�v�FD6��V��Y�9��F��Ɖ���c�G��`O	:Jl(xhN�F{�4���c�jB�0�T��s`pJȱ��Q~^ύ/3#���(`8��M";�^�� ʛ�1B�S�I0,�_U�V�cvH� ��S�-a9�y�-A�A��(%�(�H�ϊP�����HW��7k��B�����9�"ƽ�3�R�?<�	`�Q8�F���w����=]'����!����L�ciQĹ[�o��p.�"B牊�gH�
¤�y�lO�� �թ�-��|��"b��Q��cg�g��Ձ�v�7oI�:�}�e���&��.�3Z ��O�=��"���)w��\s�]����r�>��(��K/6O�{<��W�ő��>��֐[�0]���/��YcX/E؅��������-�&3:U�ơ���M���:���� b�!Ȍ*�0V��LK�G��x)eu]�й�#̊<�s�?�"�F!�#���,C�%��q��ef�&mxQ�[^�Z��q	s�3m{���6L��r���A�b�I��H�=�Dg�m�ցgH�KF�D dZi
YK1�ŖP�-���Y�2�ե�2zab��̇���b�"
B�B��a@+Q0:?�e���֜[���m8�����O�e��.!��F�0����GP��F�>�Rd��P�K�^-d�YA.4��`�Z���~|vB�C��S"�����zyV`}���	����UX����Q�.��4��T�.(�B�z��C%R[�	�+?�!�X�����a���d�K��=q`��v&�3�	A岆9�B�hOm��Z��ƵT�����.��qa�J'��(f���3�xF'b�����/�=���o�L�h�0<q���o㹈K�GkT��!P���4�[�A74R�7� ����R�R��N�<#E��QD��v���c��B}rg8J�U_NS��Y�pZ���z���v�B�-)�h>��Dqn��Kh�M��qm��q��ܠ�gK[�S�=�<�����-%�~��c�����L
�׆��M?�*���(3���`b9G�}�`jXt��X�������%.,�-: ��	�!:�F�����kac��G�^����W^��'�/r*�W�Ť�AC�j;ĞkÐЪ/t���y#�o?��mk��mj{�ON^�B�#M�.EW����O��F�����B�v#d�.���y*��+��w�{XV$+rڑ��D���#p2�2K~��i�Z�Fa�h?����c���wh����\�4����Yk8����\.�eX����ִ�S�?"K
^��s��\�)	�+���̆����1ωSMl��wt��<��}��ƮaB+o����g���N,"��\�me�X�@1u	2�Q���g��,m�2�{A3�c٫���?�k� �e��g�`Yg�ѝD�g�[��3�g��rp��l��|�J{x"�P�'����]2��"��o����Zk]N����ā��[��T�seY�\**��؏Äg�ؠ�8;-�r!�F9:� ���ئ�nEE-/#�D��ݞƾ��,.�m&$�H2���$QTʫ�-�$A��!H�3L���s�h!��B�O���
�V����执o^|���Z6�Pm�+�_	��r���=!��b6�|�F��{f���f����\�"� ���;���h-���������ڒ��g.�L�M ]��(�-���_���ܣ�}X9����="QT�ܳ�Ŝ_R��7�|#�(�D�����/�H�����P:���Q����+BtCbS͓g�Q�����l���5he��	�y��n�v��w�˸M������ y��d�?���8����+��dO?`0�"�j˖״o)єN��P���q�L%�Q	�r��uY(㓩�̍��A��y��:BAe�x9=��وN�y�l���3<�E�k��6�-��0|zG���9��9:?�ǋ�G���ʽϔ�!x������Ø��Q<��'OJa�!���怊Jg�W�w�i�0u���FYмPre<��p~��6�K��1��x��i��7�1���Xd��zNS�X�9�evw�B�Ԭ�3&����_�=�rK��-�AZ[�T�Ph*�V
2�&+����J\�Ut�� ݴ2�����p׆'P#�Z����G�S&
o�&��oA���������[��i=0��n����º���d8���̅���*����U��)�L���H�L���8�Eh�����G©�Z	y-"�Кe!�$�O��T`��K���m�2�����IU�8!�w昪��L?>���1�]���-~E���U�A�q��8�2R���М���(:[���ݕ\Q�+�^��jk����V�n����UH����g��5bj\�j���NK�~���A@i��jS��7�/_�o�rQY�Iڤ4�U)#$lS�&��Y ���8<~�d��>> 'Z�M�M���n� ���!I�N먤�0J�����{ӷ���}�a���xM�������<����%�klm��0���-�?�����j>ƈ�*a
ր�4 efT-������9b�щ�����)0x�-D�r�k00�T��:��ů���\�8���JԵ��t@�x���#����i�pn"s�>Q��?������c�U�>����o,�聨qS������� �=/~r�3R0�Q �s-�K�3�� )dip�sxL�[ő��{1t��La�I�h�;�1�0<��7ϝ�)�P�#���̽U�������"4�_�O��j.�Bt<q�G�#�����܆�S�;<st�X�8� �qR>�4k�.//D1�?��tl�_
J�Hg�9�'�qU���@�L�j�	^���mr%	G9��=�R �2�Jf�������A/�p]r��H�f�׉Y;̞�%&K�e�Ѱ6u9|0l�CJ��I��25���mΟyR=�8{J%�Iv�xs�ʭ�hn���Q:T�Ji����(����\5k;5#d.j�̂��������U3��oԁ��q�~�=ߧ H�J�5�fm�����0�c�j�h�Ʃ�u Q��?��ӡ\PŎ���Uu�8��t�������s�$?�9+~!R/ԐY��|N��	GmL|L%�.�?����垓q?_����t�h�9�^����ŋ���٣��e!��x&+*�xJ�r����A�G�֥�,�*��.�eX�9����W�hN9�p(��H�P�h�JҒ�
0N��w'����A�n	;ߏ�h�R%@�!��}����p<̑��׎$�(�#׆f��w'{��{�/"��8��1��1sMSȚ�I�8]$�(Ѩ��a���3�W�O�H@X��/�?2�lh��f��4��
=�w0W]��bd^'�؏�*Th��A)��_�9z`VB�V�Z����33u��<ٻ�֚�+��йtL�V�9�ga��G���F>���W�K��Bo&��Zڪ�gϚ�X��9���E� U�hI�yWNE�	���8�c��,��'cOFPOXr��T��zl��yYjG�h�8�7�l��՝�i�(�:  ��W�B�M+�9��>r(� ��x�<uK��<.FL<���c�j�¹�?�`u��\�#J�81K[���H,Z�-9���kсf�~FJi�s�l��V��_f\^t����Z&��
�� l9��!3[�	_�f�5p�.B;׳�P��+z���ܦ��0'U���~��}���/��9Q-��|���>�A�F�P���m�w�ƈ�H�����!�A>�e΋��k�@;1?��N���â�s�f�yd�_�y�e�%�wL.I�^o�P���bb2%R��vD�YT@Q�y�a3, ����7Y���ߝ�˹k���{DUj=8f���c�@oX�X�Q~�6�2EV�u�}A�Ǿ13K[�o� ���o� ���*���<[TC*p(�d�֮��,Q�Es�]+(�k�w4��W��^�T�3��d�@��U�k��`!�C�z�9�O�%�ۊ/���9>�l��]ӌ���.�P�j�5�U~ml,+�X���#ҳ @\�lm��Ւ�X�,�++�̙�К���:@��0JaZ��-AG�̀��e(33�B}����$�ܮhQUDd���	K{m:e�
�c��ښ�=�FQTj��b7�����N��Hbʱ�W.�f�P+�"�j�X	�!@gTI��2�/�~"	݊dT�8ޓj�t�܉�gΫ��3Ѯ���w��l�ݸ�jFi$�j��Ջ�2�qǢ��&Vk�&~χ	Ղ2B�uݴ��̵�`����0{3�d�����&z[�>>B�K]��}&�ş�Ǝ��F(�JA�ʅ'o��җ#�K*����Ah�$�3�.�x5a𲲣P2�q��	E)�7�A4�Б�5,�7�(�0*� Vt@���k�M�,�풰����*z|�l��)"8��F���/��b.8	˾$#Gi<�a�J���=���0Lwl@� �Y���И���Gtd��|m��e���9.�ͼ8��k�w���ź���'����"�O���d�`s�=����jA�O+VB6`Ƃ�X��0�I��>����5]���i𵥸�)�����*WiX7��P��~�*4��3��-Y2_�\�=�ȈY�~��y�E��i�������Ц�+�<�`X��|H�]ČyMZ���4�ja��Դ�kzwY�Z�h�W�.B7�7�1��vk�5R`e5�c�4wԵ���<Z���5m�;z0��c��-�g��d5���&2�_B��kty�8��~h�@h��
�3��:�����u��)�"��Z9u-��}C��I�i�:"�j�nZ<�2O�?�w�T�p��|����R����9����i���@+�P��9ϗ���0�7f{�
%�0D��Ь�����8��Z ��1L�k��ovh�"∔���"����H~�H��7~��H�����6N 9g���O��M�HTb��e�C�0\�rU�Y s/�M��<!?��i)�����@��A$��Q�c�c���������7>;��Zs=�y�N!IF�֌��̔�P�B���[��q��	���l]p=��A8���0iّ,��ʑ��v�"��]\�I��\ւ�8�1��� ����d_S��Й$��p,�!\��[�uE(�.m ��ˎ�t���s\G>`t�Q�58q�"�Rpw8Zz��͆�s'�I�;ɸ���Ƌ�͖����p?�J$�������K���n��Yr-�:�E��bY�$�u�b����1�TUI������z��C��X���n�5�sM�V���Z�yƝ���"��������h߸]cU���u-�P�Р���n�`3|6����Ӈ�	���Y�%�;|z��>]4.-�B@�<)�- ���J:������=HO���Q��Rk�զ$�q�i������3L������j�rS~1�\�yM�1�h(�tHA8�y �4� ��brBn�� V^��1�ٚ�}%O�Yjh���s8��2F���^��G���5Ӈ�}�����ODZ��:�o�j@�����7�}�A�%�0��Z6�iZ����PW�׿���e�]Mh�Wt�!	C����I""P�/�!�d~���T����Y����iIt�_9G]��a�O�V`�#ET4� ��[�?�[�0%��ώ�-lR �ԡf0w܅O���3qnO�ũ�F]�����o�q��o��HB��4�Z���������?&c	���ho��}� d<3%��c@�q�&��w3Q����Ψ�����,]^����jv�H�8�Gdd�f>�.�⫶"�=mA���ѵ��2^�B��K(��ן���K�,	9{b&�Y �����7S(����P
*�����$[D�f��H�Q���~�7y�),��7s�Ѧ�d� ��}jݼ���G^|����=Z�aS���vB�74A���U6�ohx��?Y]MJi�亢�E�pI]�ggey�NZU��;j�t�ʵh::��M�,�
L��bS-@RU����D��ع����l�L�r��
�x\mY�Wx��:�_��\|�

��@<����iW]�h��S�W�Ps���w�P�(� 3�Z��K�%��jׄ�cZ+%�O��,H��$|3�n�%L�F��~�Д��ݭ���n�Sٮb��}�0��.�bOBW<e�`�K�t�8,�$���O��G�@���:e§�k,�1��Z��i������r���fk-@z�ЂqF[���ݽa��uHw~�,l���� A�{����PL��
'���0[,����~���;��NNap� �2��-k	D����ys�w%��K��J_�p����#����1�V?�GB�����f��P	�T��<t)(�2�q�
s�
9�&��2hz�p�"|�o�N��?KM�L'1������"
�/B�7��9������hZ�.��yK�G[$�����ʱ��>�y6�j����8Y�%"����^w>lД��5��dZq�G�iOx�2O	@�r�m�	,�DU�o���]��5`}}�+�SV�����PM)]*����Ɍ�U�EM�6	���d֖G-2�f���	 @���G�.T}'q��n��T���٥�F�/���+��{lN9f	���X�3耱oP�TP��/Y)f���O*���s�4���i.����Knܼ���(�ư&W�������äB�5�Z��XX��6�K_�P����Xë�?�Qعק����ײfꟜ�wz�(>R� ����{��O.5}�a�W��m�В�N���=J�7\%��_�<�]���ޅfV}!�N�B�:��s�^���`$��"@�L�:�LJY�Q�hOǘat��vUĂ0��dh��D X�4�M�+0l>Oa�1]�~��>f,`4�����p��Q6a��ot-`�;������6�}e�]�4����Ò�{'�;���CXq����.4��B��2�u��c�fu �F�B�(:�FB?��T
�T!Aа��wU�����H�[v������|%��{Ȃ�U�PL`�SZʱ%�R�!��iWz��i����S�ōpI�x#E�j1��"��I��`�1{�� ��C�_�U4�n.:R��5:%,�f��ο� �'2o�+��`2�kÝ-<	;ƹO�(�.`+"㋰�U\�;J��"�t��
�� #���4�ÁDT�Bac�H��g�70�>m�i�i��hY�"L�{]QE�Ub� ������v*����	��g�(Z�D��E?BA(�R�J�}�h����1S�g]�������4�_ؔ0�	Κ�IҞѺd�����"�"9UU��lR�?=�<A:O�m.<{^��.˾W�9}��F8��T���:���hݓd��kw��f��0$`�����ذ��c���uf���Ԃ���v�KDM��K�Li�� ìC4lZ(!ݙ��9IX�8kI1�ɋЏ��)l~Lm�H�G����� ���`l"�</�(&��@y���T�9&�p��.%qf?	�Z+ ���8љ�����`1��z��
��|�yʀ����
f�V.��5ME-|��j�>k��ѪgB̕� �j�	�N 
.�"�R����.��-�(b/B�bYi���>=RR��>$R$��?��z�΁�Y/��W��O'y���`	E�k�m`�ZƧy�S#g�;8)�)r+���'��w~.�2D���i����a�ŧι<���2��9��9@Prmx�DZ��'��M��|Ƽ�5����u#ٞ��[E=�`�c�_N�k�������(��t��aM"�W����y4 UIU��L���/���'3�*c!"MB�&&�#VB�RP�h�<\>h�*[��iÙ��4]�Pw� `V�9:G���zbu�z��~J�T�z:�t924�T >�>m-��7�n~���7ȥ�B�o�ͿQ{-5O�~6.N�x��F���z��Iʨz+���C��Ln&L��J�ѡ]#J6E*=�Me�# �IRD ��r|���xS���L�X�z����!������<V�z�ԃ���c)p��8�Zb1��/���ʖR>h�$hs}S���*�6��K�'T��"�.kN�W^�w��!I�'n7���h�� fu[�o"��+�z�c�z�`�0�(Y��#cቾ̰�L6*dC����AL��棈�.����N����b04���YJ݅_k%�M��R!�(*�k��S�z"
Ќ����L���[��1�Yi�D|F"������ҰU8]�yRsq��O�E��΢�e	�uz��B�1&���-��LSٳf��*Z�������yz���@-`�r�@��l�%�-��$e�}��HL�}��F���u�*tC�O��� vbB0?~�@��q�aZ(Ww��ME9;�!��0��c����j���s�I�oR�f� �Tbo�J�Z,R�!Y�j����^��NCc��Q�N��J.��#������ˋ�az�mdaj�gp�k2��/~���K�!,�V�a�����Ga�e���Ppy�?M Oa�j]�"0}D{A{ �Ek���)]rĈ�@����T]&"�i�~PJ���~�)� +BK'�RagGl�`r�. ,���~�sb�7���ڗt�A�"�]��@D�`���l!�����3�!�=,?�������z�HоT�c��H�mA:���xsT
2�k����)^����߾uE?P����*��/��o"��|
�����Lo��ho|���we�/(bE���6�!1�v*�ѣ����uY(>O39�=h�$#a�ʕ.�)���XS)��sꋦ��Ҙ$��{EX�~�F��9*��JmU���aE���j�����+�mC97��"جhcò���`���T���敯�Ҽ6��X�swn5��=�����ʽͩ!���n4��ns��jr�����t��u��#�xvG��,&q�T�(�ݍI�<�Ԋ��;����o'���p�0k�>��.���g�L���mK��:Q�<�DeZ6�� ~�-$��4�?��9��t��y�*	�))h�XP�
X��\,����: IAM�
e��8X2<E[�`�MS�a<g�\Y"j���@�Ea��������2��%"8&�;� �B�{�p����Ȓ[��V�?��qh�c�0p�FB��R��>�܏=���xWz��,@LԊ��1���[�54�u���Z��9����{!�@��MC7�u��I���A����}�:���}���v�&�6�G�8*�TȂ�1�ȶ�	ç����uY;�GB�1^=��|���\�R"P/�wpLB�B�bQ�%��ԇ5l�5B�h�S�ϊ*�D�k��#@��'@)]ˎ@�)����/���I_ �s?�5�'��3��2|ׁRd,���w��LA����Z�����]���t$���>��I���n����T��È�@1{����x4�l���J�ߠ�g��eF� ��?��������5E�4�p�(����ܤ�z��z~;�?�<���-�$(�L2���������V�$�W�Q�A$�D<�	TIR�1i�S{M$�nRW��3.�WB	�+" �y�J���o�I���͋�L����,AU���ݛ��g���vss���D�aQ�x����O����m��D/�%8hA0	��Ά�0�bbߟ!6*sƂ��	�0/����¹���q��V��վ\�aW�6 #i�(���	z�T�AzVח����X0?�m)�hS��O~�_|�+�I��zL�hN���2�#(𦻖�=��x�� !G��GG�Ж�G@Gk���'k�}��[��%�&?�--���j�Kff������ р��ɼ�-L�y�D4��e���>?dI�����X\�f�E�##}��t ?�)F��`��n%��i��9��]t:��D��s���	h:vwG��{�q#t^@��o[2v#�5�qk0!��u�pТ��a?·�_�ӂ����%[��be%��tILX�`��1&x[fE���)��sZ�[�ZOЎ�9��"J�q�"�56~C�Q��x�;��Q��e�B�ѩ�.N�n2�:Ǘ�0�/K�̔(�/�X� ����Ri�X �MaXٺ�8��9���_�,�CT9�9kA �\!�Zs�(�;��R���{?!��TPkt���_x�!�����������õ��P{2���p&�z�b	F�A`q�p'$`�}�	���a���Hw%�֐hXpZ�1"��R�Up@��F[ƿ�97�*�,�R�4���j�-/_�"��q� ���z���+Ͽ�S����|��S�?���ƻ�y��9{�|�6K}E�*�͍�}��$N�<���	,���3�P��Cr��[��`(,fmn_I���7C�H3��{_�I�u��	�Mƺ;D�V�y�����_�&�y���������0q�������L�|��H��i� `-�H��-�~��o��mF 6��AF{Y�Ղ���W��T[��������=S2B/�]$�[X�����d-���(����/��!g#Ne�߇���`��a�z>QN'�9��/��1��B��ڬ��,Ъ-�Dzh���2'�l���Y��0-4�K �l:f_�r�-Vn�>
L}M)T�P�q4(�O%�{�����ܛƹX1׮}&�Ӹh/W�q��
����D��9��ۛ�'ۮDkb�y��l�׾KC�Q���u�B��Z�_˜ 4���f�i	yf΢����y�?&���:����k,��,v(�������b]MH�(�19��㓥�~� ~B�햠v��+��!�� 
�\)
�(S���ݼ�g%&ҝP��˄���p�䐙�C������j�q�Rn�e ��br!m�h�(�ew��C������E��@��ǜ<x9B��i��]&T����*��c�>U��ۂF疛U�>Jw	�f7���M��� i�8$���E����lɲ3��D��}��" $�D2)R�X�c*Y�ձz�z���(麮�;ԍ�t�:)��l�ѷ��~�o�k�/lx <�I@r�N��{����l�sN�P�2���G�����d �K����"�=�v�M*�-�v����{�>]��K�_kP�!c"nZ-<+� r�<��z���8�>o��n�:�|���=�>�J0V�.J�������b�5��ΰ"ñ�,��=��ҷ$��5�s$�(��%�:j���	��׿�u��TĆ����R
HS1�h���}`=ec�
u�,*�����j���tJ�;&BcX�7�˞�[����M革�|�Hb�7c��5���Z�[a�jJ���]=]+)Z�|7���cX���(ݐ_\+OQb��e)�/.����%�/%1�J_� �T��(?|֝ @����Mp;��
I᩠?�*a�`<sG���B�p���&oN���8�>*��p|&��ƭ)Ҏ��U�q���m>�|�y��y���3.�l�� ��ƹ\7ϓ=�z�6s��gJ�Z�-U�����'�v�=�5�mEI\A�T��������c�Ö����)9I��ZV�87����z+��
�t:���O�cs����O�v�VT�`[�D������D�{?zR�POP%�٪'stiy���Q��m��?��^���2�;C��{�wm�7��&������c!�����	7�y4J���n����_3:
|�o�&S��8!Bnd�8!/�!}�P�R�L��k}����$��
����M@���;->�z;8vapO��J������b�B��]�G�H�
�Wؼ(�.6���ݗ�h�_����*�FH�c�Ep�Q�	<�߁x
�`A�AT�;ܐi��(0k��}�#�,����_AÊ�ȉ�?y�φ���"-#��wP��C��� GNF�36��N/N��{x{�
�����i�w�w���W�Wo���1�w��"\��%��MC����Զ�����y��N�[�ŭszu(�G��yRV(�+���\;zmz]�#�5��+�>l���;?��u���ʽEqD��m���Fĩb�o���~O��=��u+�[y`�*+A;vPɗ�޼_)��x�/̞�Mo��ba���id����mҍӽ�&|)��Z�s�t�+�i!m�Ӭo/���i�|��	��(H����!:�x{nC ��gՃ2�f�ӖN�q;���q��zZȋk׮�GD��j�2��'�ϵN�@IZ*��X�DcA��M�ȴ���@El��B;���x��vl�����|k<�{�UC�|�y�s�u��M�Sƭkf�^�z��ط���!,q�\��8A���c�g~c�P�I=	������� .�,]���4���,K�u�V)VΠ
���Z[Z�����N �v���,���M_�?-&���R�7��	�0���L�}/*��.9�b����7�����kx~�����o�;X���׷?�_�7H؅��o,��--Ua$�J(�U}C��RA�ja��R�q�����)|ݼ���)q�a��u�Ӌ����[1W�'�2��Iv0γ�����ޅ/J*<=?c�	7�c�	)d[������/��z�99Z�O(�'񦞝1�E�B��ᶴr��;
�PrƲ�tf�w����+��;�0e�G�P�ROln�׆�[� ҋ6�w�t�i`��u�O����C(��S�$1{�`�L���J�+�6
Mc̹0>�mC��c�e_{�N<_����vwHM:��|���U����nDV��}?[��	�V��{��2.��do��[,����=��.ky��'��c���w]g}Ŝ�'�ȳ���d�˄�OP�E'��j`�~�����˫E��n���������c�F�0�_���cZ2rqai�/��)��qzwkV�1���`�d�L����-^y�Xl�|�%�S�c`[���Ugr)��= �����4=�x�8��_��Ԭ���H�G�<����Ɵ%=��qur���5�9����c��QE� ��K�Ip�l�j�*u�ASIi駁j6��ly�&F��TT���N,^��Ry�b�l6��o�.�������p�ls�5���p� �g�1���aq�X��������ߑ��k��_���H�,H7�� F��=���[��L�d�y�_T�i�!%�U����
��-r}����C�>��hE��<F'%,�(��%x!Ӥyh6�j}����'0Y6�x�����^��X���ZC����24�`v/H�Rk_߻3�
+�+ �ϰ`��VΓɸ©�PJV�Y�g7\��C+X�u�9��d)bsC�����*�UFA?�2����>�|�qT��������XK�$ާ����ȇ^��F��3
:�����u�8�>�<�kn�
��箣�RS��+q��|y?d���L7�w��~�˵�a��e�<���K�G�����[��ҹ��&� �;��94���4�;�Y�Q؛Q�Q.s"�j�U9.��*Y�+%��s����_G����2��O:˚;ӽ�߇�G�B|����5RJs
L2v��-�XW����v��U�l��s�h�����~�ھ����=Ǡ��P:^�p��1��:+���p�i�_��/YK�����=d�����g�P��s���	%)�E�M��!��vߺ��-�
TrGt�&�I.p�n�oT��o��o_߽SF�;(p.�z��0܏�#d�L�?d�'.�^W�E�ɥ��(C7{K�o5�N([�,7���Y��,D7����M   IDATN�S�C� �����ǥ���IM��d2��e��:��*�K�^�j$x�. !����*E��<���������w��v<X�YL�65�p��2�6G!���"	��"q�{@��ҏ�M��6��Mӏ1Zq�D��,�b��+MZ9�o�izڪ�ku��(������}~>�ה�Y��oo���
��<��������]�x�}&��t�pN3Z¾��x�Pne��l������\l���-���/A�pGh��^qXȱГ*��l�܀շ���	��q�XD�2�<�y�ru�_e��S4�A�^H=��g�RZ�?���X�(J�Ė%վ����굫�o�ݚ
`��S�1r�����<��œ	ZP��0Wt���M�u��!��;
6�]����l�d#�xM}	�QY� 	O��9F��?&V�_�*�9Q�.���q��Ƞ�yT5�D�����<Is�SX��y�g*{-�Х"��Z��n\�4���$�����=�������(�36f��R��;h���Pr�0�'������%�������mֽF�1�c��*j��^�
���r��͒;SDZ��V��0P!g2=��G�`tV���^�C>{�?!/�(���Db$=y|�8��2.<�י��rv/�����`�1��4�VV���
5=�� Ճ�����qȑoF�o܂�qM`(��MOM�/��H=BΧ�"�c��IM2�2���drVr$����T.g�}�G�L[�D!a��!�ѣq�*���O�6K[�k61A���O��:���\��v!h��{�[�bkf��Wy^\��F0��"�����.���J��&�ٿ����n}H`�	�C�6������a{�3ĥ�#�-7d�tbu.�@�>[��{�1���q~@�J8p�)�K�M��7�s�ζ�m�|��Vr��̝����HzȦ�?{���-d+%i��b�9�-�\a��J�:[ج,-�R�<ޞ�!���_�v�����kp�,�K����6�X���瓧���>�_Jd�{i*�������v�k�̍5n�k�OV�5�d|��0D`,e�����8��+o�q�Ҳ��
+,ʸ�R��k\�_�S�9���Ϯ�.�J�b���t�vM�qi�陴��b�Qb���5�Ey._*%Sf�27!o�w�z�X���-���]bd�Ō)x���o+��L!��aˠ$>��=�ߎ�s�\��W� ��xL�z�d���M��>�'Ҡ]=5Ϊ�e��`��J�nl�m3t����4���/����D�������a���~Ha	c�>K�]3µ��kyz*�&C{�C9Jg��w�)����)h��H��Oq���^;�ica���@��Xd�	�1۰�i�W$A|'`b�+�`	ʅ%`޹�"~��z?K����2kV3_��x��5��<C���!c�f_�}Cn��Y�'�eۛ'�����"ǽ�����:/��Fw89.�)\9`rv�y��fm�f���.t'�Բ %O�bTOx��	#��U�����^o��9,�Q��7��/��j���ot�tI��Y=B�!���&�*4��C�~�����nS�
N� �p�U���V������R\e�xd�) �L���FأOu�H E7���M��B�k[�]���k>̵RH���F1�N���{;[0ߍr�
F���o��(�
AKhP0T�nҎG��^�o�a���D|6�)��_q�?!�_��a�\*(�������ͽ�˯��h��>S_��a��� L*,��1NԄhk��w�w���4vT}/��䷩�S;�߉�y�d�+�����Q���y|����+��ʸO�:��{�hK[���(��CZL���ӧj:ŭr��N9�N ����l��$�=z^�c����	S�g�{���T����[�w��f�y��[糌���}��*��y�A���4m�$Hg�t�T��������X#�TI3x�*Q�W��3Ȳ_�(��iA	�����zc�8�y���w�}o�>�xb�)2K1Vۏ�>}F;tN㝇w��*;�ﲶU�~�x���Y�`y¶�}�ؖMV�
����?�9��?�2�U��?�T��88Gk4N��`\e}-_ZŰ�ß��x�zI�3S�87�,���EHK��5\a5���ͦvy�I�@i�h���87F6q�puTAm��)�G��<���j=�`	�c{��&&>ł].x�U���Ki!kl��(��>_A�(���XmZ0�����W��^ƣt�lR�M(C�z��o&#2��gb;�I�.Z<�?@Z��Ź�* ��)�PO�3$����#���Ũ���m��9_K�\ ��
�VO��GV �~�bSg�5�����{�}�,�&**M&��QE&\e���QfU��uHw]	)�T��g��P��b]���L§E��g�t�t?D?��X���=f�ϼ
EM�2l1�F�'1a��2Uv(Z�*#�e?O/�l[�#Z���_Ni�#���x�3�sג�6�{�W�O�ROS���U^�/D�K��JR�Q��d�6����C����q�=��>SU%V�Ԏ�(��	��1�2��{��(�*���ޅ���*���"a��kIòR
�;OYO�a	[Wx�V��!,�`��b�k�u�[9��lƄǪ������wp�Ӗ�w������"D�������
c�}*��U	�������=x���g�Y�,���L�������}��mlN׉
�gU	�������8_���U$#���5@4�^/#��s�����_�h���p?,vR���V�bFf!��.�2�W����.r�*F�x�A���+�9�7._Y�$��ǩ��Ct�����	���;A��;�NBy���I��wY�
tլ9;FX�F6)�K~�y�c7̅�\[Y�&!%��x�&�XL ��5^5 �T@\�O����]�6�겄�sL7��IY�@�B�*:@m�,��arMq�+tF���.����T���c��*5y�2D�u�'��l6f�&Y���z�Bꌍe�e�X-j7\	��'�uۘ�^S��Y)��g���[�|����r�S�WpQ~%�-P�o�]�Z�9��'�]�%�ۍ帩�f�!DU�a��Xﵾ ¾�U��V�YY�]��R�.|:4��G|�Y�����o����D+��O`=�N��21�F,���ކ�;J���1UX�3���Tr�i�%��LSQ ��r�>��8�<9v�A�������{�x�����,S��{�R�ZP�c�-�]Ks��Sv�{P����e�P�A�}#3�$1Lׂ
 ���sV][�{�{���^��~^m����q<a˧q�س�.Eȱ�b"�h���d�$�.�'��X�x�������Q�i�Vd�V��sK � �ܡ�@����ƾ�?��������WOOC�B�r��V#Y0��=�����z��C�ڕ��
OP�b�_����*5>[�� ��l�3��^��CNJ(TYWo_D�p��т���cY6�­�mBs�w�'Z�>3y������&����и�r/MNϭMNϞ	��ڱ��ƠQ&��3�~�h�f�8�.|1��Ư�@6��Ym�(���1���H%x4'�Xo����6�a~� ל�0�ɍ[Xk�s��9��MR����Z��:�~X^��V�U�Zo�I0_�EWM_C�߷o�S	�3L�	֋^���߂�3�G8
da��hW���0�e�>��6�dLh��;6>c�+�@ub�����a���	��i��v�xF@6�j�H�++��`�!e���B�{C��������8��g�S�5e�#1&�r��fMՍ_��?q�v-^CVI�������﻾����M��y�1��w�<U��a	�w�]�/�]���D,��H���2�b&��W��NȨ���u��sgEiB�~��w�=��|���G���b09f}�%W�!�d���PB����3�Qp^�{R�(D�7��"̿BU%X{��
y�Tp��B�I�0iD1�XOE�T�I!�Y }���}Uh��3.����M�g�C4F��������a���1m�VPB�IT#�"=�x��O�;��i��6қ�+�8�X��9��?��BD����ץį_��*~��.jr]�u�/B�-�9R�	{z�=����TF��sal���]�M����0׎�ޠBt�c���c�V�I��zʢ�e�j(�%0޼�:���-��$��� '����<��ף���/��YX:������ȠW��!��G���Q��ĪuS,����dcb��L��]����bA� .̐kF���'�Gw�⽙6�D���}�H�L�E�G�,�o��aqA���"�`LQV�^��>!m�V�o�C���������
�R�p�&P����5��<��v��)ޱTC*���b�8Tܱ�m�|�p�3(����5�3����5V�����+�����C��W-��|ޑk�u��|�ĕ}�Z'5��q�$�M�����w�Ll��pnMS���;�Y�_u�Hr�þ���/T���%���2�(����h4z��Q'��]�w�bH��)���d�)Ȣ�
��~�ښ~ǸN:�{�c�P�bL�j�&k�y�-o�H.Z�]�3y�
��ƃp`��^#�^!܊���t hTo"�������y/�6
���\�������x������;���;~�FX�q.{]��|1��K�� zI��;��2��:����j���R�a�7o\R��4����L�Ѓ[D���
��uy?��2�� ����a>�Z�Fa��;�����-h5e}f���iKU�I�.�_?���e���8`�)�]?6#��jW�b˶u�;l��T٭� i�{��!:G��s�(�P�����#��j_|ye(щ���!&^LC�� �����p��7��D�XƁH��RI�.� &�m�+�� .�T��0w"��x��1���B�n� �Ϟ���]�
�RL�S�yQ�Y`˪"S���`�{ON�o�cX�G�ߗЂ�}㋲L����lWg��Z�彚�.=��
17������ I����#�eţ��t�g�Fr�j��!�W{��/�EW�t�ښ4h�	��*�4��"-��Ll���l�Մ}q<��^�-�2u����A�&e�؂�BY�Ե����8>o*z����,��9ϳ�r�3�:��L?<�y����\ <S�;r>�$��z^~�$�BH<�(�(�\<�1��y�1�V MG��_�e(*a`���@ar���^Q����6��t�HU����;/�}�0�G����:1���1�=���X����V�4ű�VB�Q��\��1�=�;��o /ܓ*������P���ރ��aZ��s��J�Q��ز��1���������mb���@���R��<�]��[�n�߱k�M���������**�7�����O=89""(D�2���8�>�W�K��ZH�Љ�i���Y��gN���.yb=RJ�&*��k�{�ڀ]$�Ҕ�ބ�oZ�Jpfn�gh���e�²��N?��o�����9C�[L��	8���|<���193��T��/�',�V�+�Y���^R�}Ȧ䚲(���#L�(�����6��*߬z�	�������!� ]���q�R2�i��D� B����!]^a��k�SH+��U��FL�#�a���ƍ9�U���V�i*ϧ�e��KTv���M��XA��SqA�@�[_���Φ��~�_K�W��U����_��_L�����S�����ؕ�:�E�R+�?n���PY���ѵv�j��%��s�R�e�	��擶�mҪ�op��,�^��j�v�(��K<6?����yp��R���x��	�Y\��_�+��|+4��@�Σ4A�*J�֘E+�%���;Q{+�	�%h�V��S�����k5(O��xi}ơc����=��D��YU�!�M#N�⵽G�aU���q���3_�ysϙ�]J���1B��(����x�~��C	�(]cJD����Ub�z|z>��H|�.�(8�I�ewQ����iҺeʞÂ���d*���{4%�g��� �S�Vt����*���#����n4����`����^j�����'����H77�<����n�]UP��`a�~�߱�<d�2q�������f�-Ǔ���"ݓMl�	c���8x�=
��Fȕ2 ,��)��$n��ԚC�c.��H8�0�q�YaY����铓��m���J9�����K��^6n(��&q����ڙ}�4$�@��V'~���,�{03��3<���#�p��B��1U_�=~>ؠ4�	�£��$��
�+��?�<E�N���Ke*�����a�Sy�RiL�	E���Z���X?>ˢ���<�-aL���W!/���g�a�7���
;��O6�2���G���F&֫�e�jP�U���&�.r7U�����E Fx��MFK�rlVnG�;����&~�'��x��\��Qb��V�J���e}atp��M�R0s�cjͰ�d�Z�_֚�-��TS��}w�?G\�/�=��P�@�hZ��T46	�:�,�S��"�!�l;�kd��+A�6����1�v�m1j���*y}�t0�'�@�=�.%dH]�%�^Н�'^ib�I3��x�i��c��y��[-'TH/?I�yb���zܓ�koJ��r�ؘ|�}�3�o�F����o��t�1Uâ�|0���_�y�FO�>�h����u���[�@˙���'���m*�[�v����^ڧ��|��z`��p�E�iVS�Q�)�W(�r|�u��&�$�+�+��-������k=}����O�t���Lw�D=����v����@~Ș���mხ�gW���/���Z,������
���ܸ����sW�D	�&��}�g���Rd��u�C��e�GټK��g@�w�~��W�op �Q�s� F�y�������%�:��ܐ����'��Ko�JcШ��M��$�ZEN�t�b>a!$p���+G�'�/��a�����q�XN�1I|Κ������7�j#\�J:°�y|�.��v���&�(�|�´n��T��h����ɕ�k���Pa��$�5�m���.��y�OE����6��z� ���1���t�k�0Q�r���r�w�	
��#T�����������H[o�q	��������湒��ܸ��k�{il�o)?[]�Y��[�0J�O>p����B���cb���n���2��z1>�q�X�o+��2�����2	
��E`)YN�U3LH�`���C��@�Q�I�	�3����yMT�c�Rj�yLP��}�+�� A�P������-አ^/~<K'2�{?K��@��_���F*)o�s�
�Jޠc�����E�x�[x��jM����n
�y	�$��,��������U�7�S$_�g侅h�ܿe�u�Y֦��F6�v�O0 �^O����"L�^��貜��d��X�N#�r�f���Z���ՠ�H��.a��s߅*!G�@����
��������g�}Z���g/�����D@[1|e�������
b�
9�Xמ/�i$�ek&v�곱kar�%���5�@�L��`8���A�~�p�E����x=G�N���Yc����	�QrE8���<��y���b����'����8=B7�D�e�c<5��`��X��vl�M\�E��Y\�K�AZ����6�1�S�ź9�{�#h��1�B~j�kSʪň`~Rɼ���F2hd!6;a`����K�ӹ&ͱB��K�!̷Ѽ&��ܠ�p��8��v���d��z�Zs�]�T�,�FQyC]	�@_�E��-�����R�ݍW!/L��i_�����w>s�Zq�!P�ϝ&�~!��¼'(}�o���B����1�_5��Τ��@Q�#���g������
"�3���SȒ�T�ذ
�����g��<E��y�	�FB�.X7
@ϭ0u\=>FW��IS	!'�Tcg*�:�[��=�{g�q�?>��typ(���Q�),�
NE��`#7|_#�r�ʀ>��qu�r]�t2�#O�ߔ�Vy��}��7h��`�*^䣲aOa|�_%hn�&ZS���U~**�ץh�uίguO�ؾ����>�ǴvT����*���������Ҕ����Z����Sy�Ny�/>�F���(�>����g��2��ڮ:�9���CI�h+	7N���@ᒀ0�'�|k=���um^n���`��@�s7�Dh�<Q��U�ɟ��^Q!�����Q��3X�w`��&3A������$�F���
p6�b�BM����lޑ�Ù����.�ިG�">d1�1X�,\�E��2��F&��Xӛ/�%;NH���C	L�1B.�)�#*W�۟L�3hȎ݃������~S	�Ҕo��`�2]��V�'j�2j�i�©�2L�JN%X�A=�R(=G�/W��=2-��k���)k�RqǔI8�iɼ�gY4s@'V�XBpT����U��Iv� r�f*<�͎��@r��������~����y��X�·�e���aXz�W������X}�j0��O<��hB����!�%v֢�3v
�����C����H:1E�s�zd
��'��Ea����i�İc��]Ij<	�	���#��u�q~G�D�:�d���/�Б8���:E�=늂r�}/����/��%jLJ4��V�ƫ5V�-�Mf#���x�)'zR9��S�rե�jutFH+���1Ce[w�t�N��b\Y"�P��S��9�4��E�d���iڋFk탺Rcɚ� U��}o����@S�������^�f�4�5L�}�7���u��6�L�^v>SR�y����_|S^�c�Q+)J�l��CX����	��x����#���1(tA"W�X���=�, cE3&A��,(��R��-#�e�a��x���P�x��6����4G[;�^��ҵ�!rr�%�o�i�xR#y�ϵw@��h�qgrv����̏W���T�.�c�a렾 ;M&w��&�VbWI��och�N�j%X{��E���4�k�*|:
c�����w�HҚ�����[��*�f���N�m�Ϭ��$�Y.���R��8L��ȥU$�Q?'j�sbQhi��U*��-�"Ԡ�W��*�U��Շ��^6��嘸��
!���TX|���v�9CX
��3��q�í
��3��1��RNс
�]eo���+��OY�oGK�'�.���l:!���mEؿ�&��V��r1iMp
:_%�֛Q8�����T�4�(���<�����uc�Z�AW��<>Ɛ^OWf�e��CuMy��W����B1R]�AB��{
|��H����,��^RZ^X�T'��V��ޓfo����]�<c{�Y]�~v�����lZ}ϔ���_�n��o��TfcR��$���xm�$!z�����w�(�T���x\k(�O���o�I]S��8�G}T��}��L�Ӎy3�B�۱�y��y��e�k�O�S��qj[�E�l�@��D�2>T�����۵L�2�yX"�(��yw�i,����f�dΧc|��:#˸{�FU���K��^B��OH3�p�sةx���~7Ƈ6R_$�8q��`g�h�
�0��R��
y)1�p��v2C!�щ�����n�|����<�7��F=B6�e�T���3F���, ���7�&�&��I<�PАI�ڠl�	#�ot�)�.�7p�}����a�1I�\��ED�&g�������ߖ@�ʉ����ܓ��{>B<�R�-�̄9`�1�VQ��%��rV��cAG۳ ��kxVZZ*GF��y���9�轺ܔ�8��r��o�gw���`�*�'�/�"$ӎG�!�+'&��"F�5��΄�Zu��i�gQ ��_���F��;��|��&0{��Uw��;�<��q��Q~y��|�݈O�c]��d��Ť��$j'+�%����Y+zXY31�Nc���R�PBO){L����F���r�4� �.D�y�I0דH��$�����Sv$���2Ub��S�{��(�b�"�'��E^�^��{O~�=>�
�0�i ���8�Dt�CS���@j����ݩ��"���\�:����>���а�1� ���w�A����j:���<�?�@*�by����,^�]׍y��UxO�1���u,c�M��gJ|��j�.H.�a���_u�ǧU5����;�ZT"57� ̅s�T9�f�wZ6����kɜY���5#�! �E�W�(���Z�i��I<����W_ѝCE8WC�ش�Y<ѕ+��嫃��K��Yƞ��	�Z��f�@`��Y,t>2A�k|��ҕ�ͫW���卅g�5A>$�jY�n�X��Ж�]�0q�T���(�X�.�(ʪ�bRr���Zr���3$�75�{N������������yȤI�%�������4 ű��SI�Ҍ�BU9���=�'��?'��d��e�Җ�XF�7-���`��Ě��F��'�,���,��ҫ툶@¢�*V���"N/�5�!�!������Cܬɵ
D긅䠒���w�욑��n?^3A|�*>[�Bb�(`�S�z�Vq�;c�U��_����)!�(Կ�������<�g`(��U��E��c���g�#��1�~K�`-#��rW	�����9�o_b��w�<^UR<��òd)��~����dy>���z���~�c��I��
0]�*���BH�����E�$|v��}ϲ�],4�>����@�z�^G���C�
2��o]`.v��{N�kʳ������-#�R�Z�cC�ΰ�����L�e)!����7T�����D�����v&u����!՘ľn{1�ߊC\�4eT���}���qǪ����o��5��./:���TK�p4J�M�v�2�l��Р�~38[M���e|���{u���8�.w#kev	�u�n���E�νG�O���x=�ߢp��%�l�ҕ��%��¥����m9���v����>�k�F�ץ|��mC��N*G;��k��������#�&��aQY���(��U:��0/KG��e��xa��c�r�MM�%3I�d�6 W,��4*����.>��|���E(�b����UPqc�K5[)C��(�I5��o8����x���R�{[X�T�hp��l(�;V�(c�^Å4���Y��)(Jc �,��*�4��XV<��B�p,���*8�<.��V�V\⃮��o� Z�n!������a���G�%AK0-e���sӇK?N���G���U���̿c��c[��7Q��s+���c���jޙ�"(	=aQk�Dg}�=hh���ģ��� �󐝢*��C L'i�V���]Cz8);f�����ڞt�T/?�fR�[<�t���C��3k���;��g��[��]�;�
{t��g/���k��Sl�aTl!��~�&F���x׼JޱLq�f�5æ�oӬ�pNd�8�w�Ğ�H��(t��~��I�`=��?�9
��R�zI���7�M����bM\�{��s�J��V��cU��8
���(��O�+G�'m��ڪ�4�,ﴪ^�1�U�q|����ZZ�+�Bn����E�w�!����:�o2/kt�x [��}�x��<�i��q&�L�q4=?8��g�{<٤:��s���\�Hc۪:�Q'x���j�U{@���X�쿮	�6�k|���!���g��Tӳ�wU�b~M���؇���O!���J8�,jY��x-�S$ ��AH�C��<���y�d����-��~�!��w�&�纪A����P�� e������d[��O��}b����5X�g�O��y�9�"��\@/��w	�G���\�`�%9�ca}+5�D�z�
�����S�_�v��M.�b�mǴ�0�8��ě<���j��m<����?��i�3YhUa��M�U,��󷹐�;��ﻫ�"�%�(��<���=�x��e��U��k�S��"߉�����J��>
�"I�_b�Bf%;�;
!{'��`�sś�H�~�dRP[h�s�o�
�/<X]:�������!�)�Sv-+�F��V)O����G'��#�u��p�y�
��f�Ju9�Y�6d�[�'���fd�Z��5��p�'TV�(T�� 6���S�[�C�h��&��{FK���;<C�5�ؽz��b� ��O���:E�����?x֩iLe�Q�㊧wC�)���0���gܷ|"P�o��m���1J�\�g�k�� V�Q.�U���0Ma���M���\�9o2���������ϺY��)&� ��=�;�3P��k����Es\v����/�iS0�1��cG{0�.��&�$�h�2�*�b�B�n�tll��)��MS����"����u�|L��z�$�������"{�u�y����p��p�+FX�[��ůQ6�$��]B|�5e������2S�&��"���'m
��`�	IȆ�G)Y5�Oe+u0N*:�Y�6m�>yD�|�&�J/�[�/���F��*\*tD��ʺ�P+Ұ����f�&`.��A��56�*�4�3)ƕH�3X�����)����z����BH.>.�j�҇���N_,h'0�N�Q�N����zr
,��~��zL��J&uR'�<�.*H�8�n�k�%�w����>��M鷤�fm��(�,����P�i�I�b�^���`�ʯ��a�?T��=���ro���X���<a�������xP�>��Q�.���Sg�f����z-���>1�Uqj��D�<�yz_�R)��J`6ߎ�Q�G&�k'��b���=kD�'�Z�����>Us��DO�T�ѭz�&�sBeV])�AXߓJ����*5ۚ��4�7Z��j||��9�z=7��6$-�~�Z�:<c
�ޙJ\T�
+TT��	�?ܹ�Z��5� �m��E�=}֙���>f��ְ��[�dC�B��=����!,*a�yS�Gj��C���_��(�ע������O�h����8(�S�X��4�L��{~����{<�R�a���6��m��D���Wsj��9��v����
J�1Ja��e�a�p��y;&�i��#��������}L�.���zB��)sam�-O7���
q���{��Ҝ��>ke��n0G/X/�A�$��~���,�
=�̻t;TP)�Ƙ�yd�,�)�F\�o��*�b��Xy�kDɕв]�����W����#J�sv5'U�E��Y�u$���a6�	��(����	1B�����5p�;���w)�����,��)�s���6���-?.���M�j1�k�� ��L�Gx���zĢ���6�A��c�"`���_Pk	�"=n
�a�Wĳ�؃����ま�B��=�*�ֱz��/hj�ո���ڱ+��P���`���l�S�)\~Mxa&�����#��3��_�gl����٥z�x��y������<����p@G ���P;]X��!X?�M�6ޣ����o�OA�.:�Z�t�Y]?La��ம`��^�^�kGeS8�^�/�.!��V��^�nٚ����n�wy�(��'}��M��
z�-��5)��Νo��S��YR���L7,b�!cr>�kU����G���Kb�7Mz�]�-�ѵ���0.�z��������q�nq-O�������o>��*ʿ��Wm�6+�ORK�VIF�a��1�ާ޳�O9�>��= X�%�T{�Woa��.��P�+TJAK�UI�Z3�� @�ZU	A��tA����#����XK��ڸ��1���,��~2�����!R��v����-��������%юD� � ����
$
���My��XIx��5##��ִ�4��+N/�z;Z�{�c!���'�Jr�x��#D�n��xS۶��F�!��8�t� ����g3��,��X��*�.lY�*-6�ViA�Lu�i��]<E�F�-�2A��x�=��O^<|�d>��ݤ¹�Fe�g(�R;�ʽ���9�:���1-�M��F.T�Z}O�K�Q>��*$�s��j�	Â��*�Z����y�MD8ƺM,�1TP��;*5��1p�%ѹ?�
&�Y߳ܒ߷`��+$�Z�פ�K��`=���.&��{x%��~�g�FW��d�^�=�RjLȩw¿3��utd����;�?��@���IJ�U}��|��Q"E��Q%Zx��xJ�Z�s��M�kI$#��ȀL\9�m�4c��l�g�� }��,Y��q����-�!1$
ME�B1NfJ��+T��:*}���տc���b��9i�h�#4c����,�#=?]��-m��P${(��GKepO�Ϝ�*������cve�O���?��s��>ޱ@������rN��U��*���/@�*-���̫��[(8!�QKF��!ì}�!�� ��k�dTJ(���K4�u������UQ�B�O�?��d� ��H�z��|����<Jy%8Mw�)���w��G��@�E8:�R5^
��C,"��k�g:L�%Έ����uD�0�AP6Q�?nh��t�B�a��Gx�����-E��7z�nNd?�����ew��HPou2�4�;X��&��qS��3t���D�2;����`������ϊɹNm�뷮!��fYT�6����-��j�Ty /�,���v�Z������+�@�աLB�,4�'u�o����fD���]Ţ?�3��1��UliU�y��}v�i-d��U��|���U7�����œH�1%ڄBSc�ƞZ������rZf�Q�[�Ȋ7|d�� ��İ���`_V�b�����y�e����+9x
�������������;�xbx�2TRzYޓs�W�Br�y>Y�R�;9��[�I�%ߋ�)�w����ϒ��sT<
��yM׼k-E�]�ރ��r���9]�*M��������KN�㽄H�%Peb��Q�54��2�V�`��޼?"D�2���DkC��yQ��v@Y����_�����o���`dCLNZV�dlM�6�7�8�K�i�QL�)�����U��O�Kx9��+���Uo��m!Q��@�q
̥֓��n�	���G��cwB�C� }���k���6�(�F��4�����& ĜPf� ��ߛ����;�`r���n��`8���R��g-Ɇ"�E�o��1��!.�7�iԜF�'#���7�L�<�Q��ɴ'����ԇ�ҏ���b?&�� �̣$ͧ��I��U+Օ�Dk�t��s@XU����i�2��`-͒b���{��g��m~Rd=��W��V��,�ik�j��m��}�ut�k�6?f������Ţ1�bx�*v�=�ڍ0���^Z���l�y����m���HD"a
�aCs�%�&ulU���5}](b�Vs�$&�5�Tᢵ���-Y��~�oϗ�c�xX{4?:��tC�1ǌ]�tQ�"^NA��RE�1V�xXa�p�i5Y�����"u}�����r-��LWI�&�H2$��!�qQ��S�K�^ءz�ޯϐ���~��Utz}�U�Sed�2c�i&����I�����'�w=w�qrh#׽ޟϧ,$�"�MHW�0�4��O>�����(�7w|�w܋�^�Q�5�7�B�g��Dr�?�Lw�|�*;6��B���nmC��C65�â���D�x(���/cy��)�O�+�F�8B�GL�3K[�fX��}�Hx�8�B@@��ѩ�b����%��C�M1�G#�-�!��.w��}d� ׳3�.0,+~�Ir_�g�U`� ��YRExd�g��u��i٩��89��#<\���#d@Y��,t���^w*�0��w���؇���j��`"����8�SR�LW(!S�0,#��e�fX��B�
�R����t��,A��o>�
��%ڄ\�l)4���ۡޒh<�]��R���7P�a<٭~�^����L�(�P���!����J��9:�34��AL�������
�E ��ڍi|"�P��F��
mbX�
�\2�^#�O~G I��~�?,�h�J fN��������L:�Gyٌy�&0i�xf�r?\�W��{~��i�F�މ/׾kF2T�C�o׉��J�g?k���g-x�R�SHZ���p���9\�PYc��*G�{�0�����=׽p�V��
J�B%� H�L����)���U��ɚ|De�������Sg�����.Lp�r:������%6*�b�a=e�ý�&��G����{#hu?%����L\��a�'�,��l2^	��agK�	ƣ��s��=�15����z��T�vQ��]e+!���p�,�S��Bf>�Z�S����l�O�����Q�d�
M�gA@�Ʃ
3��8�x����u���r�@�O�܊�̶J�8��ӆF{��cN�e�y�P�p����E��N��v��ť�G��
�����o�#T2��h]&-x|^:�60�'�|r��XQNxY�*�>6f�A,�&���V�/���.P�>�ކ�7�(`�8�;WnU��3��� �����}��jmZ�*����R�!�(�!)� ���v�y(,+<;.���3�b���b%},�٢6ƥ�BK�o%�l�j�:�����vSi�a$䏂M���p�L�����U��3�����t���y�������ޡI�)$^����#N���㼸؏R+�n��5_.�-�H.��{�}�1��C)�b�SkXE�JC���^��p��[���r�}Oe�=hd��\'	Qx��۔׃F�СB۵���H�������L�15c����5��
PE�>�ZưU�������������q	
�f�*��5L#�=�F���""9�³:F��n��4.�8AnT�Iz7���s.��e��<�����Uz����5hm�{o��Au=S�9+��
�#�:OP�W9��ڰһ$v/*5�Ե���o�y�yH�(�}}��(����3�~�"|�y�5��[�&�`��\�3.�(�� ���C��.��������E��r��e�r�'���$���2 U �5ĥQ�i��2�h��)����S0�)�%��\�׏e3�8wXh�KK|� p��w��~�S^��O<��N�B&P����B�)PE����Uy�S���d�lĊ2�#�'5XƩ�eq��S�i�$Q<��=*��[pz,�x��]��*^h�Q!Q0u)�R}� �7h�?��3�l�ƠG�H�m~�¥>b����K��Kܧ���-�X�V���)Ҭ'��:r#9NQr���<����)���k.�����#Z����;��VmU �<�X�Q��w�t͏�}��<�8����}1߷X�]���<�k}��D��E�Bʟ)����@���Ƣp-$��s]�H���5�k��a���=Gźd�vD�1�g�[U.O�g
��g^_f������_��,��`Ֆ�ps]�C��S��RG��J%`�8.^���T���T�	�L���S�4}���Y�}Z�Ayx����$$�\@!L;fXD�R/��T�jUdˣJ� M
EhH٥J��U�aL�FP΅% -a�\QV¾��4�D�Uf��]&��T6���J���U��l�=j�z��*�)L��Y�5�A��#'�Ɓ�i�{��w���Iz �����D�U}�"�r�&S�B���t��`Y|ۜG�y����G�Yz+"�W�����`	u!�X'�H.|�?o�#t�L����醈`Mم!�:��P]����9�bm��j�^d�:�b�x��@��|�
4USp
*Mkc�k y���-c�MI�f���6����ų䧋�m�N���ZM5I��y�hC��tڴL9s긴����x�8�T5��V�l�S)e�e���*{�U8���s�dy�
w�kuJ9��ts���7&���Q�bU��
Y��Z�����	���}��^�?�ӽ,V��ӏ���"�C�}ȴ�����sƈ�Ð���w<<�=��I�ץ��(rM(�}?��
!�R�ŒVJ�5����g��q~�^>�[����儊�*��Q������7��ߔ'���x��\��"k��<����P_	����P�~�2����Ln���j���n�o|�Rt]	�`���<X�����$��hX��K
����2�v��N�e�P�Y��d��f�,, ce���j�F�|�q��s=��Q�#�ɓI�P�u�<*[?�YZ�f�ȋS�<^�΀��*�<a�N���=��o�4�}B>'�D;���\��i@U�1�UWTҋ��T�����	�u����sx|���W/"_>�A,V��'3�O��VA*��z�s�{p��VL%8 ����տ�W�����ⴝ�5&d,�X�!�$���U���4�6P�B��/:�JG��f��6��T��R	�ڊ43����<27�9ƛ���7;F{:T\Z�6�Z����o+hh�������u�9��ňEe��V-�=Fr�e�F+U�c]����pJ6�lQ���h�'��El=���w3��Z���z9Ǝab6>c�9��pJ���t�L����9U���33g}�}����\��w�b��y���]�~^瘾B������5ܿF�O�����O����74�;�(	�	)��+)*3Q��+��kBᯢp�����K��v=���u�i�޼����T6*��V�&_5PfUI�z�k/�������%���f�}������<�˿��R�>���j1"B�����^\��.5[��A�a����Vs]�:�[�{��jN|���F2No�N=+��"[��3���/�.eYlQ��wM�Ϡ��I>�RQ,Y�\������ߥ++�RN�J�zg��;����l�<�G�T8����n|Oy澗��{%v����;7nU���t��?�K���F*��#E��!Ɍ��(7�z"���Px*��cd��"9�G�+P���'�����q���>1�w�=�:on���id�4��+�a�r�ϳ:v�����e*�o>���#r(7�{��)������W��3�6�u�i�P+m�`�^덲_[��l�(�X��$���/ #|Ē�u�����lYܦ�x��ed�VO�b!�[&�^q����11?=��+9Hb������i�4���{6ߵ��tG"���c���V�B����Q��ڽhݔ2ܮ{��m
+�<7��J+����7����Ha��iT@�BF���s
� �2������zޣB"�H*��i4��Y*�B0�\
�x7}�dX1{;�J*s�߯��~������yaa�L￿��w,�&�J6ʰ�0E�K���:�)��v`D�F%r�8T�*�'�;�[H2�I��JL�s�e�-S�9�h�{N���PI�atf}��s�O����������n�Z�Feoj���{!Q	���ƈt�F1�q�8���g�|Cr�6@�}cyf��I�^_CA�Ӿ��g�5Q&+��Vu��1(�=hln���KWm�De�<ۗ�k�) ?=;e�^U5����I��u,=��e�4Xn�g�v�J=�&]��#j�};��t��
�ղh�x�s��"��O�@K���K8 >���QlO
' ��OP�&�{O�B�ؔ�B�:2�u<,v2j�
w�7G���e�m��9cu�o��pg��,���.�O޽y�����r���%-�k��!H��޴x㊐�n���V�]������c�&~�"����� a�a�\u�(M�b#���^���=F`K�-�����1��.�I؜'�X �LY�VH�S��WI@�FCa6�DH�U�(+M��Tqk ����sF��CNk%�7�"�Z� ;V��X�o�{�Yr��*=�� S�y?W�)���/#���H�6=c!	ě�@�\��C�Ë3^��+ξ2|բ~��yo�U��+�ﻟ��:O	��n��Êp���U�|��\�s�=��R�*k+Lϼb��^���F����~?=ݧQ}c�5i�.s��&���\��=?��L����߮=���5TB���56�?�O������޼�$�{�x���{+�\b�1BV�gcY��������}X�q�P��߼�V��9�=*�	Z��M��ۺ����E&�5õ�&D=�x�����	^���߁14��A���iB�V�FNL�5�S�"{�r]��`���Ҭ������
`���3I~�S����z������&��Q�;�x�ixdGp�Qz2@7�wV�"[��k;{?Sv�Q֡�YF�m%�"F��I�yiao,�O�0�MR�ֶ׀Ǒ5f�X��őes(�rq¶3/ �@��֚�Sl�����I��X�(s�wh_��[qa�a�S����~�<��
��G����N�a���_��D���GK����<}�֨.��n���t���pE)o��V�G��z`+D��5߿w7�?.�l��������//�͢��
C�f�T�+�VA���DE��oZ�z��W�}⬞�ؐ�L�@kZK:�Dl�ҷ���@Z�{�¹??9����G~�S`QX���5��ȹ/�T=f����5���+��!�s�cx��$�UW
�#Ų���5��xZ*�<�
��5��N��b0yA<���pm{�!�/c��p{�J���N�����x�=���wEATZ�4�TH~�k����W�Kg�z��g[�Xs���ء�k��1�B|,���<O��2i*Af���$\���b�T��,��0������u����.»���;�G(�k�rL��#[T.�h��4�2�0-YO�X�
f�ã'OIX#���� רv�n
�^��E���D�OS\�,��{x|*&(�m_����� ��0��R)U�k�b#��QZ��H�j=�1P�Y���F9^��}�6)6W`���������B�z00�&��#>�3إF�(�0O�ۥ)�e��Uc�`��������W�eX��'l�.NkX�%B!�b\x.f���K��c!g��W��R�����yU_-��̻S������Kuʰ
�`�+O��P��4�L��W��Rɵ%z"����t>K��� ܗ������NE
��ܼ�V`(P�&GA�E��0'�J�~GE� �;z�
��I)X����̚1G�?ދǤ�E�ǹ�\��~��B��W�1��Bz7<֯���c��5|�Y�Q.�;�c�<k_�<��r������'��]+��;�z��|]����/}�Tʪ���?�9g��DY֧�����8�_��t���w�P�$}���(j�!	�~�W���C��U����Œ���W�0`�(�$ī�C������#����8L���Td��6(�/4�jK�~�>y�"li p#� 	
�j|�zLSz�f�2���i�k�E�à���.�9EH��"x�,�@�G�IC��X��҂ڭ�$�R�dOVsa�os�ua7�n��G�m��t����2t�'�(^��K(H����)��f�},Ѧ7���T�N~򞦐�(�������E�ǰeFh׶Hՙ���ݦ��e�(s�b�m\
u脔�kR=ׅ�S�$���Yt4��.�T핳њ40�ƒ��ks}���l���qhTE��4�nօ��R?����9>�7i����4Tҩ�
<7j|�	�Щ �<���
��]icpn=>�CA�<����4��5g���Z�:�tμ�8��o���I�y�Q >�pI���xLJ�y�ǅ���I���1T��-��hۄ�%Z��(�(6��uI��q�'n$T�wש�
�/�0 ��(;?�o�.�Ͱwu��SJ��m�lg\��{ծz�b���~_Y��������9�~��@��R�����I_JZ�rs�y�0Jz��"�T����\��G?�q���IʅJ�������tO�T���:Wqk�yM���w}�X�Qi�6�b�۵�pB�#M���$��8����'����}xLA��BU)��҃�����E|���[��7��3�^/�n-y�KE�Ϙ��~��S��G�h����42Be|Vz�y�(��0"2U9�����e�ւ!+wz�����/�m�.�k�QR��8瘊x�VI��Q~�@���N���3�ބ�p8E>`��Y�س�Pw�ǌ�BQ%Y��	�����=9"����!�$�*2�L�
^�(5O�pܬ3ǽ<%ul��Sx���(q��,��1a%�]���x��̓�2}�5���͘8v:a�m��xSޒ������97z����+Lس�R�";�X���"d����ƼRt��TD옣]j�e���:��SP��J�T(�V���_-塝��0*��xn-ǲ%pt����wl-���gS��
����[~PI�,����e�n�ef��*־�֠�{���s�{]�¢3o������-���y�n�3��뮝����^o���vc�����a�����7F��ǹM^\��仮����/����@��E�Gi�UJY�-��X0g�b����V�xͬנ��u����e����T��=����9�iz�*������u^�ZrSm��z
��S��빼��H�٣ ����A��#jk�C&������z��/��H�3ͭ[�V {/1���q���F
�bh�R�:��\�b�W����Ji����]-���<d\�?������m�e+#�3Ul����z���W#��G$��ݡ{���t�#�0��,�kal���^p$�d)���ٕ��Lנ�+^��$��� /��/��x����M�p%]^���G�_�pE��,�k�ҵ�s��Cȥ�DD܉�v	�h8e,ak���G� ��Y[����o��+B��F��ե>�ǋ���y"<]�Q
 �M�m�ƚ��t\��;�T�)HaW���*ќ���;��Rj�'Y��me�uJ�Qcl���R,]x�f�������^�K�Hv9C��G����(}O�Z!� �\˔$r�+<n�H��1��xm>�B�k�[��Ax��y[m�!I6���R�6�K���W�Y�o��{�[���1^h��?��	�{�Y�m)��@��W�Q��c�:���*�Ķ\[��ʳ�z�8`�Z�K���ؙ
!J'y�^��>܇-P�vۇQN��
��TBWz5�R5�|��_�Eݓ�s�X�T��8����s�=a�T���{��+s��-��\��C���^A!�'����lm�:�D��n�;��^�z�i��%��H��zGț�I��5�+*m�ƔUs��/6��֧�g��������"��EW�~� �Q��)I����Ӑdf(�?��#z���1�?�_�h�bN�Cwl��Ş�tT���!����&5zQF�(Uکb��&�]XQB�}�\`P��.R�x�t�y�3�,
B�J�g"ҳ'x�x��x�y�7��nn��� l�F�'l�>GZ�c���h������R�hK���OBB�d��d<B�w�蚦���%	66� �ar1�U
O�D��g<���_q�Q�^�n�N��٘^g��������2TC�F�J�u���M�:;��)��3�;4W��H�:倶�4��?�`�ć�;��a�UМ��YöK�?tv��PKAⶱ�<�
�6�2c��Z�Qb�OkZ��O�-��[�ȯ��X�^7�^e��"� |z	&�{_�{��Y��^��U�C�L��Z:�'��u0;0Nd�����ވ'�U|��o�K�J�j�c=���.A-4�q���\�G8��V)��X�5����;;0�z�`��7��;��>��{׊���rХ<h�V'�L�1	�~B��XKE%a#� �B�0|�z����s��0F���~L�Q��(�tn16��*�8�^����[E	&	?(M���cRFq�-�����hFK����h32H'`,�����/�����y4h���s�<��s�F��\�i�~3��f�-ܡ��b֤a�l�2�]���[�C2�Sh�>oAlLh�?Q6�e(+T�Έ�,�����N�
sDmP��Ώ�,S��Ԉ�-�����ϟM�V�� ��4~����}�[�YR��c^2SU�G�,���o�����ӿ�3��
^�fS�lz��OC2����E��r6|6u6c_A

���:�L���8�7mu�ψ1�lٖ�d/T�a�]��RP�+�e>�yyn�3iU:��F��V	����bܰ�=p�.WT����EF3y�>i"�����M�gyv?S0�Ąy��E��r�����S�Z,W�G�*�������ʲ�^�Y}�T�N�FbK��SZ����f�:+ܜ�x ��#y��w��y
�\m�#{����ś�6��HXBUV!i��q���pMIvfR	�3L=
���mH21,�V���~�g��F�Xf^5^6�z~�%[n���l�祒
�u��˘#^�VJu	6 Lc<�I�UΏ�,#���;-�r�������M���ʕ�$����zu0���T��*u5���o�:����p#�iJE�G��v!�x�V��F�vy��01�ˋ���|\M����3��/����^(���o�[���zo���%��E��5�%�P=7��4*�7��	/Z�q�KWRH૊(�I(<t�l ���&���o�L����Ҙ���[#m`k���@��(��b����`%7�"� �7�y��� Y��Y��B�@���1��s��<�	~ı��=?%l��d^6x����6k�( �F�@�PG��(�?!=xs�������U�M㔌��T�yt�~�V���y��7�_ct�|:f��,]�&�ֻ��s[T���C�;��E��-��F))=�712��s/oe�9w�}l4l���m
��X��������M���{�S�`���(�|�m`i��@X�~Kx_-��`y�����llǜzݽ�,�����|&-��<IN�_��T�B6�V������&ש1K��"zj�J9gc�p=N�������P��9Pa�[Y���EJW%�����t�˸�W�֏��f�{������IWġ{���N}C�3��B��o�.0��[29�C �g���ȵ���\A��
+�Z���
X��/��ZEIora)��G���ʹ�+{A�]��^���\IH�>|��	�ST\*��Z��^.�L8T�����3���� ����2�zmc1�y^��)D[<ËtQ'��w>����do�r-�2PY`{��^2�Pϵ�^[�	�l�P�GU�j��-�S�4�2+�l1.{2>-�Xqu�n��>�m�JHQ��q�ԇi��X�S�Y�f�q�R���Bi�,��?&������(��)x��R۳��y��roݺM�l�SxQ(w����šd5�G�l�c��}���M!1�t��� �cr���a��s�2�?�����_�Ge\O�)`0hwf�E����㴩���O:�py�vO��9�6W�L�	mxt/�4�4������UA����k�0&d^B*"����ެx�Pg�F�'}w_(���Ou���.}E����g���q6�����o*S�hD��
��>�ԇ_��9,�sܰ���u�Jh�	�Z;��y�ʻ2�����r�g��"DC<
�!�8E!
e=�"���j
nh���l�7��-`{�]��ʆ����E�����S�i�+8{�Q=!�w� ?�Y�W��聣�3 J��W���}"Ό�>���q)��3��j/;�>�0��a![���������N�(C��ӧ�F�*F���o?�FQ�ݸ�T4��B��i��x���zB���F�r=Cl9pE$�T�
MZ����kv�l@���z<=E����������[�{5Vme�!I�B�b>o�[�E�+M��i�k��WTS��\��k(��@x����_�l�Y<]���-z�M����%a��*B=��A�p�������q~�Lh���k�Qs��'�%�f;�-�)�u(tۚ����	���7��L�Ob��kHxB
��j4�m� d���]�������_���M��l��s�Lui��牽S�zcg!R���� � �C�op��K�B��8�q�	8�����l֝˃;��YX��v�A�Y��Cb��9���m���<1#}b�g��S6�p�9�[bLa�[�Y>n��D����%L���S`�.�Z o��m(B=B������{��,�x}��������B��%;>���	\Qр�Q,��`�Se�u΀��aX�e�Mᕄ�5���2���%�:��k�@��>3>!�r��F؅��eFg��:)��= 
o qqn��Q�/�O��E�g�C��B�Q@�E&����-� F�gn36Q����6��eJ�Փ5~� lA
V�/��;����)H�C��wf���X��h�-_��ř�@���qNUh�k1�5Q1��y
�/P Y� E�UP�j��2|�±ۂ
Ta�Z�C���6�����@��A��T�F�R�6��&�C��̳���J7uJ��!�E�+�/dj�M�U$�$���,T�f�¤���)Y�J.Uى������6^��Jy2��yF�@�#(��vtp�bLJ�90�O>�)�/�r ��,�w1��?�8�h�������> I�>���Hس��N�o�#�Sc��x0>')�6-�x�a ��BY�"�Aq�~���Y�]\���1;���逡'LJ�Zu�癀7G���_�z�T�T��8B^QE��s� oR�*,�Y�k���`��&�  �0�� M�]��[��oQ���*�GC^�򧬁���I����~��{J�?������h��SF�(�a�L��P��]�99�^?9��r}���%�����[�E�
����#,�@��ne��bR�k�EAbC[�x-)�ς�#v�/RBK��z�^abl�F��9���_��=w^^��YA�g���{�:W�c<�������׾���1T~a���
�F�@8|S$�O�����D���/��+a�SH��F�3�%�Jʠ�Y��bϩ��yx��� �kI<Ǥux\������/����s���|�	hHCߣSH�"���U��=�MݾEwvW���G�L�����[B�hqC<��G���x���R���2����S/�e��>�s_=b�$�^��imN��
�m�6T!�Ӱ�g�<��$*��UٹWhv]��O��[�S� ��i�˯�n�����D*d�zI,I�B�O�>�^�a��O>�%�%���р�Y*�Q��=,���B=M��e��/A2S	*3,d-���iB�(����ώ�f%)����[��fe��	.�ÖKc(�c�IG�lns�k@�w>����/�?��T�17�ߓȼ���(�
b���}����:���R����g�I���X�æ��IQ��s����_06�H�G�rn��0U��ʄd���ʾ��}��ʻ�����`New���C���n�>|x��`����"��9h\:�l��L~�z�t��`�x�;MQ4{����z�:���}v��ેip�F��@1�ABΡ9�#(�Qư1�	����	qO_��'��'x�?EرE�T�}�Vs+�����`�n�>�(I��(�fɪ-���?*C�wsٟ��Ep�^�5CS��)B�����ڎ�NT���w���}%�s���և��.Me!u��׊��z�ِ�Y)�T���/��������f��f�Ǜ��K\*�0^kbU�Y�,<�_=��D�3��ol.�ľO	���E�����FS�q.|^	Y��k��8OM��1c���Nv[�	�@�ޮ�[3�����0r>�z�}�2���6��Ŏ�������lmgIf;Ƭ��b�.�\F����&��]���^�n䌰�-ǈv�z��-��kU��΀�hJ����F�_�mB���EJ z!���=���3�[Ϻ6HvO��v8���zyX����R��:��2�%- �N��� �U�Ps���*C끊G�/�w�?��1���!�ڍ��H�����s�x�F5��MJ����IJ���0F-�Q�d�KЭQ�eEx4�|�8�,� I��%<5�E��M�]��n%�مmQުd�K@�&ǯC6��s�#u�o��^�#�j�� ��������}�u��ט'�����w�1��qc��D<;��y\�|@й�0Y�A�<��3�z2L��{(鯿y8{H3p����m������ ��6F��1<�I➭a��i���q�5d�jW0���s��޸G��3mB���X��	�>��W��ΧP���:�'#NW��
�}���[;�
�[���^�,V�C�%Ji�s��J�6���'c���.�$Ĥ����u�1
G���dB�^'�i��g)Ӧ����|%���t�
$1��b��б�1}�|{�kޟ�J䠱E�[��}O��W���f.����.ϣ��uF��P	��WS:-��cZ �n�/�o�5�������&;��x������b��9ú��j��<B<�k�I0��6vh���,�*��X=E6���5ڶ�lP DH/V>rM��<S�C��ן�>q5$�s��B�2X'�s7����biO��(*�H��������
}������1.Wp?rÔ��v����D�[�Z�C�����d�}�<�m��;����k$�`�3܈��\&MyX �J՗�YRP��c�r�8�����EY�P�l��U�U�+�mZFq+'�ގ �,�H?�Y͑��I�V�����H���Ĕ=�󬗼J~� ��c��(�Kzd��U;��߻��׉o�kC��c��l2o�u�z���D)���<�8��~4xz�8o�Ll��A����#P�q��1�]Պ6�e�sKd��Y�/R�u�rľ�(ĊYN��LMlC�z���÷��#|]�շ���� �N6Ա-�r[3� �D�������H�u�9���^ӱ|�!9=���Ɠ�GV�BŋO(ȴ	�G�*����l&�,P_�;�TG�&��ӋL�'������b��Ա�R���K��gP�a��̏���M�'�{Szg1�(¶l/Ɩ�{��}BNA���̇�w>���� r^�ߧ��\P�?��f�ӕ����z�=��װ��q�hXb���G �*����ԊlE��7|�`5V���c�mjk���ձq�H�k�	G
�
��
��J,��&}Vyj;�k�b��9/�:��4KE`�i�?lKjϸ�E�H9���1��9���N���-�Mv6J{�{6~��ʓ d�H�=���1H0��]۲IB��}a�ȶ�t-�m�3 Ӊ�U�.�!�����e���Xґq?c��[��](Յ�7o��^��C�ޡE�m��x�0zMז`�JV*��Ґ�[0P�e1z61~��w�����G����@e�%����#�?����E�$wefd��KHw�/���i���#���+<��?l�qRe��I���!��k�<�?C�1��wx�h��^-�������Q�i�GE��rel�n��uH� �fj�NO�k��ym�r��!�����j�W�X���� ��nu�Q��,��[<�~��E����h���������>�4䛖H/-��T�F|�D#��&̼�>���$�eŘT�נ��A6Xˍ���
 ���Ha��k��I��{�B��L_�TJ��a�<P�1B.:���B[]}�;���yn�/�v|Q��n�[���r��~Y�@�C�����+�T���I��C :������kg���daʒ/ �U�
��Y���6�{LOp�)�h#Z�uY)]���G����|!�7��ֻ���Iџ�$��l�
,G�����?=�d���Θ�>.�q�@|A�W�b�d�oA��*\߂YIJŶd�&#�z+|_���M�C��kƂI���0�F2�w]	��Do�oÀ}c��)�c�Mr���g1��=��������f-����w�� 3J(��v�e`�E @翼�����W��ǔ�����;[�����
���7x�_�}�'����	�5g�&e/l�������������7�a,X�F�E�`�<�U�))�0=R
�.J�)�xjv���J�㞓6�����N`�@����L��]�s��w�׸�� #T%dis���a(L:ct���}��6�ېzފ�}�K����F��,Vs�<��~ܰ����A����Qb�z��I�o����W	ė	�W}�~~�?gs�Z��
Q���akF�*s� �G \g���_|^mfVW�M׋�'���;�W�Dm���
C�a6��^�N�� U��z_���1����v���I%����E���s���^b��}�L�en�������r8U�Xb���X��sW����oc� g����H	lO�cc�� �� c��|
��Ē?��ڳX�����|�K��n 
b�ؗ�i�5s�<w��������-�a��46hA�5���bƯ�.�b�t�"U��ԓ���Y��{*~D �\���Ҿs�2U�T�3�*.خ�{�V�9����!��x�[/���oۛ����16*�K�
3�n�E�n�u.��,y�MQ1��pb[vo�G	6�q2�@�O���>��2J)��������`H�q�d�.�`��Y&i�
����.������4l���8�OP� ��U���cׁ/'Q�k����c2�z��m>�s���ۙ��P��oY�N����'��M^�>����^��qO�:���1��E�M~_�N8�����Ӎ�0@��g���jQ��@һ#t�ek�^�jC�Gx�zŦ�L1��|�%&s�v*J0��7�;	:6�!���O6͂�<�=F뾅�7��;%Xa޹���D_��w6|?����-�%~�k�؎;�2ڝ�Aog�Q�I]����3LC-|������NM8Z���J3e��^�`��V�
����U�Qv~��z�T��gM�P�/b����"�cx-?o��;��o8~�z�~oC ��[w���*J�5s�W����5�0}��~���-���$d���^�:�Bӫ�����:���ם��Raym�����jL��q"`�H�!Pzjךp���\�qV*1%��1+]W��c��m�I����[���{�Rz����&��\�]��9s6��R�1)]�m8��P���Y�/�|֞Kx���!y[��,�ޯ��Ŀ&QzvS�M�P����#��drs�Fi 5��w��
	.�'�>�zn�{y�Ĕ����(�]���PY'ַB�����/��2P�P5���?�j>B����u%,��A��%�Nq��@d9���0�'�(�c�ZL],�Cؑ[a� �k�W�@�dŢ��e�5^B��!i~c�%�����ٌ��&P��O�VN��?��Y���y�sh���Ga�.f ͺf�I�6�@�@F�|qu1 68�������x��4<B���hg�o��d1���˱$Q��݇�Ae��{R���ӈ �8��b������(�����
?��L*?S,� ��O��r�:�"y��Γz�ר'�+u"s]�9��#5st�y��g|���1�ӫ����a��;fN��[��Bz��\�-�Jӟ���U����8e���������^3��
v4�d���aّ���E"a��}�PԆm`r�@$�tī��tM��j��Y p�Q�v}�5�k���:u�@�v}7�]/t��:<�㱥O5%��o;BHӷ�߇(9�zV�� �_ۢD��	�#�1�e��$,T˜�G8.S���0���x��Y��
��������E�7���@�s�+�I\[�^�i>�2�3� ���#b�[x�_�y�37�:��-r��$핀M�㽄�i���՛��1�O���Mbu�8���(�)��v�9���g�q'x�?b���)ͬ��87X}�g�'�����1����=ݢ8�8y�����q�JWG��WExl��������P]�X-��/2�3��e�R�)���y���$�q�ý4S�f��&GOv@��_��_�����E}� =���K$Ȱ ���+S7L#�|�UM_H���"��P�C����xS��%v��$T:
��V(j��]����T^�(x�E�Y�w:(H��Sq�ߎ�ד��)��İG�����OQ�]d-�Q�a�������˿sF��ǿU"*:�[P�ݱ��ţB5	��	�ߺy�h��6Ep�)ΐ+f�rcЖ$�ڗ=j��kc�r�<���3b��t	
4���Z�?���W�O{�R��)�^�^�E�h,�zztG��:q�5�i�Be�N���lg�:�2ZѶz`cx>�K�0�j�,ϸ�7"��\/������;bz������4�Ls@��	Q�(b�ԩ*���D�1�(�~���Y�O�[��h<&f�2����Ja΢��o/��߁�yb��M[ y����W�~M���m��ɟ�	�:K�Kx����6���+�@����C���'���AA�<�cll��)�a��3N��uN�y���]'����_�|0�=������(�g�}������Į(@�Zm]��1��矱/�J��,�YƐ��.��������/w�}�e�`R]�j߽���Nբ���-^]y��켋�ơ�2�P�,�C�ڛXsWq������]���pQ<��w�0|�����=�jX���W���`g���[�Q�������/��� ��T|��y���D�Ae�B����K��j����G/����4=&Sjz�	�%�ܹУ�8�7���$Me�}���W.}�ҟ��(���axm�c�}a�\��V)p�yX	����k���
E+��k+��X��oN^�����f�LR���i���8�mn\K�]�=��N�G�y��u�����F���z�\���G�5gQ��m�䧜�؛\��T�A$ʀ�&c[����Y�i5���\)hTE8G��ʗ-��:d��A~�57Q]yj�����鏌���[�m�س��-�Zv�����1p٨|�(Je��V�\�%�Q�'@������Ijk.�I7Y�~c�2� 
/j�sc�l�s��}�6M��]z�1WWy�?z���o�
�8��t;[��4�C�^'�}oŊ�^ø�J�UfƬAz�
q��3�I-\���p�r�^d�u6���:A!��Ht ��!'�@"1���Z@1����n-�m�6���-�/��%i�L���?�x�2�a�X�pӐjF����\x��޳����2x���m�Ք;��WFW�J1vN..N_z�4;�=;5��H���x��h�l3,��
�Ma҇E���9"������.��~�q���)��������`�P�g�B����6q��Z��Pҫ3VdU-=9=D�N����8��&X[�^��{n����}�}�����\�g���^�����U����߾��WH}}x��/�����9�!��&3׏��*�Miɤ7��K�%PK�
꘣1 5r�`%BPe���ƻ�Bai^�R�Y:�73��2��^x�xTE���[J�9n!D	�&��5\%���V����z\A��N�1��b�"���$VUq}���l���G��jI�@&y^�q.l�� �U���Ek�l`FY��3���t��Ƨ9�x3ǐ���~�W�Rȓ��+\�j���&��W`�N�Q�@������cX�h�r���ާ��*]���7ȹ[�5Y�N�W���7$��\�vy���w���3�"�p�q����㵏�6&��z����������C�l�B�p3|B����q�����J(q$���E�7H�8~�<SC�꤂��b����(M�������2�u���1|�i�f(/Y�f��) �ح�#��ֈ�>�o�ݯ�0�7ߡ���1։�<u��=��+���<�89�g�>�u�����1>N�x�
��7�H�_��:���J�E��{�*��U��U����c_& ���s��㽗�W�7�mxl�4�e3,hw%�ևK�X<�L�������F����t6�~/�T��0�3L)���Y����h�����������C�A����k-�F���Ǜ;OI�勵G����<z��m�uv����N]Y�ƹ��zP��.x-��kȨ0��9�
��xˤ@8^��7(iCN�VuC9��?ϹA����J�6T�_��!䋾�׏�X;��=�C/��SY*���rc�G�wjR�p_:?lv�V��]�{�$�J
f������1�$�n3�1<�ʅ�$����I�s��w�e�F���c��~�!�T��#s�t/!�p��k�n�s����Sٕ�<|I�����%�~�����[W/�%�LIa���{��_�$Ů/�0���Z���8ve�W�Gn	�G���g5��|F��*�e�c��Q����i{�w�56,&Nډm�w�����.�]��S}H��(�) �~��4�x�&�[��"�(b�Z����>�4���h��s��i�fʚ�@��(�_~:�����Χ�lP%h�������/~�1E��ȃ�G}��B�
��Pؠ�����yas�c�U֕�9�މg���/��xs�;���%�LFyGH����9, _6�Q��eu���x�v̊���S4J(^E^�;QLas����S��T�	�y�(B�i,�"L��̩����U`*p��k{���C֫�����<������f���wξB�����?�S}�ql�jZ��VV�����kO��!BXƨ��y��I��9��P B�B��|���\��8��,حU�w�d�:���1�\Xҵ2c�j�3jTf]j�bkI�7bb(�2L-S��Jp��x<V��E�!δku��[����Ÿ���,꼈�3��T	�q:�(Q�xt��0�E�sx�GXuv?G������r"%�XN$�-I�%���v	����Ͼ|�i��j0��dS��%� �\'��|�C�Pr�a�Z�s%�΍+�/{��	͆K_"^wc.��������������(B*׮�`��J"�C��(�K� C�\�1=�
z
�R=
̣G�x�0���d�Z����(2�/����yF�H�s+�j�S7���#�X����`���۝+ޅ�s���/~�__���~�)�A�Y�jr��w?�����]'VH�5J�1��m,`$LVsc!��[�y+����,�=2)~�[t����Ӈ�"�c0��}��s�C���[��8�L�����]�~��p��g�����sF��x<�x61�w�;����y>�
Lf�M�/��=%"0i��=�MTs.�kZE	��_���1W��\������a��=ӷ��/S���W���W��u�1M�6ɿa;����q>��Oc�c�aD����.N<��S�L�ɠYKaJ�qMx̝;�G�j>�P�S�t���@�vG��冪����	�v(�<^7Շd�z_�g믱����@c��|n7	H�����q�|���,�	:5xL������Ͷ�[
�)�S���xHs��y��<��H���lf�N}Pa�I�VVhd,c%���f�7�侍���8����Y�t
�q���7�!��2ʆ�9k�c>�ٹ<�	�97Oww�g02�Ȭ�x���!~��ϨڂB�w���>
ƽ�����p�>��;�!$�hޣsFl�>����ʛAp�"��o��g��P����|���vM�+�PxwV}��CY���
�62g��Z��&K���Q���\�!�,Rt%���_b�f(���]��?(���9�*�W������lm��g�-<.�Q��n\�.u�dT<[��[�y+���|̂�bQ+;��8���>����2%3lq^�|�ǝw��c^�idCG!�﷯ �q5��W聈�Й'�B��ł�w��%��0A�f��5��G�m�}�w��$���9�^(�7����{���y�W=}�C��u�w��2�˺=��o{:�k�}>;����@��2�͸l�P��q�E���H��0�,i���/�T� ��<�*�G����H%P�]�][	u� ���ڡs�yr�*u��F����=4��ul�N�?}��eF_9�w[w2B��� �Qrd�V}�-�&�G�����)j=	�qO��8�fi�SG���k�\�a9O�[RL<�$w�������O���MnqHVQ��o\\�y(��
[yN��Җl��7���D,�j7��&�x�pw����퉮}P����Q>}Bn��w�|��rp�g�n���G���?�jpx�ك5�#	< 3�������)�R�r{r����:	�[���k�(`��QԄ<"}(d�%)%�l�K�:a�qb��2d��8����K��	ٞ<7_��O���5c��43g��-sx�(�)R&�\w1��~����/~��+ز�8�
W1h ���Z�N��q�|i����!�>���%K#௾���ш����y+��EN���>����x�2�C���j�sV ��}߳���	��:��,Q,�9�+�eq�X՞+�xU���w2��M}���x\%>�4-ŧ@3���כ�{Il[��I���.��{\U�y��YQ�x1���:��}��F����<6����<D�d���y4�ϢՎ�Uz���q�K�m� �����au�6����`�����h�q3̭�_�+=0�	��}C�p�53;Ԃ�#��;�3hC�平�c�el�����1�b&�^��HA�ݚ��*�jR�g:mk�i�"�'L��lTK���2tV��#�7��vF�ts?��2d��9���6��ݑ�Gk����f\I\EA}p{�z�0d������/eHR�l�j�+҈an�X-:���u&cw�rpW��#��|�E�����{�Z��1��=�Ўkxk<eu����Ai[� �#�g��C�@��0\�ɿ���z��W�7n��7��ކQ����1�vQd�1��j�]3ƙ�����ئ�͂� Z�&��5���Ø���2%�VW(l>����H��N�C�=�����ƣo�Un��N�����-��\��&��
^��w���zw���ߧ���W?���5kw(��|y��R�^GV�MExȢ.ɗ���Q%�:�C��[���c��颊��|�Fj���H1_<�C���C>�~���0�]%�:iíy�<�����X�c�=�T�%��9r|���N����^�N�����#���9�C~'�yX�u��z����z�����0�?r^וk4��׊�د�f����<�^�����WO"�}r���R��F�O{���% ��/֪3��+�iVo��B�I�7f�y�T[˒�k 9���%P�Am���J�?+M��(�͛,o]�Vj�.~��� �e�`)�Y����:=B������io{#�@�{�$�� Q�
�E��Iαc��_�N�E������ܸ �i88!�}/�*4�xF����u�@y>������M+9��|/2��ٽ�/_=��8�ۍ���x�҃�W�$N�ty����(�;e�N<W�r�o��9Ò%��e������	o�fQ���)�yL�����Q�����Ms1�����ᕙO�芅���gɿ6�{h�I�y4�"��d�	��m� h����`���p�X�:�9��[�.�b�1Ɗ�|����2K>�U�Q�ݺ�^���7���zۢ����e����[Q�*@^�w�Ӈ��{��@x�Ӿ-���ۭ��2����׎��
��{}"KZ��>,�Ab'9�B�c����\�s$�,^`����"4w�I:��wS���E�J�06�d�@d!�d2���������#g��w�3�HO������W�a��F��M���~���t>�/��\饫+���B�y����*Mk�ifAe���̹���� ;�#��2.��"5�f�͂�vkP�ʺ<}�.���<5�;M��wμ�j�-w�z���V�Q��<�2�L!D��O)��%ӷ����ʃ�	���}l�B�?�w|N�n��K$v/Ppz����:$'�e3�A|�@�P�����J�)p��ߠ� �d��c3�-�>�����k�@V���PxW�O,^�F�^��3?o6�A����� {����c��m�E�-p߳��W�]�q��;�#���l��������-���9fl,.>ʽ�=[b͖�K5%���F������;��p]�Kf^gH���ݠI��R!��%ȳ���e~|���<���=�B�xݤ`1~�dn���?���� f�\]�!��[�P�v�u�i:f=�C�V��K6��¦:A��ʗ9��#�<���*%w��y3O�*�5B<B��;wO+�^��>������*��)nJ.U�s�xF�Dh�L�0�K��xt�Ƣ�2'!/�p�8{O�0�<u^�Q�^�8Sʰ��K4
5
>��4�,�B7����73�o�,�úg$"Ј1vr��<��g��y�A�'k4�(2�Η�#I��^��K;�����x�M���w߫.�����ԣlUf��7�f�����>�xb��>��gh�y�X�[�^���������*���+��ɽ�8K��ϕg���Sá;��V�(��6l���1����Z�*N[�������� 4��T��.(�y�[��>d�/K��c�潫X2=��
�X�!-sr�ql��6�4��`�?5A��1N�/�%޷KՔ5�?��.���Sd��aQ�y��
�l�۷o�\��Y�?��S<�;�W�12����X�σ���,tO	��`)������{�J)�=rFLz�����H�9�c���B�/���!��!�f��]5��{�6͸й��7�>�ǿ|���?�_���������ߧX;���2���#ތ#=�B#�ۤK|����������T��k�&H�q��C릅#�WϷ�oo��(�.F�Z�[x��>e6�˼��GH�#�r�C�!�D$�ЇUC4�+�(�a��t��R�G�W��a���7:r�|��(h��:�>s�*FcK~�k�s��%����#�B��ä�����n�U�+G�}��c4�#u�hz
cK�1h�?�̓�x�y�B�l>��D�b�B7���K&��U6;�u�v�Z1�2<�bX�P�q�!�YWiy�爁��<���۬[���Q�3���~3a��ɐ�K)�?�%��!�3��<<��(���W�NA,��. ����7f
6�� ���oY�&���ݨ �*�E���m(��e+�ܮ6J��/�n� �f����s�u�e �9�2a爡�C>��bZ)����9m5%�t�l.�:��o�ާ�����`~��'��S)�G�4�/���Hx���`,ЮG|KD�{�bח�j� ����_�U~ ����`�
0k$�?��9=��}N����;x�ݷ��c���m�3\GW�������z�g�����71��G�G#�����NS3���Rޮ��y?oSZY�4Fx�{��y����y��XS��5�P��\+�0��~,PQ���������{O}.
��`����TT�a�&����(��<{߫�c��� �_
N_>���w��CL��x6���䳼����c��P����+��J0s���m�)�L���5D&p���*�Xj��6�g�����_�H�J�ӫ֭�R^�%�P��7&�W��)d�P�O9^�M�z�A}�3�S2bM��az��u�`n���l�$�C�g�> y��A�"l��G��کA�P,��P�D�Y�5KggGaj�޹}F���+���G`w>\�5O�eb��b��� �k�ݾE����Lb�p-��j_�:��2�|K�EW�+̓BdzD�n� ^H�s�;/7�Vj@�3���%���7����sܧ����;�'��d��N��(�}���E�J|*YLY$&�	�/H/Ӹm�M�g��p�)�F-�Fj�ƃ{�'T�Y���l.۪靫T�!vH	��Pb TU"+�l�߹9��?����?F�_/"�k�� ;6�������)�.c��� D!l�1�YoM8�-Eh��o�F_�e�s	��]�ۂ��+q�)�3�v��H�{?"
1��zV
�������\���3M��B�)�1��v�n����a�x�`oϭ�J�A�N��`sm�0
7��뇾� �vLt_�^d,L���@[?g�5�y��W�y�x�}%j��(S纒�16���Q�%��)���N�^�b۶a�,c��ޞzN[@c֝5]�����8�rS�ܺ�^1 eIβ��r��doN,z��{˺�^k��>,C�Dv��o�b��_�@�:�BLY5�{�4��z�
w�����ȍ��gh)���*�X�)�8v/Ă�@�Ma,��8���z��������=J�s���7g����F�hb�M�<�yr�v^P���j/Pρ4��+�2�lI��Vf�<�M�9��[ۧg�TZk]%P�׉Ѿ��:15=��cbm���!��ಽ�X��(+�C eXXk�f�ܯ���Q� C�Ro�"�%�,�KU3J��b<f!���iW�}.Ͽ���W�:D��ą$!~���
1�9�qݳ���M<?_~�/� �y⮇�3�;Z���CKS7���Jج����"^!�d��Eo��(B=A^�,�s���Ǐ�0`{�ӟ���}�,#���8a��~K�Ok1JO"��[������(��aq&(�j��&��[,лa�Y��x��n���P�s@`p���F;B�����aZ=��I�6bG땘Xb�_e�%�j��b?�]x�/��C^��E�ǩVt}ġ#}����?��ގm��K!?������eܨll���!>C��\A��ޡ�d�����2uNlg�'��r3&(�F�RE�D��[P��æέ1�D%��H�P�{��t��"���֗P��Y�_%���k��}�ɔ�D�y�*��������ޏK��D�[�E[�,�J��-sd\���7HkH"
^<J��#7�iod)3�9�!z>�Ȳc�x�>'��D8�����%��Lӛ��ßf�0�sO�}�%yyk��$���x��C4���.�@�*�0㐣(�]�ܳ����jn�wj^s3�X��t������KV*a��'_|��y0x��?����T�Y<�;4�6�d�^�-ldǒ�&�hR�
�~��(r�Q�T��\��\@�b��r��@��K���
6����|��^ j�N�z�g�I�[x`�JSg��q���*��>���xz�4&���ƾ�J��le��W&���d��r>1�=6vB��m
y�5U��!���2'}�?`��R�e�2!1,�ަҌ��5��5��(�<G�^��qc�xN��ｩ�T�G��{��X,�Ғ&d��9Kk�mN���Jo�?�0PLA=>s�ʺ���d�c���뼙��y|7e�o��w 7�����7���gɣ���<b���:��ڼ�o_x���!���졾���k�=GK_��m���	�hUꭷf��0�<�'u�3E踪������I�aS�C"%�d�z��ϟ��9d;���JPoG�P��n����?!������-���i��bbP��"�&K�(L�w^�����Ϻj��(�U_
��ԢRl��_fcW=�u��;$NyH���Be�=����^�����T�seB��>�
�K�q]!C��U>��sei�=}�bp�.%��I����Q�%/������4�CX�;���RAO�sK|o1�a`ɶI� ��1��=���HL�1�fs�Q�z\E��|�6�z|
��̶���B�����!:Y�k
�_��3��ھ���J�h��p)&>	�PK��q\�����'].�P|x���X��3��@MZj�����}m��r��/[T�9�A���5<X�NZ8�,�!�5mĨ�"]��$Y��a�bP�̓Y��f�)�pȜ�.!�S�T�����s-��n���-�����ˉ��V!�GX��a��ѷ�# .r�oS�)�ۿ�(�00C�;rc'�ω�Y�S�\�Un��>��SyZz�� ˦,碓���y@�l���J˒����"W]�E�������{x���`Sr�Eo��g�0���0Jp���c9����@(�m�V�;��e�d�a�iX�f߸F�x��*(I1����<���˹1�����z�)��I<�k�@�����K��g�1�M�?W�]JT�z�ěX"����X�@��CG��a�]+���rHc����=�T��a��m�z��E���q��CՎ2 5F�x�SH��|�2��r<䜻���Na|���5UߧQ�zadZ��*5c(���%���9н"���s<
��q?K+T���-�w��&jX>��؄a����6}	�Σ��"���������{�e�J�{,9a�'}EQ��(=��?�9�˃ǐh�s?��@�#��K9����P$�CC�V�^�� �
��2��@�\�����j���q��؇$��4��B�T�YYZ.#{����d�<^K3�`�����ݨ��(V���D 4��Ϛ_���i�jd��d��$[Y���i|[{�m)�t��쫔�Rѽ)��?ϰ�{�}�\b}�h�������,�M??+�*f�������TL�Xϫ\G5����W�Q�-��mE�c��S��(A?Q&;��J�����Z�o�Ê0׊����7����Κ�y���g}�y�Z
�L�~	��B���oK	V,
�����?��2�\��L��6L���>�����T�5����B��,�������u4�6|�Q�mR��/3~2^�(�<���1�@�E~q�w�(�Ň�?�?��(6�-J��h �9s���(�p��C��G���J���4'e��8�!)#��&��g�-���h͑�8pɮ$*��)�J��# �uznW�!�#Rn>�}}p�*�x�׺I�J�ɃGU�7B��<`�n�{���R&(�����~����s���M
�OW�ޱӸ��Ce�$xt�^�����"탸�qUb���<���/?l=y4]��<e�./�����ÜZ�΂@�������SU ��2�Β��KQ�sM!*�Z���}#�5� ��`����R�ߖ"TsKE�P��r�){�	�<[�x�?7�������3�B+�5���Wz�����&�Ρ�a�DR�V���U�7#K��Dc��ſC��e�k�y/
�(�`*��=�����9Νp@6��q�=e|_�3�� ��DH<t��a�0f��
ʒjzs���8��,M��X���S���I<��q��L�7��g�U�<�ﯠ$�8���8�l�!9��x���|��~�3�~���o؏��Ǫ�笌��U�t� K�j􁜰���'V�[S0,%�K�N%��1�-m�TH0���1JU�&^�	iv�7Eav����j�9+�E��tl�A2^��y㚖hS�.��"����KL�q[|u�'Z�� �L2�^_ų'�[e�(x~�
� �Qʒf�K�$�oEg"�s�U�dYN�4OC\X0Kt��S��1�ޞ9��;� ��;_�?P{����[��2T��<波�]��	WI����>$��u�<r���dY�a�;!��l�� oQQ��4�^��C!��peey�u��J������/�[��a���!���5��W�[�{�r�x��Ep$&�u�����g�Z���M���\Y��bAI 2®]�J���	��L�[�R�e��6B�7��Bv�����S�$e�Rr�c�,��2��|�~��m�˛:�B~�������HɰA�1k8�u�����5O��W���r7����1����O�iֻ)<x(8[��kιR��U�s�k�,I���P{a��]�Q���@�7�bu��2�2�lq��u��o.e{�� R�����l;�j���b�f��1�Zh�ZI�#Vk�R:�gH��2-0a}M��U�Z������h}��1�w/������|��[(�+xY7/_�X�+��9�_}�Y�K���}U�$5���6�[M�y�j�V��Z�,Q�<��8�9�(�cR��� 9fz��z���&��M�'4�ݡoF)�� ̹H��⏫��	�� �RF�,Q����&�%
b�Gա���T��:�8oA�B�JǓJ��r�#��gn2�=��:�#�����Տ��}����ֿ�#�)��S>�˔����#�|�"Բw�)�ױ6�>�fc&={ڰ�m܆K��Hz���"%���[�gG���W�s�B�~�����S�YG����`�X�����ux��!��3��^]Y���ޗ�E��珿UVd�~��5����[�2�g���R��w�>���T�	c@9��/��˴�V��=�)��es�GR��3� s����k��eD	�"��e�.���I�$�m�P%x�7�E��:q�=��2F�
r$�F�h����fŭ<�k�+����@��F\ Nx�=�������X=㷝�'�~���]�H��&y���b�Y������9�]Q������&��@���~Z��X������;�}���lv�����ˡ�?�?8����S7��D�^����y�B`Cq�� �:���%K�\!�c���|\���B! �~'�`Ei)���Y�ح�f3���"�!@/$^��mɈ��"0�y�mn\e^�>�m=ȏ��}�/�{��Cg��t)Fɤ���A[����yE��F����~�̄��U�Dk�Kg�Z�����W��"�t��w
������}p���	���x��;O<_�g���<�/����{����~O�_[��FF<��k$���ح�Kl0��{�_���e�����Hx��!� nU�����v<�0�k����z��2/�TY�9
�Vb��#�[�Y��I�`���:���E��6���.=�-�BG0�ԋ���D%.xb�����wܣ@���elNRm��;2HQ�����Ė�/t�G"�!��0�%QS	���-.� ��K�q>'>�_0�?���q����a����UX�i�DQt����qc�z�\�gy��	����i�>ןCyM.��EaNq�U�wf�!Ǝ�,��@����N���j�n���p�
�K��s66���߁1j'�=��YX�7o�|��/ �|��m�ol�4	l�6F�*�(Ŭ�����B+�4t�ɚ)��j���0R���>��֋�TJ���V�!pOE8{��S:_�\���f��ӷ�S���0. ��$�k [5�����`K,�P::���3"Hp����F��;���2�g�^�~�Xy}O1L��cX�Q�� �`<3�������>�M	��{��o���hK���A�O�
���7����祬�FhU����G���&|?u�5�>F��>��Ħ���.���g:S�F%�T�ϯll�q������y�<��}?6�k7�!��Se�s�ݪ����e����4�G(�T#q��x��VA3�����Ġ����[�bI2��i�5A���#�"���Ự&���1��g0F�6U>�4��a���C�nƳ��S(ow���G��&��^���e�H՘@1���>����7(B q�7��wф�y�(W����!�D(���B��H�8�xNl�Z����൛?�F��8½�c$Y;v��
�ڭ�w?���O���*�ȴ�(�IH7U��'�ߟ������ ���d���o׍���Q*�KE���iy�4
;�e�����,M�,��Eګ^_��$���@������h��;��1k����V��>�+,�}+��UΖi�aU��f*ž�i�Q�l����9W&�v���Ş�O�z!a�ƛ�<҉%�������l|������g���M���b�3?�^����ﳦFk���+�ׅKs~����t�ƦkC���-����)��~��*�����%d����,��U�"{�6M�#�L����e�.ڥ�uV�_F����]�c��ay�]�`�^c?��s5���̚�"��k��v�>ch��4�VK�#a�n
곡mݶ�X���H��i
ݴ�
�#�`���q�H�%;��vHuHa��c{
{^�����!"Y�z
��"Jf�r��$�̦�+h���iU4�d� @�g76_2'��W�l�� �C�P*�聚�IZ�4�"^��>\K��=�:,�-Ϊ()0ɽ���z����_����!i̼�P�W�/Safee6Bj�bu�Vr�i�x�����<�_��~!F��>L`�U׌e�m�d(
.�=h��s�z�*��G;�1�-��������ߞ�b�Y�>��''����=)���my�v��Jf�/���soG�e!� �3S�I�G��n#잎<-�Gz�I�Vp���+7�M�x4�9Z���*^E)�lSR)��v7�@����u��ՠP�Ca��T�8v��Q�c�Ê�
c8��<n��G.�_�8�����1^�T/��#T���{)��ͺ&0�T$�� ҀQ��V����yIpQ9�)�yBOG�f���Q �Ih֭4�܈n��ؽ�т�Z�hն��*XK�t(��t%��?�Q���I�B������j�ĦR�X�戠��F�Y�z�5�j�HA�(�8o)�@�B�|>a�>q�M��G(S4����C�����<2vF�Ҿ�+�Ӄ��Y��)*�N>��yLb����(Z}m��`d������|�J�mj���w�s�����
i�N(I��mis��~F��!���ߛ]�����z���p9$	}����Z�{�U%��>���_��ޥ&͂1F,Py�{�C��h�r��7n�q���閱��qvM�)�B���h�����a��c<�yNJOP
�cB#mM{L�����FM���C��ֈ2^�(B������<��	��s���?��]�S��;�u��kN���B��2]��Iw��̭V`*�	�mg�qX\W���D�RlBF-^�ՕA��Yu)�P?#�S����x��i�v�F)�J��O 5m��^�Eď��u��~�#���s��54�Nr��P�#���tn����"��E��d��O�xi���{��ڵ��l!���
&���O�@�0wUOB��$uaЀR�@�Qv�1��<�%�c������^+�m�.FR�w�F}�y��@�i���&���6ՙ�#�0��7�`��s�=� W@Y��ŉg�Ѱ�B�P4n���yv���F֞R��
K��2,̙髕´F¯��d�+ʵ70,���iCc���K�I�8|�PţR�_��B:ߏ��O�V���%��x�
�p��������@���EB�C_�70�զ���-�]�fw`�,�xeY1[J�>|𳏪F��[�N�7)3@��2�8�I�0��^����0FO]�b��pΌg�)�@�γh燷���u����V!���.`;7k�un��r��(��8�$�bX	���Yԥ,��`f���s��p�*iwX�RWl���� 2��F>��7Ρ�h��HMm���ڏ��&M�T�9��ЎG�y�G���z�^����t�y]��u�I{���k�f�<��o�Ի��8９�a���r|$�RmT*/��U�!��¼�^���S�g�����T�LL�6o�H;���蔀�V�
ɗ��5J,�߮�}���OQ.��_q���=cm���y��YӒp,�����(�p��ŀ��gU�'��ݑ��¹��=K{����$�cf�i<��(��$��0~��|�r�B���i$3B�xEzgŸ��πH�g�O���eR.���ˢa1�ѻ��w�J͎��.���K��
w�6P��2Ů�MͰN,����GNpo��P��9���Nv6��j��ۧ4���`嶴��d�����v8fcey���U���͖�~����V��$���W��Z��8��0�2�[A����a�g�d�nr��ph�ci2)���`����G���������ޑ�m���O���5B2�A���a�\}�0���Z[�&\��z� dWi+߼I��p�yU��4�,h��a���m�OϔG�A���ϒ�}�x�Ý7"��
�n��M��^Ӱ�A�?�u����p�?a��<S��>�e��$��������0�>qe�𨹂Z�*M��h�G!ڤ�J�٪Gb��a������R]���5�
����͋S�
�R,��f1�)�O���W�Q�96��[k_�h���˵���Y�Ʒ��
q��i�����l��ORfͪ0W.����`O����j���˼�`L������q���Yuf���`]B�6�bSV7�\�h	�)k�Nކ��7�^4N����w�jޔ�ʽlY�/{�L:�b%�x�lc��\�xT5C��R�9v/�<y�x�+vwG�L_��8��	�Z��6��<����!����[���J�a�~��k���{~�
�[����S���9W��6 JPVq?:��~�8LSo��5ĜC�ĩ�m'�����[K�w���s�C ��H/����؆y�~e�b1_D���1}��=���B,�H"I+����`ޏ���U�Yߨ���[KY�h,�Yk_����^�2�֠u}O�y��}D찔"������@S-�C �T�d�"�t}h�>G���=G�;�y���:��q���7k9&^�Y���w>�����8�l�}�f{Pw�y�B�|�={ƭ?~}%�xa��=(X&ISQ6��~�=�K�*0c�����wPx�����,�
��]Z��ơ)�V-�f��yd��v��~�F��;�;+�x��=�����{h�X�!�VT�I�ɚ93������Y��}['E��P�OC�Be�:IE����x�ia�cJ������Ur�Q<��!Q��j��P[F�>^���$!:4<&�ɳ��i�)�N!���]�/n��3z�{(�l��=i�t���PmCE&�^��&�!�-�@5�1���mr�u{ e�ݣ�=��O��1�L�(�G\#~�f�[$��ڭ��:�N'
mh���ۃ�b��_�r���t��g@��ۆg�n�6���ʂؖ#�9=IZC�	��%r�y�2��K�2�.Foւ��B�J���Pt�sk|�k�|]:�	��6��֔��*B�Q��b �m�����a�<,X/�p_}\KP�Rm<��Q�z.��I�w��ۨ�����N&�V�$�b����h1S���F�9�z�!�jXA|�g������}��<�γ�� ��/1�7�.��_6
�nƼ�)�^��uR�\a��H<'��b���e�^*��|5���q
���^@�Z
�2�AB�2��W`L���@� �4æ��1��(�䖥)�����=�}+�|�ֽ��"��J+��7�P����H�!��d�BP1�>cZ�d�^�{뤈 ��@��$1����������(�h��*+���3_��U�_U^!�box�s�_�ܖWۤ��s
�o�����xs��'�ai������"�# ϯ�����[b�k(������e��<�K`��Jś=��.���E�4�g�g/>x�=<��>� x�sG+(�t�������.;��c��K�v�إw`q�2-`>}TqF׏kK�)�fl�+̚���g��=w�S�/���%Q�s��:���[����xU����S�����)�l�a!��� ��%. �V��
Vr�j\`�,"���/�RU���V��f!a	�;E�(*��#�4 S���/������\��J+#�O���M���J�� ��#!�q��������ҁ�_	<��BɊ/~W��Q�)�d 
M���i^`Y�2����k,���Rqj�ΔTE�a�]���2� �-�]]ֽ��WE��|7�]�,�ʘXp�%eBie��w�^�T������)�+L�L�=���c"{���Ww�\�k�G�*��"�U���zxb�On����ta���-����;��>|�<�9қ檕�	��0
 m=���C�(���x���ٽ�����DQO�h���Ttc(S��x�;(������}�-��wy�?x�ֻ�}^�����:ic�j�"FO��Fk�[6p�Z��"�z�(z��*/\WZQ.pid@��k�5��I�J��B�
�n�gց{�dޫ���y���2k����o@��'�UV���XI
.F��L�O�&�.�D��+�(�y���>�ŕ�QN��
0v�6�������:z+<��]0���g�G�����g}�^��)�<S=�_eǘIڎ⊒�}ƥ�]�k��U�
�ԥ��BN
�0��^<DS!T|�x2G��BkھJLF�-���o
J��/�S	��za��Y<%� w\�S0/M�Aa�OX����~��3*��)6nŝ���(/�4WVe���*�->_/�$|�W/I��B���dY-m8fF�/p���˳>�@b����%��q Cw�����5~n�^���5Cw�Q�g%�`�;i�c\�8䑵Y�6q Kt�r�Z��O!Ԭ=��bpou�傄$`Ж���[��X,�vieip��M
 ����>��N�<n%�J�!�g���G��򝞢�?0+CSc)�m߅��X�˷��q_��9��҇���M,0�){�9J��u��(�5M�[�H��Xe�ϛg����[S����eJ����l�W)�����E��9w�����}�H �%��w��fLs|	Y��ELku���z���*Sg��B޳_�pE���E9 ���ުYiW,��~
�*k��y#�r��	�~��s�㻿j`^u�$ܟ����yY6���:�)B?�C�1�W�Ͱ�{QQ�}�!�Oak:B�_�8`�x�ʻć� s��owq+���=���^�����^��&woCtY<�Y�<~R��J�*���5@oG�4�E8{z�YQ|�l%�uƱ��J}?6���Z����o�>�1;���,*?�4F����sGx��1��WqI<�	��N�=�_��wL
E��R*0/%�xs�(Y��0�P�G�>��>�x_�}�2CZ����aj�[���ޚ�9'��.`H��HY�r���3�B�؅LO	7�`v�ȃ�O��p)v@��'�`�X"�j�t)4*�~��U<���ч�W�H5`$�Tcz�a�1y�'�Kθ�O8�.�����͒�w9I��&�$3�0������qe�sU��K���_+��HceLq|����4i�=�U�1v,�ժ����ݒ�X�#!ܼJ���ߚ"e�vyU.a��о�|�P~���~� ]�{y������W�}(�o_�:/;N�T��ֳ�r�״W+t�^�A,�u��>l� �%Qw�2N#t�ffWp�
�b 
)+�t��U8dZ�x#�����o~߇��ʥx�B�:�+��ח�b6����+iU�߰��5��}��N��W�4�',���JCO+/�E���q�(�M��z�rv��J�w����{e��B�s����C<<�n�_:��Ve��G�;�3�PkkD���\�.�������"������Gֶ��/��j��,�%ԯ��R��`5�]�%Z�1B!�5ne�5�K�*'�`��ojr��P�}�O��'x��NPLWv/Sf��0HQb��EI��pL��c�FP�X��}3��[Oh����x$�o�����RX��K՞K(�y*���o܏�� >�ܬ���}��w?'^�3:�_'���#]wS[��,)��1�67�<�g��䞚�V��b��D�ٵDjlt<�����ulƬw؊5���&�8�]1Uz!@���:m��GPP��W�n{���=� �r���?|�sF ��pEr���}��kώ�ē"�����`�M �t/��7��<��3:e���22��?&���.�ν�/4�oa�r
����U������=��A���S�T�0l:��o��a�u�������ʰ���	�ڽ����j�Yg�=Pik�Ԭu��~#.���`��Te��Z�AE�5|�$�V~�5T�8�˩�${D����c�D���%�lPݚT�P���{��o�߶&���8�m����I��>���&���W;��=~�9�O�$����@��Q�tn���|�<���>�;$�XU���MH/*�O(�F�I���2P�4��<����v��Q��l�M��X�����rup������&��.��\����2Ÿ�,�����r B�w��kgzc��e<�]���:��&j
��H2]�8�s�7x�b�G�Ӏ�}��]����b�F�%�0�s�Ys Ί�缜ì�8���2�<t%B��Û����y���?��	�a��{��Ƹ^zc/�`ћN�	���k�P���9=Ϟ}��`��
��̾yj��S2H��r�;�nr4�� ӎ)y�%�}��b)��U��/b���<��+�x���a��C�)�CM	�ϱ�uZ�%qA�{~'$	.�r��Z���$󼁒��ň2MB岍�|
d'���F����1.�W�U���q2�H�-ā���Q���x�yD�I�:G5C��6_��q�o�����tW��*�m���FġĠʷ���!������8�D(�D��Ё�
iՙn���?/v%�K���= ��x=�K}9\��N��7�s]2C���q��d�'w��x���>�P WvԼ��؄2��&'��,��X����������}��1�?��?\������2�^:
y��C7����~��/��+�P�����n%�g�ҊK^X\[/��FKx��.kt-r����s-�I-*3�)FUb�a�
U���$�	At��N�?K��t!�"<}���H�������N��O�>��X��^�]�J�k���Ky�������r[C�Y%d������?��nY�%�|[�xZ�,�};Eٳ�)�7u�H߳臟���������{�E�;�c�_`Ҕ���2�Ƚ���r��5����dy��^R��<-{
u
���W�*�f{��?3��5TiB�v��t���/CY�z�9O�p�������ib�q�V�Z�|)�txK*Ī�Z���U���ګ���i����t+��m���L4�*�����(���*\c�03Y�v���;<Vi���T�X�lQ{Z��9c�YE��y��5G'��.A�=��Di���P�l{��`��=��S����(�ԗm�{u����Q�:��{����c*�T�����8���)�h�{����<��>�w��3$�o֘��� /�;x���2}Ħ��vq ��Q���x�Xn�$-�݊�������������p�%^��J��0G�~�Ol:ŵO��jSz����%��#���}��ѷ���9��Ӟ�+�%��ȿ_% �S���y�'��s�>J�o��Y�BsX��Z���/�,�J��٘V��⬉7i �n+���`��zx�
WQ�nh7Ȏ^�E���	<�)ηm�=���.
�ƪ�e��rX(�2����l^�ٓ��z�<������_C}�#�N���Sc1V�0
�_�<_��䞆�*�Oz{B�Z�*�~y�ıQA�1%İ�e{��w����I�%A;��D�E*��0T�I�(%ƚ��o�ZQ���������P��Y����H墑$_I���i)����T[��pm?*G�]c�"HE��h���R��A�k^-��a���2UЗWQ!�l�̾m7+�}Y�����S�J�2=*�زc@��	�:{6a �l<C��#�g��5j}�}��a���W�7�!�,� �:Gl��T~o�ax붭�t�cܺy����#����Z�Wn�[9���m�%v(Z�c�I��Ʃq>#^�?;cv�y�����}O�f�E��j�k�)F�!e�$�L����r
����s�����B�	�0�ևKSx#�Dˎ�t~�'k�!�S��T��ex�< ��-��Æ�˄�E�y߽��y]!;,0k[V`��Q{��??B�O�V��qV��;֗���r���cݟX��c�X�z�l�+�g�y��x�����ցi DE���f쀪��1�=~�wF߮&�W>k�rL���ߧnh���\|��m:^E�y�b�}��d�cᶡ�v��[��2����ᰧ���Q9�>�|�%�M%�"�KO��t
!k�z�o��`]�Q�he+�6I���J"�c��mZ}�=�U`��$g_�RmQ�V��)JaR���ʗ�[i#]��V���9��8����Hv��cd��z�J3c$���V>7$�y�N줎x��}�/����4�i��yl�0���ڟA��Q�t�|AO���CLyrߊ/_W,pt�-���:J,q���KTᙃp�`�l�ow�8<yHE�c�]L_by��;��`y��b~�����C��iSv*'o�vY�?�������1����w�_Z����QhcB+��C����2��m���쀄-��h�ԨI��G�Ibxד�\�VaEjt���{��IS9h�4�suph�q����k��oR��y�X`�<�nߪ�+�a/�<e5��U��2?t�_���SZm���P���+�����N�u��{�m����:�|m �}Q��X��<|�͝����Y�$�r��:Ў�p7�p��0s������8��$�1Vun�.%������w�:o�{�)��׷�f�������$c=���z��"���Ga%*`C�)��{�F��5L:�,�q���Kg,jOD�N��F��`��u�р�f z�tݔ����.��}_��Rj���B����%��lk�A���mF���m/Y@��?�U`~��V��w�w-�qb�&)!�F�C�L��Bz���W���ܥn'��tmX����%}��|M1j�-���^�o� ����H!��j��**}���ps�c��:/]H�=�K_�t�0_Q6�@�������Ï�[�ZF�=J�m�lچ]A�h���8e�
o�L�U��D{=�	<Q�V�]��8n��j���(�"�L�^�Gd��D&e�;E��R%��H�g��;9�Q~gʐd�$z���^;kWG��������A�C�6��7e�L�{�Q?T�]��Â�U�n�a�h[^Y�g<¾'5<�R��n	lW>�f��X�B[;��0��z��Ƭ�����W���r�5'awwm�Eۭ�!#�*��v)�e�Uf��x5�潦[���+ƌW������&�|��������
����^:�>ﾯ�^v_�;Vv�:a�&F��
t�TR�������g���=EA�4�3�����Y=�����K�?��h.ٔ֙���-�R�%�Q���W�rR�'I�i��p��I�c{�3|�}�L�ak����H8z����?p
�ߣ[j�D)R�
\��-9�4��|C㖦��la�Xt�=��۷G��=�p���;��x:�[��6ޘ��.S�E�o8QG��^/TXQ��؏s�e��J�Ht�d�G���Q��/6i~���q�t��@I�[�}�C^�c�M<&�i�=�
cԤ����i̿���X�qH�\f�w��]#�aͩ�O��B��B�q*j@چ��=oH�ѣ�Y3���Zc��2�A���k?��I�{�#[]�:O�Y�^�]���N�O�#�a��c ,p��#TMl0�d��f��E�E��[�?D�]DH3���r�{8(ܿߌA�p��;�r���7!X�=��(�����k��/�� ���>��o*��kJ�Va
�H�8p���S,�o���(BmE�MSt��b<�n%�L�|���F���f�!c�������}����2�A��D[nVS���r��� ��s�`_������1*<�t�>�P=@�����e�y���=c���[,R?w�e�z�ֻ���� -XG�=~��z��^��'�H�0iA�����A)�J/xRa�קWwVv��O�6��L"�+����:�;)|W�*��*[Z�g�#�6��B!�T�!�:���~���Mӵa
��t�s��w[O�(��ٳ'�Ac̨�ii�K(��7�RUg��ZKs��IV^���Fa�V��T�c}w�<��O�0���Pj*[a�����u����%9Kz��9��7�A0Ag{�@����X������v� %Ni*�?�	�L7�.5ll�6�5�o�cܸ��Q�c]Y4�7��1nh^f�qO׎
]��	T<� ��VI��(�T�ƛk�f��?|���ګ6�k~�֠Q6��m^<���X��#
N�W��.r�E�y�qz��+���w���W;h����<�b��B�F������/��+8ZE��v��8=��
湪�����]�W�/]RT7�\��x�}�o�����g>�y�N��3��s�Y��}�w������JQA�DA�2�|���u<~�D�_�uͭ�NK�:�1#�7����Q`�sIƩ1�A�r���q��S)9+� �RM��������x�Q�!f��Q0��F��|�l(h�;[��|Ŧ�c%���_�)7��%Qo��o�'͗!����ű�VǇM����&$ďQot�bسx��`�K�(+�^��N˓�x%��w4�T��2b�:N�(�� 2O���߻�2��{˖i>@���jףo����	�s����>��Im(Ú+<ƍ�΀h��1�^��ۭ�6�i8��iO|i��� yѪ�R�햤"=�C���S�$�C���:U���V]ڎr$����ze(k|��P�v[~���6�N�[��oM���oO�����0��E5�C
'4��|7�����u���Tߓ� �B�{��s�,�ֿ[��;�ن�
�����:
�0S�ͤL�-ϓ���Q�j�zI����f���<G�c��(�����c�2����jl���X�?6gǽl솽R�ݔ�}�ZY,�{���Bժ���(��	!��4]&ǟ��8n�D�Z�P[.u�f��w1��X4�L��
l�'t�X<قԸFU3B��7�Ma?mqg[+)��S��U�i+�U��<>��
�a]R�%Js
�� Lbl���>�C�h������K�^y/ ����)<���eH4���<�I<�Υ2�~��J�s�����2hM��<�&��GTuR>'?�{��@Rcʓ���~\g����h��	rEt�֔����S��z�R�8���q��a�5F������\PV����WE:�)��g��Y�0�N��k%Fr��)L�֌�?A�<G�y�SM����$ޚ"��p�_���M�oـ�����X�F?u�z�G��羈G�͢�
K��$XK�w�}��Gk�F��(�M����`�s$\´N��W
��^���Y~}e�����}>��/��~Ț}�w�<���
���U�_.�j�G��8��KaP_��M*�̹����uإB۬��'?mF8fb�A��[F�s��0�}�#C�޸�B�B((�]�u�Jx�Vh<�2:��S	��Z�ڣ��Q<c�A���.D�����u��0��5�;�is\��$�����8�='��0N�]㊓(V�*U�H��	k��r+�AMyF�O�>ؗ�)1Y	.� 9i'(�RFVx�#t��>���r�=#UO+F��k��sj����Iߏ�q�k�'�ȩl�?��B	Y� 2M,�u)i���_i0�>�^ե�������1�~7�0F�!c�~��#�-��i�O�`0������_��K<hy�!Q���~��mH�N!��}>�+��������P妐�Bt��@oݺ5���^���x�]�?��̯���?��?տ��;Uv~7�E S���°`������|��E�_k }ϸ��E湏+پ��h�<��J��2��z��>��1ކ��1�,;���~M�C�c��Ԃ&D �㨵o����X�cL��;3�m�˗W�P�G���g%�w��;��6�0��d�.I�~{���A��A���G����@���B<Ċ][��2���C)M��F�G�[ȽJ�)�&���׌�		��gl������������}G�LI�	�I����r�1V���s��(��J�[��>������Z�b��
J�sc?�S�fa�K�}�@Λ��׍��J��(�~�Wf�j�;&}�5rP9%ф�Z5���������o���������A(_c2� ҺL�nK!�O�E�B���ʰ���}��{�����w���y�a���������*�x�^�g<�|1_.��K_�'X�'�t���s��H<��"Pc���#\�B��(��4R^wMdm+���"{tVs���@}�tX���v;'.2�}�~/��R�z
���0r�<�s*�J�y�z�¤�Q�8��������֘�15��ˀ43QJ�r]]��'Գ��c�^����؂�`0���V� T����H��\���م��E۹[�E��L�3Z���ڥ��>y�����̮,��D��Ph���R9��seU�)��nC�~��)���g0�'��cc�>?l����e����M�C�YC�sJ�L)5��)"������X:yCq#
I�*o޸瞳��k��{������Ŋ�R	qs��9�j)��������ηvͦ��-��e�F�/	��H�z\`}V���W�����yr6�w��ċ*�"��h��+v<l���*gڍz�:'��+|�^�Ћ�4�eOah�H�	�dh�T�'@�e�U���5Y;��y����}�.x��Y;�~��)�|�e۲9��a�o�t?T���:�����$����ݻ�HU�z���VT(V���N�';73��ho.�Ȍ��8� ��	f9�f&huE	�-`�,�	cc!�E�͎;�Mm9"�i����g�z/x3vv���yG�X,4{f�9�s1_�k3Ϗ�ό?ϳ�x���=K]��w�8�z��8-��Y.�c���
F	��	�k��Q���(�:�j�5�4Y+`�3ce}�9�n�cEx�V��ׇUrxV�q��SRŽ-��bX�a��P���RGFƕ��L)E]n_�N�R<J���3�
U �4�T�+V����� �τX�f��8܋�VP�װbV�t[�+�G��WR�Q��U���9�ϐ�������*?I~ |�-�BE}J{xP���:�dP��<G<��懚i%��LA ֊�x�����@�zp_K�H`�+<Vu���5���<�e��ϴM%\�.�Gx�=ε�i��v#�O�o�Fht=j�*_Ե�d��s��s ��o�����뿾G���]�~Xr�&{��,�M5��H�9w�����M�A 3�,u�s�{ld1!��6�%@mL:��[�A�07̑xA$Gv�^�0)3�[��=���۳�������y��u�&��d@7��@x�o:�62���q̉�a<�yYʀ12�T���-�v;D�&`�0;��A�5Hm a�\�H#�b�B-+fk ��Ȼ���M?3olkH>�`0h�GeO�7$C�4<B�i�
��9��1�MH���Xrd"1*���������
bgר�UOH�����J�v��h8��bp��y��s��Ca� �1y}�>t��_�́K�� �q��]���眨�^�?+�U�Y}�D��"=���vh�fӃ�;k|�v(ᙴ�7��'��xa������ϥ5N�G( n�ªͼ��-�y4��O�����,�Y�j�yg�|D�|�<Ic��D�9fs�,��|�#c�����7�&��"ܽ"H���j���:g�i8�n�uMUWf�ߧb��nâ��g��X���������b�۫��Fp�=���L-�à��C�N�6'��w�S
���� ���q\nӓ�����ҵ�\�;���[��*-33�
f�w��� õ�? �N��nҳ�>qf8~����Q�&"�$e�N�J�0���O��
6�Rʧ0a�5��f�����JRZ�6ەc��P�����	� �p`P O��n���+�0yx��q���R�l��)�{�4���M1{�����T�}���wn���fI�L&�����޽G!��^qRp��q|�1[
��%sM�j-i�A�X�� ��\���%���Y���Z�ڞݮ+��%t�u^KYj3���'ҩ���vL���f^�V�[�����Ѯ%K��l��]k�8��*�Śb�D?'���M���_��U�&�������?���k��oz�v�h�+<�I���f�i�acyV�y73W�9St�Lp2�蝻ݒ�W�� �*�� ��1#��fq��G��tZ|���I�x���U06v�����3��W�Q�~8�.Դg	�*T~o������Vyjg����d��RE���0�۹��y-7�e������D���%�~d�����2�\�c�s���l�c'�� ��P��-�Ӫ;2 X<L�U�veHYK%�-��veaxr�F�S�?<0��bΣ|Q�%i���UЏ*���X=" �a�{.AzN2���_$**(�([chF�I��R@�O����S�1U� Л��+%�[�U)�֪R;�Ww������uۖ(ctRtxV@�S���P2�}{�G�Fd��Õ�����n)�D?"ś ��L�1�d�j�d�)Rc`H���^����]���i�y2�1�^�^cY��D�UT�(^��r����7�7��Kb����YC�-��F��r�fu�|rm�]5T/��5ڋ�|��|:�7~�gvDA�G���i��"�t�w�nh���3b���I�6s\��5�I���n���6��]&f�)�lvۖ�m۳$�Tc]NZ�7���"�F�@m�S����z�3�����=�覢���l��_i��Yr`�m�s�L�9���;`pϘ��'>K��C�U�l�V��^����yU����g]�W�q��9��et� W<�:F�M?��7���ݪ�pP�LnLj#�U5�1�=+�O��THQ�cc"��1*_P���xw�V�N�ed]�s�M���o�UA[��ݨ����$pǝ�un�~�@�lK�;������g�<;�tCJ�(��( �Xń�+y�d<�tx��=��Sz!!"92��fg��>Ϝ�wv����sM}=�[�d.)����;Kw�z����A:V�ҤU���6�ro����CC�~����V�jl�!�v3�\@~����/��/~R`xD;N����D�[D�%V����v*�/ z�La��Xf�W�سT�X�X��00��l���:5֋��s4�fQZҙ�Nzk&�\d6$R��l�x,z�egӄ�x\>�~]	�f�zݳ)�5��4˚�<�ɮ�ǋ٫�>�� �5&�;<�7k�f�	�18�3%�cŋu��(k���=R��TDE	s�|�l��d`��Q��;@	v��"h0|y\S�?j^���!��$5�{��ް_�S�H#^x�9�gO砤�S
U��.jW��q�R��s
��q�G��:����!�[nWz4��]/ivmx0��V8$ _%O�ExP����r�R�i�[�(�	����2U�~����Tp�����L<]{f�>4��6�� d���,������ {�2'�W�%ϙ%1:,-m�a�{�6�k��sQ؇5w��
���l��mĽ˸K�1NEl^�B�D��/hL���L:ׇj�������_��_~VǇ����:�mZ����γ�{zw�t$��T�zh���j\��L|{�:X���W� 0FK�YՖ�=�*����E������y�!�8c�.���`�	(�l���m��L�t%�����r}��l�y?��~�i�͒�B�\n������s�� �$jt���B�������M�>��-%�dH������k�O���V�^U{�٩�9>�t
�z¬İY� I��ܪ��^���/t���<�*H�fY)k��O��7E@��f]s�T���h+6oRh�ڍ�m)���ƕsd�	(�h�U��!9Č�LB� g~�����S8ik&Rŕ�������,2�R�PDUr;b�t
�����N2|7��$N[�|�M*m��=�5Y;��w� oq׆�Bf�*��K�V�r=o�` ͼ�`��c7@�
(��ΪͲS��׼8�L������?#���zXEދ#zp��w��_��I�"e[��e֛6�l� 3�f0�3f�ygo��_h�횁yCa�k2���&s�|��	�S͊��Tc�/�А4`����h��%�,�3�+=�J@��!ɛ4�k���axp62�3G>��`���~�����Q�׋B����Q1�� ����\�̸x#�t̿�AËP��f����
 @���)��B�ˠ��۴qSg�jl���$@T��ȋ�w٨m�o���$�-�NR	@0�'ʎ�H�*.
܈t�6�E��Y�@q�!goHG�D튗�±�!�FS҃a�,�:��0�&4��b�>�D�w��P�"������6#���	�nj�y4��>�g=�[ӞAW�(�aUi m���*״�k�6��Fh�s������F��m����T�O�{䶅�����W5+�G4��y�O���_U �[����_��W���e�?)uڟ��C�^\���Mp~�Qb��b�H9y�}�D��̈3���g��qx��f.f`V-g@�*%�ds4�]��;�q�</~ ��AՆ�t�߸�#�"q�B�r�6�f:_��i�1��и9O�9w��d����K���4���ę{�p�1��A~GJ�}�Ё�\���\Ü��M6%$4��=���@u9�x��H}�3��vv�©�ݹ%ż�C��|�f�j^�I����:�Ⱆ���z��Y��~��RY(�m����R�&�(���[%�ѹ뮻�V�B�5	� ���+������
���))�F%���fQsFC���B���ݔ����!�x���`���G���m1(�����H{x�VG4��[h�������3{x��'�pJU|^Y�,%�Y�{�V�"��`���,���l��<ٶ��$�O��s�y���; �:�7Q��
��nL��i	&�pՁ�N������������;w�GI�okB>"��z(���&N�[ȯ�W���l��Ά�n�#3#�y�1�&ý�<|��Å�!�2{�2fv�f����Ҫ�8�����2�z��e��1/hg������`���H��!KJuhAz�4�|�H(��1��5�Y�\�-��Z�lx��ެ���A��ƋD���j�`��D�.��E;�K׌�";�߬P�|Og�$����:ON�uuu)p���C�*�^El�ѩTkg�tsF1���+V(�Vy6W�R��@�|�K��oT�@̫]��	@C��
����H��/ɏM0U��	�!26�� �!��Mc��隥1溩z�f���?�!��2�gNi�jN�lz�����X�z^W�c;�ѾA����ͳ��5k�!�&oY�>��nNӫ- �#���y�������ߓ*m���h���"���eV������ٹ�fS*l��L�f�bV!�6�*�l��L�{f0l��)�ѻ������3d�eH�^���+�l��}�4�)M����?�"���4�s�ݹ���J��m�ށ;f����qJ���Ťlˣ}���L/$�R7��J2�A���G�,mD�y�0xMY������T���[���I/`��PϞ/�@C�����TD����$��yH0&��ܣ�M��e���l��$I_ݟ<�0,J�EN�
z��k � ÀA�p��Xb<����1?��ZCl=Kh|�S��nON�yά��@h�2M�%���mW�Bʹ͆�k���1X[��q�g$Z^��^���Vֽ��н6l���x.��!�����׏}�����;.��q���4���H+��O�2�w�L=K��5�,�y�s�Ң��,c �l��5��m2��^�&s�f�J�0J ��"��w�o{���<�Uӑ��n��Й7/���D�%�!�Q"lp�`�=�׮���:ob�L,��c��9�5H��U�F�A���>��߶i�:leH�K�!A��/��N!�>%���G�"aV���x-�x�}Um�)(��ȡc�z��IѶb��W
4�CY���Ca j0JzU�!���#	p~l.#;*Q�1�EN����R~-����j.��B	�z|��Xb=��MY�������U��N*��]��� �ꄿ�.L_�������v��f��F�x��ɧ���<V�o�⭊Z	�{��=� }ιp�!����>6,'��5Q�&���R�&�>=��,m��3�ف��6C7o�lIa�0��'��*�~����o��释�-�Dg�.G+�m�3�.�����c����1.�p�#�Q[*t�WTK�������y͹��a��t#�73��\���e�j�������&f�W�����?L��~�e�YM�xUq�9*�J��Ĝ��ɵ���Z�d��f���A�e ����xSb�
՟� VHնF�c'WF	F�{ yP�0$�
~����!a��9���Q�(�d�:'7�+��[�?�-Z�9�����U�Mp�Y�$���z�<$�f�Eʫ&��m�J�DD*I>�;cp�)tÓ�O�{~��  ��IDATc��9�-�qvEAr�2uΛ���f7^��	��������5!X2~کv9f?;-���He�ip�!�]��#yJ��y��ɬ����<:��yV�p�2�K|~��:a����O�vf��w�;�kD��H�f	���ڞ8�9O���$�1���D�륗^�OJ�;*5�w����k��nf�f�R�|���z�_���H����ߺ�˪n�f�@�O����鐔��m���[��?*.��ۭ�ou���I�̹�Q���Лn�[��`�gP�}�j]47���T���s�����L�6;Z,Z�"���!�$fl�q�sfg�H���E�-)������X����N�2%���V��P�p򨉖��_�O݈��Y"��kKjQix�t�T�S)���bu��0z{�/B��Lܯxm�&�c0ռ�}��3���!5���3�k$d�p9^�){��<ړT�g�+{��E�U���E�'5N���$�Q�,ő��NJ�qнC�����L���>8	u�6���e��Ϣ���"� Ҏ�z�y8;�a����5UU�an���T��L_�@Ȁ�Ds�_������[��������Џ������*����۪�^���|.c��b���L%�<�y��F��d�Y�g?=� /Ǆ�ÛA�;x�ߪZ�Wؖ�tȃ�.u�S|qOmg�P���H^3��f�5�~��X�v���r缻�K�q��ldK�Q�P 660h�7	?��]���Nb�`ʑ�E��R ���;����[N�6erA�<+����ɏ��fp�O����4��9��.�˒z�+A༑x9'좒��� �qk,��1n�KC-��Ν��B�x	�G
ZNev�@���B£})�K�쉑M��5��������nY}�ପ���y������e����W�Ϻm��?�z1^�]c.#WjW��RF�&#Ԫ��|�"i��C�M���Eڨ�����1R+I.��3<A�M�в���؀�ц~c��i������.��T��5�C?�C�D�?��x��O���;D��׮s����}�w�1�Z,���۝��c��)|��ݒ�%�~ۛ�<������g�d�d��L8�:�@�{<0)�t���7�q.�4���o0:}��l�x�=s@1�b���넑lfH�6HW:����u��^ ]�΋]��U)ҙ��;���,HR�޶'r�m9�jRr�ֹ�~�Rk+�(E{���&��ݤ?RN�$�i4w���9!&��n�(�٤����7Y�'MΛ�7�d�J6U�a��)f��b9}V#]?&{!^�����J��]6K�b�Efv�$������x%?)�J	4�E��>�0o2�����mG����Q�>�gm<��/��^���c%4���	�!0G����5a��:)�KT�Jv;�X��ώK^��,e�B�q��YJmQߑk�w�u��\9G�8�~�R&TB���hcAK���?�3?��o�����d�dxZ��517�H�\Ue͵M{��NO�ѹz�Mll����,��*�f�{�����d��>��s9�ݼ&?��]��u�Y�凒c���FM�! �ߜ�����ņ�,�z�-�>[
�E��I}�߲��78����i�������P/�7�G�>��M��Ɓ�0�� 1��Û�������s��R���혳Q�^}Ӗ(ć)a����O`�i%ݦ��7J��áB|�b*���`��@2�p��Z!{��� �~�O�,��;T�Jz/���ܣN�kl�$A�l�\?VӜJ�*[*�+�$�4�"��rk(�X'.�����`Ȝn�^����	%��Gl��U2:�[�}���ڼ6���=����l�ހs?Ǝ4Ҡ�j�E��|~�Vl\*��՟0gԍ(k���f]����+�����������5�������w\N4O}�S��dH"��P�k;��»�����e��TviM7���d�5��_�)�\��,]��^ �T�����.���H  �ȧ%|~�`x5��۳7�A(�o�q�Zͱ�3M lJ�S��7,S�?�40C;����?/�>L|�ʒ߲: t7e���1�MZi�����G� L�v�կ!,�Ҫ-����GGF��Z^���I$�FTE5�*�M�S'N��U2n�A�� ���F�m;T��=����(�$P�P��fHN/���n�@L��&6X�G�0j��kES�:Dxަ�G�_d�Q�B������ZT�}��z���VRU�en��ԯذHw� ���I��f ��r�D����b�R��iu��Z ���l�Bz�@����5 �W +j�ȳS��uT�:?6#Ć��5�8i��l*a��O#�j����io���4�D3��?��ϫX�����m�1�&�-7��mc�w�yQy�d��|�H/F�w�S1ʅ��л�&�4A�)f����c�ݫy��]#�40EK�9�3}g�
��&��I�ӡq���خdM����Fz0x��S}�<��b����VYMU6Э0:kUl[�)y�HY-����f��0g�!˦m6*+k%����	���tx��Π��*4[���2<�v�rvu�T���� T�k !̃$ݫ���ć�H�m��!
�8$��
��p� p����\�&�p\�B���=B�]b:���K��6�ޜd���� �տV13��7�1x�y����wP�IT�(�)����h#1(����j��o�Ѥ3@�=%��&�X��y��L���Sp�ڛ��J�+� �+(��M�ן��E#$BJ��8��YJ?��?:���?~iǎ�� �z>���nx-&��3�^�)3����Ͻ�9���DJ� H@��jb�m����ˎ�����]oԟ��^z�W����"�y�]eV5����TgB�~����M�����*������%�n�Cc�[��xQ��cf�ٙ&�fpl������R�k׆�OL��Щ���JjT�|80�d�ݸ�7�/K���2Q%�q�dV�q,�p$'�Tr���w�_��e�Q���Ƀ<�˗��f)��*�6 Г��C
bo�k������������{f����9-R�EORñ��^��4/9�0�i:�y��!S�|IvN��VԔ�.�u��r)�Y��EE
vh�c��oR�L�	U�՜l�8ϠM_��7^�g��7�B.­����G~�GF%�Ԯ�����)">��tsx���e��yfƝ���!N:M�9_`8��d0� �㽀��kJQ|�!�aq@.*P�ѐ��$�vub�nF��*{�6Ǚ�kfll�^a�ϙ�e/�|������� V����8�1���G���L�#I[' �s]d����jO������O��Y�)U�Ȁ��L9����p|�]�jL���۳f�y��h�$԰�0R � 5��x��Gs�da%����n �י!�g H���*�`�Z}���h�,�����|�u)ݖ�-�C*~8��u��t�lR���K���:W�+���W�,6;t�è*!����	/]]㯛�}���%��2��sù�ެ��ce�pX��VG�#���퍄���68���`퉤�-:�9}]S6�&%$�;~�'�'���=�����u��mb���R�*!3��������;���,�K��Nђ�\�-K����L��df�6g�*�e�0o>h�v�����k.ՄT ��#P�4QA �Cޜ���i�h����s�/٩Vۊ��$֜#3;��D�7�� ��Q�`���o���nvVޜVq�/�}Y����"�Y����{��9N�X��76j� ��ڙD���P�˰)������g�3E�	h���\�<!ur_Ԟd!B�
�BB5�?!�7��>��%gK��.j�a�H� �MK1�r*)����j�*� �2@{@IV��T�=y��F0�b=�)��<�S�xy.-m���*�Ji$�uC�g��~Q�
�Pa��H��8ό�.����=�5>�	LokU���J�Z/
]�Jt�6 �V�� VH��ߐv�Q��������¶JL��?�kv7t<����@}Tt��Y�\c�O֕�J0=I�[��T�����������5!g$9kҾI�ݮT<��/3d�����&��=���I��6��$a��X�w˴c��0�]�vE5������`�0g΁i:T {��5��;��Ь	��ՙ޷P:\��d������%'i��W�#����p��@;$�fTm���\ �,�[��8EXMmТ����t[�y�f����Qi{%�9�	}�4�9���1��ܕLP	�I+�|�z�z=�7�x���F���(D�;�y3���`{���v�\�$ߎИ�p���)�j*�Ζ�f��M��y�V��p�Z!��v���$Ă6�Kߚo2�<��6Ϸ��k%{�:4��������ƨ>1SF���+寜���y���0��E�[���\N�fI�y6�d��%���@����伩���ao^Ӕ�&k3�:K�<~(����r|���][�$�ީ�n�daF�%r�3�Δ���y|�s��z��5;�\�ޖ��d�q���c�f����(�Ù7	���k'&v�"�r��eC$��|��R�Gp;�dۭ��%�PoV[��>�kp��p�t�y>��$��}����`�+)����Ίc��젨L��M�Ѧ�f�?�3�7_�;y^����y�	8������ֺR��_�a�n&�1�Jj��g��'`,־�ܧ�C�z�ӕm�1^�VA����a�:7���h3E�ty�p����]���>c:����Dd7<#��˯��꿕dpN��o!	�X�f2��t�s���	�Ҷ����{��n�ٿ̤�\x(`|x��P���d��P�F\�^���7,jR��*�*�+�RY���4���Z��ԗ��f´a���sM����ڴ�j+υ�����5��׹N����ޜkI��AШ���1�g +�7��?�#�]�{�ʶ�s�TI�̽��dޝ�6Ki�h�W��%_ڰd�~3&!����B��j�8�D��7�h�g�cVkN�y����ľ��"%{�L6?oj^|�_�^u���ϣ�|pK�u{��>'�ա&�5ɮ���y�X��1�'��[H�)��qp�p����Y���2���~�=H�_���!�vM�}Z(�-��M�꼠�b�oӽ�TL2�!����4��WS��ŕ?���d���f�>?�&3P��'��*�<n?����0��+��!qu
��w�l��o����_�`�W:�[�Ɨ��ޯ�&��n[M�K��gjJ|y.� �wȽ�I�ˁp�C^��yk���gUae�"L�ߒ�z,3_�V-�;6תT��-�[�j �9�%�+"X�����;Gلa@�QrO�9��ϴk�U���L��5�^�?ӄ�����p��%�:8%t��{f�1t0���HA#KE��kMSB;��A�R�����й>K����A$�#�қ�ꡧi�2]V7{��'�zEw%!�P��ܦ`��y��Ǔ�������f���� [e�藥���k�Yf�QGT��uM��פ�?���Bܐ�e���M��� 6��󛠖����.t����������m���^̘s=6?�Ĭ�̪%3���~f� �"�s��n����T)���-U"�CI/�!.��&��[�H���C{�����F|��z��� ���C<��iҾ���c��62fxV=�s:�d�&��%d��7���%H{�h�c̅��s���g��'1x{r?���@4��.�	���Ì�du�%�ө�#��Yoh���@1ᰡj,��MYu��.Sd}\?^��>s~F��b><�}�V�.�c!�1:�ܰ����ܠ��JԽV�ۖg���_���d�gq2T%�j�#tebA	��0��]'���&�Rn�6���V�[���I�hT��:�J��.��y*��;қ�����|뭷�h¾S���&�&�bd��2@6��g�i`�,����5CȌ��s[����z�m�>co��}5=2M-љ���D��1��`�0.gq� ?X\���l�MxR4o*Y�[��D�_������gN	�]�@�u��1ߴa���=<W_�����t�f&�<3�^m7���~�4m�#���X��Z��7m�(O��]�4L՛0��A�k�����L'\cO����E}@�P��p�q�S;���I߸�s܎�A3M�4��7T��!��� �
5�5�LYu{JEz+KN N1��g�����Z���tk�D�6�~��k��Ṷ�C�	}�IsF���	G�3����5�=W�bV/]ەļ��Y��7�
�e�z�X ��AC�l��o:�Β6;	@V��Z~�&�����*��k���1G�m����F��ʚ��O��>�K�@;�c���z(��vz[El%L�y�`1~*`�@8��2��<n	��`0����4[`�ɘ�)-��&�7}��a��U�0/?���X}�E�$�͇�y��㴺����.ڤa�W����5_�5�T��W��_}��7�xJs�bh�C�E�*YF�Tb� ��y�ț~o�--e ����nˀ�7�9��Y�V+;��1"�� �J�<V���Z{�� v�ѹ/��d>�c���N��4��I 2]�bе���X=N�VW���}��4@�'�O{ ��D�1g�I�,�	��Z��4�3k���A+<�P�j ~�^���D���ϻi�,J|�� eI�Њ9���j� ���Tni�*b>�)��D�̉�������Q���	�w�:�&����藃����ω7�V�p��ت
UR��q�;`�J�S-�~~���+�DsJ�'5Qߦ]߭z0���b�#13l�A��L&IM�'/���ᅔb^���T �m|N ��9���6��`�K�]�dA���zŌ���R��d��G����E1�Ӛ�b4I��������9��o�{�������$�[��3�0k��̐2��qKK<Ȗ�2M���k`�T���6:�ڰ��w��#�A?���w��ӧt+�����֒���v�1��3d�.6"
��\�G�A���ӊi���ǝ%�5@G�.k	ɒy������a�M��zƅ��#�5���` ��c�W�^
���S=s^�^G��
��8��uF�Ƅ�Q}�ƥ�]�=���n��5v��F��cE���6ٲ��Y�BHj���h�h�Y�F"Kt��	M���v>��� -!�wM��H�3�T4��߯Ka/�(��ԥ/jq�������5a�(��̰���s��o2�^��8������惕A�L�^��Ƚ@��f�>��{1KK�
�qC�Y�XF��$���ĻXK�]����j0����gV�o��o�U���/����������"fz��Zkp���qq��$��)�F3���6��������0���^��l'3�8@y��Jb��x���	��`B�vt�׋	����c7~3E3xo �j�҂7�y̌��*kǶ1'�v�AK�V+���u�R	c�JG�
�6\���8�t�Tj	&?���ˌ=g�:��)쩶�F�f��B�(OU�J�lYM��5���8O��1�M�`��J�A�dy��0@7��E�՚�"�H� z�����7�P�A�5�Ro��|���Ο{O���B�,�a���"�w�5Ѓ�"�cZ@s޾�������w�g��*.?3m�df���S?盡d n2�&ò*�*L?x�����g��A���,r�=��.z��jΔ���2=З�S�ſ����_�ŏ�^��ݻ����߇�T�g21�OjYh������4�@��/wN/��@�4����ҍ�O��_3K����!�R9�8�ޙ@2Cd�R2�5ɲ�A����׈�g5����:�-۵��t���ċ����k�Mh*��ש���p_-����sgWH�:#U���@f/�9�g��t��7m1Z�������[��<y���`ـ2V�[$��G�$��F���}�A]�!V�3&;Ƹ�v|b���b'l��JE��k(�og׏�؏�HUvT��P�����sT�N��ߔ�2�]3������wB�1�6�����������l��D��}�^4�y��CȂg�n�����,�e�ʠ�cz���͕bfSn�~�p߯�ʯ������[@��ù]�[i�q3�&�<no��Rc��^t�g:M04�2p��c@��Bw>�J,���� �O�x!Q6��`����w�j�%ɬ��]��Ds2�Zr'֌&}�a�G�8S�XEkON�zc܀$�zm1�Yz��`l�}�|��"�Y�/ka��0��q��,7�		lt���~{Cm�Խ�"FS�7��|;a������h@?��k/�.��@��u��6M=���R��[Uj>��k�Ω��x��+��}\�s?�s���(=���ߠ�ئ�h�w���fF5S���2���>����~���y�^�����Y��w:���`.�΃�yg�KU�.o&r����>��н�6��#����������Ey���8ħ$�~������M9�w��M���w-d�i:���*3~�s�텉��0��X:o4�! ���3ڷ�8f~U��I���,Z�b�ms�~v��Z��v 4ۚ��� �x6WW���Yl̬���g�Ôk����v�ݛ�ޛ3��C?�e}W hjX�#܅���R9[C{U%i�[]͡/�i�k��Zz�:�e�=��ؠ*VX��Hb!���N����!�y�Y��3��כ]���F��Ц�������Z�A��>h���*�{Dv�/���K�	��U�mZJ�^�y�][~0�[���N7;v^4����=3�������������0v�)�j����m�|���:��Ҫ(��&��f㘽�t/�(<4}o�?� 
�����?�|饗v	��b�_+FH�Zl]ɖ�0&��{$��fI1��������\nsӔ�z�M{�9EYE�v:5�R@������<>~���n���Y��,.Ҧ�28��7�Y�
����*@��Y��ZT�8� !-�?��8@��Y���c	�(�����a�������|7�<��Q����!����z��j7��һC(��d��t�w��!��K��f%�^��) bn)]2G��rKx{�@-���J��;���p�R�z�{cS���q���3�������PU��6Z���Eu���nx�~��W2���6�C�Q=�wjr���Y��w��O��04��&���V�|�w]��&�d&��;�#tvr���U�����'�Gd�B��p���[��1%�{�����:���_�xJ�b�$�oU�w��!��,�1ߟqgIv��N�;�:��z�`lI�j?�L��Ѓ�*O�؄jԛK�#ٖ�Y�gNm����	 ������V�q_�3K��ۣ�eP"�Y�4��`;px�c��R��5|ڛ�`8a�,�����|d)ԉ��h �NG�s^H�ʆc���uL�#[�JS1_�CHa*f�y���; �\XS�u�ƈ<�Q�������(���.oP=_|��iG���:�Â�U�V��9���q�yv��<]7�Dh������/��/�����U��&��(�$�f�����x�C�iq�trSz�D��^�����$��)ھ��43S��d0��y������փD�i!4��G?:�O|�yiN�����Cjw�����Л�,����q����A?�yW���vZ�����l�+f�R��sf�����	��M����a� `����ղ��oX�I�q�&4��m�y�=3`�8@�~��Y��Dg50������8��k�s�`�����̜�`V��L^^=��0f�Б9b����ydĉ��M��J��u�Dw��d�OM�^x!�������0���X�P֍�4����ATTK�޼0�����X����~���
��7Ʈ��3#�4'��J������w��߽�]�����>��5�jb�Z��u�W
:3���f0�n��觳fzI�����X�a��~��{��]���*>�{4ǚ�*��1=����8�~������ |i��Ν;wK����0n�?Σi�m��@������sۆ�ڄ�94 p�����E��������ŅO�!4�i�jI"Ϗ�,38��ux�rl�����m{���$��~�Yǉ���u�����h/d�z��+��*@J	�^�B�pԚ��1�K�G�XJhǅ ����#�tUuY�E�W�)o�&[+��a'�y������1Ԕev�b�k9N/�1�����Q�l `�J��y睝|�!M�1жT(�g
5�b�]����-(��۴���hWVV[a8NU�l-	Zsa���D	�g�]:�~�i��a"��~���٣ ���P���wja<���h;�gu�d��_��wyg���c��l2V?X�B3I�'߫پ���/ Z�ɟ�Ҋb)�-Ec�G-�z�I}cU�]��&˶��42x�U�	�Z�g5w��2�|��KC���?��?�W�I��X�	��V���1�݌qX���i8�z��.�s��|��>��b[��l�*�/��&6.8k�� ����a` iay�%�(���b��A�K�P�`��.V���02 ƺ����{+Y�xe�{�Ri�Z�7CMGeҠəDYi���Y��N&����3C��
{�0W��Pi]��a@�}M���:�r
��$C�֤�5�N<�	�\�����3�d�H�]�@y����*��2ਐ��a�}T6�uU�z�"ђ�KK�`Ž/ P�zL���f�Ν�_T
�a�K�u}콝G}���#���E�ql��Nj��(�K��P4 А֨G�$���:FU{�
��+���BɶuF=��l,-c��=t�8E�ak0�- ��߷���{��+��z�V)��+-�o�	�M�=z��J;Yr�Ɠ����Ǽ�2]"6��QZ���<L6��c74w�n�mL5�ݦwr�3���>����Y���`ے_�Jumv����5Ь��*j�R �c�& K�y�����JewF;�#:N��ϩ��.ᮩh������N�����s:��#G�����t�u�*�!�������dӶW���~��8z���:����B�#X:r��통��Ҽ���b�E��jxX�y��H��bE����!U��C���[ �Ayi��+�g�E�P����p��Hv�mr��r��Ϊ�2T�jcpYҁ�r''�"���u�|sWdE!��S�y���Jf=�95r�sN��QU�P�FG�@3N��SQR��AI�l�X��7k��E�A���ܚ}�|�@��"��$�Q=?��=�N��7^�lTW��lݺ��n��$�$TxWb�z���[�;�(�����;���>�Y#���������|0$�5��@����P���Q}=�B���(�����j�>6Z<��<\�qH?j,S?��?6������fj�6KV�C���o�}C�j+����vQ4:����i��yJ�vX`��W^y崘�1���N�E��H6��4���B�*̒��һm�̬�]�����(����پUf�9hW��3~���ßv:j:�6�	$�ci���/�A<��c����umN��j����n;"����?����.��_֦���~@6�/s�Ւ�B,	����@��N�ka:��t�W(�7:9��d[�C-,�YE�unoP;`P*�Eo|�Fg��c�a^SV3:�'m�B:9)5)
�S)�B5�Z�{��p ��e��r/o�A�����S�J��K8��^4~&Q�bOQ��[��U� ��kkU�љj�F��[-W �D�LGoZ
-ʆ�{��dC��6�w��w:����;^��`�e��~0�voV����JЎ*^���{���~�4�1�9�+�&k��$ώ�Bζuf�#c�N>\?@��$�x�3�"o뾭��Tk�U����VL�~=�J|�&gyfp��Ԋ�x��n������\���g��T:36N3��m0��a� ������'6IK�|V����Q�q��xA��i�j��d�W��������9|ɳx�T�g�uw� |��o��q��J=��f6s��ϛ���_�kfI�kx  bۗաfx�b^v��CE�f��Ve6%X[L�z�os�%k�%W(���$ G��HR�%�P���m۶�}���K�Q�y�j�)��9�]��U��K �h]�ţ��8ot�oI��y�������e�X?��8' ПUJ��������j!�51�.Su���Αc���z)��'O�-�G>��M�6���E�C��=T�/�k�B�Y*�Xc=�1m ���M�=X�m���il�A֊�����qI�О�����9|��M���)������(}^��z ������=b����0#�t����c�3�y7h)13�&ö����N0.?Ȝ���S��@�{������f~011K�z���-��I �Ыj����[��јǗT��~�7�)�kc�E1�?����f�}BՕ ��4��h\鐼&�������������Y�q\��_�+ah0m�<q4AmCc���G'k�@�s�r�j�ɣ��B�U�7XH�s��I�V�@%����<>KU|� ��|� �3�=q���`� �8�.L9�t��Gh6q��1�Ӛ�j'����iJ݈���DrР#} �aכ�;R�wH
d�m�|S�;���6��N���c����: Iz-X�I2L�̣���zm��n���'��W��e>�U����AH�HS[w�"��On���I冊����?�O��=���ު���3zGܔ�������#��	F}t�]��^n����=�l����çU^�E�Q<]m�1����Aa"V]ю�&$d6{�����6��n��9�?y���G٧<�W�3����t��_��_;��3���ω_���6_�;h ����TVf�Wҏ^�z��>����;tw8 ��i�;�q�$3<���%���8����W ��3<\�@yc�t�Fq�) �~�N��G�!L5��js�;�#T���S��jV���1x�?�vh�q�V��	u��1�(���7u~�aIS���8�9*��|b7��g�ʩ��l]Yq��X�IзZC�Һ������?��S������D����;��<���:<�Px�"����+�_pz��Vy7����7;\ӵ���%�Y����2�3��u������k���=��v�B�����������ja���?��?��_�K�?K*8)F��_��s��$�֟��*�&(��q3�������R�d@������A9�e5��)�+���a=$�z0F���k�(1FIa�ۮ�vզ �<��=&��R[_���Gڽ�*����d?㟯s��;�������i1�&�e����b�w�q�3І{��� ��\�3o�,Mٮ�v��lf��$�M�m� �w� �m= =*;�s� |���������F�ꇳL���HJE���T���H��`�4�Z��R��y9X0��ٌ��1�巕+W��jP���5��^,��ԼRK�{]��MwN��7σ��pȤ��(��Q���⋝g�}�sT�~���t���������wݭ~o�o�����4��U�VY"��s;�.`>fI�tg.y��ܔ(M������Y}������݈���t�|�����??�7 4@˿�����x��uR���4�[5iz.J�`3=�����]>�	�y,~hf:�&6wj^�M�d�0���V���Q�;�_Sܥ�5j�	1���ض�
&�Cl5L�8^LE#���H��>��������������L1��g������=���N���Đ�ט7k<+l1�3ͯt>{$�ۺ�O6iHB|rsH�x.�c�$�e[�m5�p T mp��9Ʈ�f-b�R�,�-�����|U��F�.�9~��'�D($E�x�-Eeh��T�'g,�ʷ$J�v����/Kͨf�.�Yr��*���'�U��z����X���.�����H��Be�X�꧆���I�s���wz���C�Xy�1I�w�sZ�;jQ�D�J�p�����D��'��R��ͪP��f́���aʛ�@_�g�$@��Y%��g�n��iU����t�?�����>�EA]ÃZ\ߦ�u�� ���N�L'�z��_�i��<���&Z-��f0��,R�lo��&��:������y1�礶z[R�	1�%z�CEo�֟�/�y[Ծ~Z�uկ���j��w@�u����s� ��u�]�T�D�/����w���]�ј�U��	1����HVk:�;���h��w�����Cw�Q3q�'��TD[��h|��˛<�gɐc�ǩ��Dl��kz��GU�z-�G�<I���Xof!ը۶*���> ���nܴ1�_܇c�GۼN�M�'�#}�V��+W���~���ﾧ��W�
m(���A�H<P��x�zsg@�μEo��J���h�r��X ��Нg�y:����w�}�G;w��6�	fY][���3�.�����;���O$U��e��
֚����z�:L�����X�
������鍴?ݾ��+)"�j�}<����Q�@8���U��S�m����cZ��~T�:eu��1�Mf�?7k�������L�`�k��ܾ�mU���sX�v�������9*����v�O�Y�zǆ�
���Ù#������%1X�����R}_$��-1���t��u��;���_��Y��k��w���=�l4��ݣ����������(zc�X��3�13�ڵ�lK�Җ]�Ռ������n@��h�wq4)R��e�
�c--@�H�t)�2�l}Q̐�f���=�SF�	�����hA'l��48���ձV������B���D3�8r�X���!��(�ٽ'6xu"8�D ����I)z���H�^�-C=��R�Bs�^=v��o���<�y���߹�y��^��x�V���g����{��ڗX��@�+�-{z����:�O�	-�{�;{�k�kk�|����j�L��e��䄜Ev��S������Y�k�5�O�Ӛ���]�Ż�,}�E�]5N(�Q��L��%B�^sGf��Puv P��7��"�����އe'e�=_�����'~�G��s����޹M�S�%��3� _��+?��'mk&�Z�(����_��K�吘�&��61�-����[�<�b�O�튝�N^V�Yu�ޒ/^�����Z�\@ê13?��K����e�(ڳ�F�3Z�k��D��Ƀ�1���G<K�9�7�}�]��a�	�~ zМ��֖+a��iU㐲�G�r���B��T<*@B:�}ZI ��H.1wUښ�D�5NkUM��G�^Aꡇ����%��q�p�)�L<�w_�j� �ڷ^ς���(�JR��e�%F�c- �d��U=x�A��o�kț�P�G�����&�~ ���UV�J������^��{���;2f��N��4�_����(謁x�������z����;�}�x�����c�AP}8- ;�����g�����r����������������i1��=�zgT�?�#?:��0��n⛿��ٖ�!���#���E�A3 >'��Y?`?��)9��jHo�����&@aU���i�u�챙Ui��p�rer�g���v��fЌ�q�"A�b�"|��89����^� S�J-����Æ�	�	����$����Cil�r��P+s���K�;���'<a��� er)�*׏(� 1{C5��z.=���M�� � Cer�)h�J��#�T�X��b����|g�c��ZL<@z�Ub���UM��̇�Xe��7
�����A�1�2 ��zm�Wj3bm��B����@�S��:�������_�k�b�g䲍4�z0��1�)������c��wS�C� g)���H��Mƙ�����ҧ���v����N��!]�����\�����R9Q@y� �'����_���T�ӧ>��5gs���A1�g�,�\of^y������J�5��r8��=n~g-8�ުI����б��	U!���yfp�͵֠�Ѓ�P��Y�3����I�UU���k�#���)NV���k�s��EJ��֐&csWu	�YK���qI"*ٍ�T��7i�:�#G�w���/(�X	5Y�j�T��`�R�p��5�ۙ�#ӂ�m�F����l+�	�������Q'O��"���2����.H4&��jqK����9f�K�/������y�X�ʝ�k$q��P]� ��V5:��u���'����㓒Nj�yD�Ú�[��[��y'ɢ������<��>��Tr�,�w�e����8O������zc|QA����<�c?�c�f���S7��ϊ�{D۳�}�^s7�:���sndF捘C ��t�Mf^\8:������w$E��,S�O@��w�G�ig)KV��X�4{����\���-��l����.�έ-�E1�#�
iU&m��V��t��ޮ�Lx����Fn�}o�Ｄ����������Gu
�Pr��"��ymnbB���b��0e�P��.k��Ib3A���E�|�ZEIl��j�jw�tMU��̓,��i+׳)0�{S�q�ڭN��������Z`X;%����d|�����ol��F�Cm�������iU�WN�KZ����������	OS6��hw�1�Uv~�CĢ����p�×t�Y�� i��=�YMa	Ӫ
�λ ���~]���}A��g�&f��O��O��e��p͉�2�\�3oN�,���<��;ߒ�A�50 F0��a� ����$cr6&�ҡc���X�5�&�a�9���MVa�EEk{9 �Z4� ��!V7��T&p�"�L�oH߻��J׬�{�q���;%�4����N=�?*�K�Z����ӛ�ù�|�ݳ���6��E���
UР�D�*�f/ը�Ϊ���D�8Vr��f��Q*^�VF��
F�e2�+��m\R�T�@2,����'���"u��K;9A{�>���|���<���ot�͢�ݎy�MD�v[�WVi�5�us��zݫM�}�rП����W�R��{��т�SZH_���ftɰ�hlO�.-��g�Jc���3#�NZ�-��11�=j�Ry���/�I�P8Ȍԟ���e�EsU����^j��d�ϪƬu��=��g}9L��m|:ȝ�r�!��u�h9J&�4���S�YR�$�5��Z��fv������Z�Jǎ��ox���rN� 8�ɦ ����2F�E�ľ�oǘ�;c!�1/��zR�	>�#�T� 
��w]<��H|�JHI�lI�u#�P���MC����F_��~;T�cs���c������x�q�5]nàh��8��T�aK���ul^�R�D8��2�S,Q�P���%���z���v:_�cs���C�w�^@<���{��߬��A֌����Q��o{)W$�?Cx�x[6���ie:�4�jN�j��t��]��yϼ#��Y9��� �אm9 ����iU��M���|��p���0*�"�0�����/��E�܎��Y��y� 	G��Z��N3�e;x�:G�Mi��T��[�B��~&�V�iH��۩�֬^y8�څ��C
�8y�X�.���m��u��+���PZ`J0=6L�H��lS�W�����]�H���)��/��f:vS�*њ�N�i�����te<lH���jըA�&f��ͼy�M=Y:��&�3�lHϪ:���go~�jK
�>$u駞����~�b�Q�Bɪ��p�P��I-2(�V���4��9{[���Ř>�]�S2����9\��A�� �M��\�ր�k��D�3ۛ`�^G��ժN�g'K��3ڀ)~�����=����'�=8�'�;=��1���,#R���OֲcY�a�R_O+şc՜��rn�K,%Ь��S�Z-�r|��<Q����YM2�5z�J�oj�m�vsgH/���3��⳥@0����`ى���`��R�=I�7��;5�)m$�
�WI5�E$ҎRL�4�l�+��b�-i��e��%Kms��jPox(��0"������yYr�A�������h%¹��ڗ�1ř}Z�tQ;�Q-���t�E�,�RZ-�����]VV+X
���sB�S\�O�8U^�}� x9��* < ��UMZ=�^(� ��*͙�Z��2����cTp��w��n[�m�N�mfg�%/��2��6k�km��:ls$�^�n��f}7$��K�ZM	%I���#(���?A�J%�qIEb�eK�M'3���i!1���� ~w�7>��I�6I��S�OE�C�J����t����Qf�<K��T%~�j��1���U��2�{��:�%�ڠ�\w��X$����_��!
ޤ�u�q�B=z�p��T��o	6�,�,((��Kb&��/)�?H �]�1֪�
�0�g^�'�xRyl�tE~#;��^Vs�F�I����*�Ro�P��X��|J\m�.�Uc�kR�,���휢�#�%�}ZY*N�1��M�mz��\��+�	yG�ݻ�����Ppp��e��5��i�}�ޟ��o���k@���)��,�͠k��׊�9;A4�i�k���������m{�q�C4Lo[�5v�Y.ɊJ�ΰ�=����]=C��b�+����9�F+���=��9g�C��]8	�vK*D9���gN��Ҍs��m���ȩ�qݏ�}�� ��<�4o!%9|a���2��]��pv	�D��A�|�w�<�p5A�ǎ���sϽ��L�Z<of�z� <`#"#�q��p2��)~*�&h�Z\}BE]զ^S$#�T�C�ӿ�4�j���<�������Z����d�W;��pf3�p������?�S?�y���A���w���i�J(\�f �������3:~L��z�Y�r}I��9��S �QI��}�R����-;Ra�3*K�s�+����V�:a��e��(B@�f�E[��s8��`3�����C�(��a�+ey`ެm<0����g�N�
��1ۤ`>��0�eZZ���&��'@-��2\{��K�;V��݊]�p�R����[��B�a%�&�)թ�L���}L���,�"[!��쓄C�L��ٸ��c��w�z���Ït֪��
��t�Q�]�Z ,�;�^̱�V#��y�P��Nc.b�*������iq"w�2$A�4l�q��.���Y���s�yE[���!�q`^6�j��%<��G�W�%U;?��CR��Y-�G�(V�!���H��؋�������pP��eb��p>%�ɛ���Iu��u)P%Ai���nգ�u��fI
�� u k��<;D�y�>���ʞ�ӎcm�|�e�N_\��pRQ!ۢ�]"�q_��Hi���q��Vg�3�#��B�@b��h�Q�Q9�u�1s�5��:uR�����,-��Y��Vtn�|sdpU�0��Y&$S]���	Ÿ�)I�9��'�~l3�{j��"�]���I��?$��R�.�
��W^y���t����巗 �����TzN���Ӯ*�$Gp��T��k��8��8"a[݉� �1�?�Kl�Q��<-���wٔ�{���V݆ZOs^���+[E3����(�o�<J�B�2���&�1-��?â��Իa1�Q'H�u��� U�W%����1UB��Y�Qoۋf@�K�V0M;?Y��A�S^�A��XX
\��3鏵�3Ъ������F�h��Ϝ�������$�. c 6�ZD}f�^W'J[0K;�H�>pd!��Rŀ_Μ��xB��p>�^�wZR$ �\�Y��8D�
$��K�5���`
7R�ڇ'wm���.��~�	��v O�C,.�<��"�Y�cN�D�T������[��k��3��d��H�lCR��K�H9&�Z$��z�Kc�ˉ�v8����2�t��BTʱ1:_$��X�>�BF�9�D�CI�5����\��,�k�y��W�����SqJ߯�����i�������ZgF�K:)������}V*�7~G�p]$����W�5o������l�iI��q�k،�mf�cn#ɀd)�4hv�qBk��S��zK^fXv�w8Ҙ�K>8{�G�I}��� 0^%k
�鋍Ό֪����dL�����C�SŬ�$��t��H'��}�>�JJ}����C��}�Rۼ��
�X�a}0�#��~���Ή�'D��Z!�g���pNc���_���Q���^v��^�ٝ�"�uc��0�\I�]��J�E�-OH�цf���@{ɀ�D� �/�v?)0E�|	�V �9��rxM$��1�2��U��=�8B�[��|�*g�wۖ��~r���6&��ı
�8p���C�s��~+�Í���(=$��Oi��
�e;�2=�[�pVh�Pb�vJ_҂���w���{��w����o^��zo��`*2��Y�I> ���g���-����cW]p�p�!mٶ��GU	��Qڳ��8��T�8��E'O�`���/�c�ߩ�6#�����vBj���ǆ�P�p!��b�E�]�Յ纙H�mw�B�7�!�ޜC�O��Qw��-0aW�x��:�=�X8��t���駟'�իGnU�%~R���GV�ML� W\2>h���%K��ƒ�y9������b�w�޻?j#���f���f�u�d�)�frla����PsM<v� �1��.��oX���c�x����l?�	 o�h۴�^/�����0�$Q�g�2��8�U_�U�$e��W��A�)�8��`��n�����MZpz�W��0�d<��?��%=�Z����#f��~2�M5��f&M�0K���!m8g#�a�"�ƛ߲=e���qܘ3̸<LF淥v���(9ǒe�,o� �[�ձ�9��.��b���l�HH���"j9�ݩmȧc�� ��5V�`IJ1�uP}��AHs����;��Qp}�#��������v����1�B�o�ܹ3�ZX�g'�K6*e4�����Q��Q VY�OK��Z��m�{۹kG��w�F!��k�I�@vE��JC�UxMLHb�\�iI��N�p�愀���R��zCo������w0�im��.�=v�l�˻���e�Ӥ�T��×*!����:���'#vR����?<�{�˦�©��<������A������b��I���i�7�m*��!�n.Yj����Ҡ�,j�U���� A���7@λx���N4�'�u8��9��9�����p���:qU�ۅ��5%K��-��C���%�Kxr�8�06�Zp�̈<'K:A��;�>�OI&�A��֐�\1�e�N*,���o��G�(en����W�n�J��aɘ���kC�ų�q91R�_��$@�.�wM��ɀ�y�:U��ߡ'�;$i���_��!E�P&�JL���N�(�F�9�\���M��¦W��Ü��k� �6,��4�V����DqNZ"53�c�^�����u�R�ɦ�$H���x���G�W_}-$n,��&��q��i�i^<�[ �#��y?��?�y�e{�Y���	�F/��df׏d8��w�f`��ˏ�ax0~^V1r��x�N�f qF~wE	�7��ҧ3���21�ի%����BI��T?�@q�9�X֮[tW���Ҥ�S=j�e*	H���\�)l�ʇ�*�
Ć��`Q�d�d?Y��,vQ�-@l�y��|Q�2��jc�*c��W�C#℘�h-��t�J9�lV�»:<�`���;2A�}��d�C�|��;$��|��"�~C*�������N���e?��zh.�,��0�p9vRRܫ/���:+�n���I�뼜�����<62*5/jO�P�R!������!��A�U	)�"�4��Y�Z�� *lѓ�~��e+��q�vHE�c\�va$~�+��b�ś�lL�m�x�� �0���ڣp�ݑN�(�/Z��D�Sz�a5����n4
��K�*������V��s��U������`\�ΛyH9����>�Uu�o'`��K��b���� �/�%�СHa�I�|)5�L'%����H�l�FG��SL�k�����v�Ƈ����7;�}��۫:�������B���޺u[[ ��w��Fڸ;U�wP�ek ��]E}Q��r�'f}V@-�X�zJ^b�g���؄��f�vw�d�!w�_q����Q`�AI{�;[n��ټi�򡮗#ЖΘ��Ȏs�ęn���U+�������i!=��y�.��!��4�ջxQ$PU�#Yn#�u�fG]JB,@@c����y BԠ{�hc"�5s�zSt�Fu�iI��bj��J8O{mK�� ��0s����q:���( ��A��Ź�Ȋ-o"�&�Z�����h�%m�oK�x<�r��״H �K����:)��[�� oU/}�-�O���\K�5<+��)|b���g�}61`�������;+@����w�}�8�l8����b� os��)�7�K#T����F� uHOI0����2O��/K�,�pQ?:|$��|@�x��^�;f!����ȩʘ�g�_o��n�Z�`Jz��A��s��I�@5�^�J��4hT�v�Q�� ?擵F�Yr��ڵ���/(��s�=��B�޴�X����p\*�S�l�e�Z.�R�Z���/���k0)3OK�f�Y�]��Q@)�7m�r9$3w�F�w��u�m��#�[/��Әu� &�ڣ>Ux�h�Yq��n/�v8� mr��x�����b�oJٵs����P ���;J�e_���|8b"�#BG
��/���)@�?q�d�)$�r��<Ӈ6&�1�u��9j��VW0��R����v�_��ڻ( <-������~�v͆���b����#�ET�p\kV�{�D��P��Q��#2휕���a-��c����oy��P��>��Ϫ�_���v2}��1I�紾Ƶ��s����������-zP���K�,)ͅ�h�u\���X�+��m�fI��Q�av�!\��ͩˬ*u��.g)�6.��_�"��֎.p-����P�IE�M���K�<T
�6 A�K{����9��dxL�A�L�j�������QH�y{$G�Z�H���j8�Ԅ��[� ���p�9}Z*H����%�Kԣ]0��s H^N}��d`��_2�X�F������(�R�y��){ꪠ1���W0�<7Cz��h`��h�����h����ܒq�XO��W,��cR�?�@ި@Ylp�C�T�v��k���/Qi>��a����e
TF6¦-(K	ӽ����9$Ì��$�3�F�t���Ϭuߜ�����*8���-%��HM��� 1K���C�Ch�D�
{����*[q�)Yi B�}��~I��ā*t�~�*P��7�@�'�M$�[Uw�&�c�",*@�����a��*`R�������[��!�ª��+�Q���KkS��<OX���Ѧc6pBR�8mP7�C�ʇJ����7P�sϽ�t]�]Z���u-v��ǚ��}��(� }�F�v@s�jtT�Og4g
�ǡ d0��eJ�GR� �_��7�c.�\�[~���ٓ]/g���.ѺX�ϩu��}�z���,�m��@�a#Ի��m��L(�U��>3S�mu2[��%�P�� ����Q*G���t��1Tq�^l>%`>5۶��3<\���x��q��"�$� 8��M8��7�%�6M���1 �v�U�P�|�uUaۍb��1Bj֕�ɏZR����7
y��?�+l�����9���wV�s�"gj��ٱcG��)D����X�>����k����@9ix���o���h������`�"N(���K�c�.-E�YGK�juk�$�rr64�)�E�$o⒇tB���t����A4����kZ �P�i-��@�@��V���?�W4��xj�ç�� �� �RRn�;܂k�!�'`��P"Z���"�������+/�;����K�;�K����l񲮧���GZ5�x�� �vOV��Rqk���v�m�ʤ�ļ!� ��c���Թ�`�^�X�;�9�X�x≐n���)�67�}7��Z�g���R��K�ޘ�!`3��п��s�^B�*l�5�q��t�&m��Y����%�"�xU�ʃ	y� !)�s<M	�G"�u�v#A��a t,��C�e��[Wl�H��uu�9�sƴa��p�>��9��Y b�DK�Lv�b(�
g�2�$B����c��9��	��㱽Ȓ�U���m0_����t�~5M[��j1VK}H0\k�	����x��u��-*��i뾇�PӅ�0�'�|��/|!bi���������#(��͒
 :���%��F% �{^ql1S�4P�:(?T�c�
	(��%%��lol<W��IO�,^T�U�*�1�pUmYp�dS��
���qƺQ'�Cc�W�q��]�ħ�%!��"�f�橔����!$�З&��髁�ر�c�H��o������Y{�i��CH�Z ��۶w�S��t��_r"Xu���j�&��x9)��Ss�2ڶ������v瀞���@���!�J&�jv����f�\�ߨM�����s���_��>����R$� %ѓ@x�o�>��7�I|O|�Wt���<��'�)�!�GGG��i��3��b�����D�\���}��T��|  ��C�SJ�r�K],�� ӝX�����j�v���uA^��R8Ȭ\!@�"���w����~B��w�ڻ��?���4q�w	ؐ�Ǖ�ༀ�[�T֮	gI�'�6vA�c5�rDZ2,0�t�|�Z%�b�5I~@���/=֪6.a��@��Y�aJNZ��2�VĆ��l��\���XW5M�9��y	�h���g�-�U5

Nj��̗����`����圬r��f[�ǅfJCf���2��5h�~`�0a'�Ւ6|̊�ap�H�������0<��:�;� |W��S
��	8�. ¹ 1��6l���.����*Kt�$�m�n����ߦ�ȡ9�K�aM6�y�є�Kx�`�`�=��� Գv&�����2Q~��d+��d��^s@X��������{"�a�{��W;kdS���;�Ȇ�i���"�NI��ӑ��FHy�=/ jN��4�j�������qp�am�C��o���0�Fβ�'ֳאm��Tbux�2�����Z 9%�Q8Ȝ�!4�[�p.8a��NeP�v�����w,�\�3�$�e���(�]���9,���|w�Ⳋ̶A����|O�4a��ZM�rMa�J�U�a�(��Y�J߭*œ����N���W�hH+_��_��0a��䗬7x<
���F�(MG$�^/��-oB.=�b�R`�|�K_
�%]����c��;o`,�v���L^+ݟ�˽�&l��M��ۑ�U����O}:*L3�ڸ�KJ��r�5�����)`\ƆB��UP��c�͘W���z��q���%��4��	j*:�^��o��o�a5z8ਝb'\s���B�q�g�7:'m��R K��ﯮ�QS%j���S���3�^��t��9~�����e��+,�ޮ,#�ק�I-��_~�W)��e/B�jm��0�M�`�� ii�Ra�a�*N%zČ�G��E�4Q�~�g��E"l����=Gl�d�U�qr�_��a�$?)��H���4��'�f�ĥ����Z��SG��f��5~l8Q�fș$�f0"	��@s�k�r�v���&��M�������̹Ê#8�T�4��7�ِ���EE��;�x���] �La)��XV��6o���~�D	I�Z�LC��#��3��Z�p�(���F� �yч���pM�WVu�Ȭ2m��*�w�(��J6��|w�5{���(��e�=v��0���2����R^K������Gj���zK8O�����&�'g�ٶ���I�B*��s�H�&�1�B���������|wxZw��P�z"����0;�H��	�����y�0�t�m�.�b��tsuN�fJ���.�b~���d��y��u;,ZPu�8�)�ɧj�Y�Z�X�/�"�3��UX��%^P�Ru ��c+`w&$�[n����v�.��M�Cs�'1�w<�����(E�z�i�%8s^-���[�p�ר���|'Si������&�`R�a��alfn0����MaSs���ބ��R�SgY�w���A%Lԡ�C�|��#;���d,Y���]���3��7v:p�z���G��q=�LGKhY:ݕ�8R�=Dx��%�����m��w���W�P�g��� �$�6�&���X�R�Q�&sJ �w�~�����Y � q��\FM�����Pk 'FH�b�,&�p0�>�=i��\ݲus�;�uE�g�a]��A�͛ �M7m��ޘ�V�jc��e�s2��[ �	��kZ
LM�K���$x95���^��	��ա\e۠�Y`P�,�qۮ�j��,2�La����'q�w��=i��Fg��]
�س�6�$e碜��ިx����h��i|"� @ e`�k�i��T�`y�}���$@�t�ˑލ���O��^hp�1r?&�s�Ʃ/��E�R��CM�''je��N1H��m��q������Zє*�æ'�P��"<>�5Z6#�]�Fk�ԅ�P�����.�a�쩓�*l����������I��~��N��yVۧE�y+E��r����
ԝzI+i����ΜM�~䂬��\��eu ���ۑk8Ʈ�	�]��Y��t�ka����5���mO���R\�^`ǚ!IC�Eڠ�=\�!G6�1����y���H�V�"W)�N����h?�F�f���14#�[�
K�7T���[�vuT�h�}���g�t�j�C8Q����ӛ
����\#���E�E:6%�>~�����O�!���=��c�u
9�\ۈ�J�*�����+Z��$�iyQ��o�Y���^�fU�����b�$=�)�r�@\�j�UߐP�)��Y����o~������m-zQ Ԣ~͗DX��%�'jF �vK���l�s��������.p�j�jV;�X}U �xҮ*�;�"Tn�=Ǖq�]�S���1�P�,�}yq]��N��%�E��' �ʏ7ޛ0]�OFQk#U�t�Ŧ:y��˦��О��L��Wʗ�����EJ�	��1��3�e�d������ӰE܆�jǞ���XJ���
0���&�1�)����0�*m1�pF:o�VxP�� �
�.]�9�׫`�j�GTnI 6����5�����d��u�x�D�P*~0��}X��F��@#6,��a1�@I����MWu2���[��R��@e���S�%�̌�����Y¤ �U�X3�	�rua�:q�����lϣ}�/�a@�
�h9��ds 4�58�f��U�H����lp�@�-� �H�+���Œz��F�\�}Q�. �\�q0X$C���~��`���Y�TBD�jF$�H�-�U�RN����ӧO���ޠUb馑c̨�V�y>�o�E��#8���#F?H��*���c�R�AX��H$*�7�ɬ�7!%�u'�^������S{��g�2_��@Jw�6e�[�T�urcKG ����[��泝���R��+0$�����E����t4([�H$A�,U��b�
ea�,��膍�;������0b9�$h�����Ȯ
5�b���`b=i�Y��`T��i]{Ts�f����`���ى�I�,��zI)N�̯7Y/͗	X *06,��_0��U�#�|8�k�nu�c�αg����O@�#��"չ��=Q�jP���W�YR·~r,��vH~ e� �d���y�"I�����\+�<��s���#���7*�-����jJީs�_[�l�d�)�1q��RQXמ�����ެT|����"+�^��Y[��Θ=K�5{�7M��e��(R��xD���@.`y�M�4�D�&��$<@�v��=w�#`W�&Ңi��;�Q3��ъ�F�K�'���#l����W쁫�&]�n��%�m�2]$Y/���yG�8��Ҝѱ�Fx��v��>J4X�ϒ�w�������;܎�ʜ���^�h��P���(ci� �S�YgU�S�e�O{v�'{ir�U�0jK����PΧx�����}�,% o�hu&����\�VBq����!�|�s��k�����I��;�oE�X���)2���� ��СL{ٲb�d�Y��Q�X��X):,u"�������*���={vwN�7r~�HhR�{��$ �;埤����P��$��Y���5@NP�Y �ތ�怤�U�W*1�xM�^BKVI"\�~�b�d��vKH���9x��C����G<߭����=�g��Y3@jZ��NW !N1Ќ�O���[�tn-�92��y�P ݎ+�)�i�NLR�	����{U�:2�l���'��{���W7�0X��\��{�{�d�ٴE���
S.N�D�1��#U� �l�|�;pmW��r��ը���:O�)��o�m�CK?�H�81��,n�(�}�{�5e�lE�X<A�cm�tx�� ��>ܹ�q�+ (;6[�Rb�E�A��D�A��^Б�!E�S�>��x�*��2�xl8� ��L)�M���*]t�jb�LZ+�W
��j,�8T���D������[)}g.�1	�ԛ$����*���2s�R�.`��������͛�wn�U���MU9�gi�k����/�I̹��?��*%/_���-��vf��끂� �����tM����ÇMX3H�K˻��}x�z��K���:���P?N�'�h�p>����F� ��.��%�MM�Kw��p����$� �I��xxJ�Pl��P����N��5xF�I���� ǹ�Dcp���_��\A�0J>fv�Y+� B�.� yY}
���txL0${
`M%T��>�l��.���)�����D��GZ y�_�NmoU �<�i!cEr$X�U��$D@́�HEH��	h�Ɔ {��8jP6+�����4�Yq)ҲU��|B
���H��2YfHW�"�[�(�W�k�82�p��ݼm�JUm�l�����d�D�c#����
F*;b5s�!�̗-���eo�X���^ccJ鶜����ܤ�!$Xт�����H z\�O�q�ҫ�Z ���g��.�7FS���D��t��|{��J��TnQw���xq��5apf��*I�͹B�nU�=D�0�A�}�=�����p�Wۓ �cz�ds�K��Aaݚ��!L�k���pL �0�&�XYQ<"��°�4>�DC;V���rB��%�Z�9q�P� ��K/�26�y��DP���e]�6����U� 5�P{�.�! )P,������j�Ssmg�Q9	�B5��0�7l�j�;ﺳ�U��n�n�F��)a�� =ۄ� �jy�*�\��#R���ހ�Є����O��-6O�H �[�jU���5�W׍h�[�O��<�Z �'B����(0�#?��v8CH� �i�\��*v�?��j�(��}s�4� �9�7mr�"��J8��\F��͞��ñ���x��H��#q~�x��O�-hOU���@ �����v�
���)����;jMW�@�� �r���x�2y5z'T��M� (R�k��. y��r^+�Î�n�x���S֬�ady��ޱ� _@��j��\g)^��F���'t� �D2ģtp�T�Ҁ4�+�D�V��c+�t�D�kkI�7�T%�{�7�6ω�C�+�Y���&t��b�z�nB �ݜ��Hs�-�1���4لJQJO-
��2er�&'g�٦ډ ����c�J��M��~7zJ�}�ҩU�Mj�.Lk"]��ȉ�[���d{�noJ����� �*�H����!�s,A �H	��`-�����2<$�Oe�9�7�*F�3GF�e�"#�T�K�������ƽ���zb��R���@$��

+W�]��ݬ'�����w �Q��I�?��!"H>l��-!"�KY$����F�@E]��ëwXjK2�C7tF]�GR���=�*�@�X���$��Q�'���n��#Q�p���ѹG�N�r���ڦ:��;C�76��	un����!�H9�S��THwo���W|�W���jϕR��Q��CGK���ȑC����]�|0��U�Vt��p�Ȏ�ڗ��)���|s�V"�o����(0�jt�o �z�JBB�s�ki��:Y�.<���O'�@-F�{�X��SHX5(��=�Jp4�A�gǜ|oK�����E�s	/ Ӡn�}�@�V	')6@��7����~��n�~���.��mQb�7��{���ݎ˦������'���>�~Y��s�%U�R�w%��[K�� 
F?*OK^���ëR�RT���#d.�oW �m�#����;��{_�>�B�H&c��Z �^~����/��SԠ��&��  g#�+`��̧7 ���j��C�H��&���wG��Eڀ<�yGR������u�n�)l��c� }U�����k/��>���ἒ���D��UFl_�`�5�mCM�����!
%.NJ9���X��*2����{H��0s��k���YMj��%RO�,�+�AƏt��<�D���L5�"`���'`��z�W*�q]HVQ�W$�9�%��7's�>Po�"�6�%^�7-�_!U��C��� & �ԷO� !�p?�L�eˊ��7x��.�-��L;wA���K̅ru�|kV��lް\�F�:d�4q�R]
(�� �����k��3�7:Ū���=�~H�|��֛"�}�*t`oMN=�@���%�KO_������y
�WKj[%:S&���7v�d�l��{��<��:���;�<�P��W�+I��տ����}�ޣ�&�-�sl����@�<�:]4�}�km����Z+�6��l�����P�WM"��5t���,�����t욏�;�#D&�Z {�Z�i� l1Nη`ؾhγ�L��v��������N2�Ri�^�Ǐ��8VO�#:���I��bq��^�: ��U� (@Dj4T�Td8%��!��O@���{<����hpg)*!���JT�	��C�'<G����y��';�Q�w���ȵ���S:PՍv��~�'xԼ�+y�q� ���:���=Gώ}Pkb��v���١|���)�Zݤ���L#�5�F�) 66$1 G��v�Yl��yD��f�rx���tux��-�Gi�]|V��'�wϼ=���@x�(���z�����>�lS�Ė�P�謾�q�UĂU/Hڻ���4K�v��1��^m�A�43��;{��Ӭ!��FJ����Lۜ��K�7��v�֌�۳�Ҧ�w����D:$v��?��RJ ��H��7,�`����gu1�(���<���ٱ�Bƕ��<�c#J���p���h�z�':o�zC�R�aH��9���r�>�m+�M� �RN�U�z�t{P�.�3?@�1�7���y.��ތ�G眍XM��C@/]~?��ب�w��+<S�@��͝�y$�s�FL�Aߐ�m3ER�Z�:�y���{�"z�[������yM{EK��(p�$Bg_qm@;�X�sǭ������2�rP{�`v�w�P�<ǝy�a|��9t�@h������ʡ%v�T�G��6l��^F��h���$l/�3KH)x\�Q�pz9��/��)�P�:� <�w)E+��A������K�})�jՈ��SLx���ݻ�Dڳ��7j����'��sC��g�����®H�69�l�iKH�H��4��	�;m���^�vwIܹC*�7��. �����c�U�I㰤��}_􏵁'뒚,}��3l�H����
�o��ڀ8sè�]�
��e�>�Fl� ��ӓ��ޫ�j�𪑾���J�ff��8s\��h��5��ܦ���7�Y	�.��0d�Ns�u��ޒK�q袽�M$K3�p��1bw��rVڇ1�{[
�"!�����df9ۍ�;#g����9H�?�I �k��"G$9���G���'~��R��M�A�����d����<�z�ԙ�$s<��X�ƥ��l&#0 z��Ӗ�0^�T}9,��?��OF�Ěu_)����*'�g�y����B"D�{ۭ�u�����*@н��;�ۧܨ�J}If��^{��O�NT�cj��k�(df�%Te$ք����*�EW��!H���������|���C�t�u_�u�~����o���e�.������^Ӛ��vU��yj��z����t���>�+�U]|:4�^�|Z�u��-$��KL��[����� �9Gh��j}A�48p/�ۻ��\Gߜ��l�Q�%��^��s��a���.���9��|�@��q\����4������D�G; "*F�cI�4m�!�T�<#y{����a;D�q�o��?l����O^��ڈ��w�5�d���8�`�<���l.����=r4����-o��
�`�܇�x�"}�(��Z��MŋCŽ�|���ջ54�˖̀�ڒ�3�ؾ	-c�Z��A�]��=u�6W�u+`
�Q7c��ʯ�ʐ��� z���%����ּR[�8�]�30��[ �	��kZ
\�b  `$�4��/0�bp�d�m�/�ؐT�W��oU���<����a�A�"O�V{:u���\�W�5_U��>s��SC���;�Nµ�1F���r������i�>��]=*��곃��\;z82�j�*�{OJ�'ԁ�ڐ�To�ת��ތX:F��bȦ
F����x\Z�L�V��I�Fqz�6m�Q�IQV��9��� �V؀E�𨍊��q�� ��RꉾY]n$/���(�f z���T� I��Z4٪b�<qB"v��lL�dX�:��А������K���*Q�����e
��^�;�@g��6gF�|$����s"�CE��Y	3t%��=J�Vt�^�f)`Ab�Z��d� ��� ��/���k^.s�wg�9���%r�>���HC��&X��� ]r��tfEBEu\�E-�@�c��[�����L��#"������)��M�U��.J-	X�BU�Eg� �oڰ>����F#�(����m
c ��^��K/+��s�M�U�%��j�b
ȶW��H�*�+�&�P����~X��x�LĦ-ja�B��@$C���̒ǫ%j�_��r��U���C�P�tyAS�r����s�3�ɼ���3��|q��>7��#Ro���)���ߕ�	�p���`T�{�1�6��L�+)����*L��w �v@W �lC\ʉ�]�k��W�K��
[%�Wl*P<��myV���=`�#�;�&�2OHoH"N���\�)����AFQY��/�D4���� �}�;��J�J��1i�66hl���6tz$OA��/UʱU�\#�X�mUg��Mx�>{(`[�bL�Ua��Y孷v�wh���0I��H��%��@�$A~�����ZH��g6d
���rB�CI�PI]-Z!I��_��TsRs�Kj�]� �\盾�.Y�d��^��Ȁ�u��5�E�T�}�=���t( �^L}LLJ<���2cDJ�-P4�6\r�����<Pՙ1¤.a�n��W�䄄��({Hrpr �vl[DB��HV���ĻuU�:� af�o\�$�nu\�n���i�K�����NC؇�A�b3-�j����u�ٮ�ػQ� !�&�I@��H�N�]��m�\�;���C��N��dGl�Zy9>*Iz�:k�r1ށ�;�TC����9+@Z�0
�RԌ$�&[*P�[ !�f���2]3&U2`v^�E-�'�?�l �b����!��U���(�IB����ț�O��UR�=r��`y�J�c�}Ocy/Y�,%�%�~�_-^�	ho]R���!���(���>���T(����Z�6TgNf;y�w'�vm$4���_�(P�!�q/Kk�C�ګ#�s�"���H��o�����J(tN`b��C������!i�R��w��,���[j�G���@�<�g�=���	�M\�0K��CQ?��b�*�~J^���B��ܡ�x��l��/��#5��ӛ;��e���#���K����Έ�M������l�;��YzS�y ��f,�Yҟu_�k+�T7'84y]A/hE� 6̵_�Z���̣�I��m북�6�o'J��{J�����|q��>7"�PLC�G.��{p>`�� ��c�w�Ջ��A�����L��wףc<�����v>�%�m ,�g)�`�EKt0�qr�����Աkeə6��оSf`U�lOQK������=�:�cz7��1�����ʌ�q�Ԑ�`�=��oI�qf���lx�J�#;� �r��u�nT��R3@�4!|������$���[;[���oQ��f���Ce
.^*��c	����g@Mc/ X��@G��`�=C� �b��y	��5��Ԝ{���y�-4l�,�_�[d? Iz@6�V5:���GK���@�G��!-����]����f��0 n�'ep�r`|W"mr��V�7�֠�����9��7C�sR����P���p�n���>L��_hPrP<�u�$�H#���k�I)�cyx��e��Zb��ռ�ɋ��p���GB<��Ti�"�O_�/�>sJ�x2��߼}k��G�<����$G�^}��g:�H]J�$�w)�p�je�Q�7m^�y�}O(3�v�+�Q,�sQ���)'�B��oi�R[H�%ǀ��3�dhTBA�=
9��Q�6�s��!�-�������|��D���� �7+�k
�UJՁ'���>��D8��nov#P@g�%A�(c�]%���i
b�cG�4WlOrz�.�{0��7��|�$��A	�aD�sݶ����l�sX v�
�� ��0�lO��vB�W��>q�j��\�L�^p6Sw��R* �6��ש�i��K�:��c[��o/[KҖr��4Xs�h`�|$:�'x|�'���W�NE�}>$PҐ�-)�6e�a���/����mr�f�K��'�6*��[)g���TsP:��NqT��Ρ#R����^aS�AF6He���:�'�B%����x��\WBB��T��X�4H@�?���lI�	��Z;_!Ů^���6���Z \���Ả@�.��]Z�͔�t�H&;��9>���m�R�>��kW��՝�3;�4��.}ޘ� G�i,�:���j��Ռ�q��i�����m��¾G�=! �-�Y��m/N8��e[5Z��FI�����`�}y[�h����l;�M����R �j��x��έ*��M��u��z�N�ޫ��~B��ܛ��cc�7��Ɗp�">0*�ˋuq���}n��q�*MP�y��ߋ/�$�Sufb����Z�Di$ƫ {o҈~�:��F���x/�ǋ�C�k�����H*ǽ��n�hl�2��w-��ԟ%%V�q�� [0�)��a�@8ho)p�R@D~2�$ ��P2�]NB̀ef�����c��!-1q|b�_�o�Ӵt`u���}��JFg�H�H�m'۫8�RZ�����I3�H�$���c�!�o8��֘��-KlV��^ɇjoT����y5.(���(���m@���V����O;�@��*V^���QX�]���Y�q}��B��ݧ�5o�X	�?*�"�'���H��"0%��T�Ȧ��b�E�_��fwt>������o��o���UicG7�)c���D�KTn)hT5��5*5�m�^��~��+�D ��Cs���,@�懝���OZ$��,�D�wd'= g"J�mRB.ֱ���8�؄W�L�Y���g��m-2^k��i�� ��޻Z�@�µ�7K�f��$Pa��"�#�b�FT'���c��֭.�����3����i qȃ=>�&��3���p���ݘ$۷h�yN�E�.�d����q06�os�cVa]*��|�����%�Ybj����K��x�s�Uk�
���c��T{� aD�:�����w�a/=���|;D�1..l̽��ώ�p�6	�%�iI�ǘ�
���eސF)<L�^�Cè��)�o@��L��WQ�����eUˈ�$�&y�*V�$eۓ�yo�λ���Yc*Q��8��I
��Q9a����Q�7��JX<�R"3��2�i�Z ��D�	-fL�(��a����pM�W�t�:� 8a;�I��� ��@yI,�~�j
خU�@xYJ������sp�4a�xrg�d`ـ-�
�؎X4�Q��2��R�1�`2&�#���lO�^	0/SY&lX���5��E�8�7�#	�b�F �N<&�(�K冻ĴIgFl��(��NV�Z�����`/L�R˪n;A�XE�i�##r&Ҙpt�Qy~�έ��y�͝�z�]����˯��(��	9��u��@��溋��=�BR��o��(���/~QU">`x��;Q�~D��� �d.�T��h�|��6����y�R�y@I�5G�6Sd��Uo��}�w����Σ�>�P��1惹`��$���ay̢�]'P�.�q�l��yNA��u)���B�g���[
��@�IE�DŧK=H����[��c���E>�,S��h���='@�]<5���!F9"[Y�Py@�:�'$^�:?��r�j;נ^u�^��c��U��&�Gٶ�N~�!s���q����8b�aW��*�UI+�h�C��(U�K	��S�2���	�O|!��4��i�H68u�|�L�b&eo#�tT�ï�-�Z��<?Y��'K�Yb�������(lmK���P� V����+;(s�Mrzacu/���:6\�8�+;*Y����&N6�T$J��SQ�8���7N8$�>y
;�x 3$�/H�lB�<l���]�n���W2����� ���
]�"h��$�&l�^��S4�W6��q������@�2Җ�# @��J/xaF�6�`g�]4�O�.���S��ՖB;����8f�j=3Z�sP��{E���qf�n\��Hv�#qЖۀ�-��� �{�v�v$qF�xԁj#@2@�H��\�|��޴�.��;�Yb�`o�^s2���v���1��� �Z�� �9�%���C�]7=�|9�xxs	�OB�-�&d�2Ԭ�c
�+��Ѷ�p��
�Lt\:�1`7λ��%�q�  *Љº��ݎ�g,� !"�)�]�W�g=Z� u���K�+����^�W+^�	ho�Q �mO])OL.��=�M�	�b�3�b�v���&fJF�t�	�'�fa΀���v��sRk���xbN��Ģ��Tk�o�6?Ix% ~Y�Z��i���Ep=v4ٰ B��"��.肾vj�ZԒ`�P	'	�CO�s���LA1�I�<6۳��ޮ�W����c7ɸ��M-�Q;��)��!��0	Iv�{x���.����8�c�0�:�+}`� L^z��ȯ��VO�,"����$I�Q$B� S8ت�Ԅ[�=���wJz+^,�QK�P�Y"�hS�f l�ߚ��j�&���M���j �j�a�P�Z�;�}�T^�� ����g��d�~�W 6���~r�A-jOJlL0���
���,�^JC6(�� %�j�<�s������s��o;���� pܢ7���j�����=>���p<�"@i)PD�f�$������p��N��
����q*{��
M���hyc�����n%$C�8��)���"Y ���W�X  ohϸ�yƙ�4>$Aԣ-��"l�m)p�)�d 1����촒Aα[M��WV�M������!9�f��������J�m^��8��(�%Mۓ8��YE�g��W3�准#�4mp�~�ܭ2�Sc�#E���V\N��V�q_�p�T����yӾS�Y�k�d����d�k����|��7V���'�����k�7c��H4���k9R�		ɜ9;z�T$�v���S���f�J=m�6 9<<���"��FEM�bF��B��s���H�l��¶�{ړ���i��Z/����EyO���o�o)����$�,%�S.�)Nz��Z5S����L�҈SnY��4G|�����0�(+���
��w��-�4��J�?����E�#�%��tHň���7�!�pMH�J�6�sp�@���H-�m��S�q,/�vV�����ض�P���I��d?�z5�Ǟ�ű�����o���=��O�%y�=el�j�E{���Oї_~9T��c�{�a3���5?x{�t�n�k�M}�C����<V��{���V�NenP�F�pI���5!K�j�p�f��>�fq�t���Z �Mj�m����r �>�bf�5,pJzf��빨�<�S	Ɍ��cflV�(�c�n��� ��B��m��]]�>b�f�	����R�fJ���������mkD<���ڳ=�$�.��I<@8X�m���>j���LK��4�ZB�&��NI�tB��������sd��ƀ{[]�6|�%üy�<rz@T� މ�G#5��O?ݡ��k����VW��@Z���.�Ny�V[���2w���7r���}��4�.�:Ǫ�:D�N�#�S�AY�z�@8��֞�R����a��ϟ��c&��w�V�9=������\�T�$�V\���*�*.�5(�Q�h�.�Te�L�!�8���*-�������T�� f��_g�1��ZT|0��OF
K�����"	�Ξ��/�'����kZd,ݘ^���O&�M���&�s'�Ze��d��9K�d�k�K�ܓ6����z��7ɸq�aM �� ER��Қ��5Nh�&���I��� �ͣ�>ڕRMC�A텚%A���G]� p�U�N����[
��f[Q���3s��͌`����S�Y���ҟ�|朔��@�sv�sx�mWn;$/ M6E���YsEYX�T�7'�@�2��7�D�X�b`�p�t;�UJ��V�Z���k/���_��&��z�Es����ټ��������|�x�������dc�t��seU�SO=�E��= �
�{�5����[����ƫ��u�&�{Aw;�x\���k_/Fv�Zj��|��oU��MѶ����]��͌�Rۥ�d��M��I�,=���2��`�~g�i�]��r]?'����̸mb+�L%)��&���Hn��$�4�YR}�** � �B/��-ɹK��X�޵w��E���,d|̡�.�|�d�d	���o�4p����s���|���*a�ǅ*;vt561e"O�z/K�Q(W/�hg@��}K��M ��F���Jy;l�1���ՠ�#��۬v�0@.[�rA��-�����Z
�I����y��d�n�rH/	�r���t�R�?���'Er*�����qeHf��b��8d ���*��^�2�� ��`�.��o�a;�`�O8��4����y�[z��X2�H/����>`VAf�e�]���sz�^�����26զ>/��Mv�ǘA�k������U�s,� X�n�L38� ����k�椩>�FOS�d(���\�,��#�vZ�������Y�W�w�Z 쓹����̨�1�w���dSUV�5u��f�2���f���>�څ�Ʈ��ݾ�>^�K�a	Q��mN���Hu�_�4g�cH5��)iU��)`���[�9~�D��ճ\C������kPe<��:�>K&��9�R���2��Ϳ��F�ZS��Ц���yc��eu��<;�]D�()�7/�V�@Q�BS;&A/נ����\�ih���,K勒�����6|����L���S;�O,�W�b�N\g@ �s����n2�gZ�9�%��I���v#$$�ػu�7�d�ϵ�=Y�O��0? �N4����@�X=���~���z��Y�YS�Dm�,*�%]�Ԧ.��%PK���6�� 1v���K�3�[b�j��w�<w>>����kp��Y�l�c�G�7�l�Q}�Z���@e��ʒ�7b5p:��T���˖�-�Z�:��kn����@x�q�v8-��C~^̀|�]{�d��jf��� }pL�m>�$�z�n�)�8���Q���� j	 ��A�RQ��d/�	�X�`��W�!|�^�.�k �/�@0��O�>�l9�/V�m�;�a� 7o 13z3���ڬ.QM6�7$M	p�y��������a��	k������t�n���iJR7���k�b�[>'hX���"�N� �D�,���
� A�kA���B��Z
��u
�+�w�~�F� */�НU�9Bmc���A`�h��Wiӹǻ~��3��ɽm{�YR1���rmkDMg;`ؖ�*�¯.�æ�\#q���RqbD�&#iu��>%�銮�.{p���lJ�mX�z�f�����Զ]�����9�Y�ڔ��V/����Z������"	G[ ��Io[i)��(��<ҫY"̻�~%���
g��r0�C��̼J��C�d����W{bZ��@{��~�i�O@py-��Z�:�g�-��ʵ��+�<m�O�X���c�B���0cI��l�-ү�WY���K��K�9�\5����Ng-�Ne3�LϦ�%�|�<����v����6z�IP�!�D��V"��
k�m)�'�b��/��k��Km�g�=F��a��X�˞�"�Q�/ԍս��%.�ͪR��j7���:�\�9fPR*��p�?���� ��P�*9�0��lT��5��% ��R�o��^��p�l$$�o�`l�����\�@7���;�z9�4Ԕ�R��Z�y�A���Ϳ]f#A����T���R�Z�  ��;��%Ø+ �M?W2�{Ԥ��%>��p�")Ih����i��e�jE�
p��t�HGUz�/���C��Z(���.�H��Dr#�7�)��B@H��/�Mڹ��V�G���R�����i�?�oV�:����Ҍ���^�������$��c��baI�jM�l��籙>>��h�u�����"t�v��62m?�
T���ҠA�{;��:��>ڳ���89�0Ǩe����%�%w� �U�?/��*T�.�ɭ�HlJ��sa��bpN��q������ls^i�¹Cא����$� p!�Fg�����,�4�9}�̰:�������9o��!�5ަ�m��oyc������}O�@��,���v)�H����J��n�3��s�k�m�����1x��م�ަ�/����L��"m^P����-�OhEIv���,�0+��� ��I��mW�PΡOc5�3 ����i�<VKAY�gzO���k/-��T�����$�����j���%m4=j{�ol�:�jtA�`�g`�Ķ��7:��0�W�jI��4@�[$c���^��,S ���Z.���xKX9fP�����b�
%|^ey��_v^n��#�wH|�"�w� N�����:K$E.YB=B��PJ2�v��
I&K���k�������ǖma�t/�m�ku7U��R��<��y��.u�/�u�w�X�5���h\K]&J��@x�.���-�������p�*@>�p0+����aY��0lah��,i9����J�*I�u��Rl�@�!]"�U�)[`��Cչ)����gx��w��ɋ�1�Y�4_�k�1�~�XC;�p+��b��˞�S��t�WE����5T�?�u���T Ö���W�W���. �l�w�7s�WH�z�uJ��k�����`&�)-�I
.*�91c	%ݼ��H����� ���6%���L�md;����$���ը��1{����5��I��j�av|p�^N{���$pv�e�:�0n��6���Z-ɴ;Լ?�9���Y)�� ���R ��O���Yj506�z03���n�Պy�2�6�s� �8Hym4י�:��d{`��h���ޜ�V��]��1�����򀷪х2m?�+
��bW�O�z.G�,�XEi���s� t�Ã�>�t��@۹@���*J�E5�wi�a+�LԪ�*R��������!��.�������h�ѢB�'����ja�V��k����Q��^�5��{hO-%6��^����$��{�4&SѾ©(���R`�j�0$�4��%">� �9f�)�\a�*L�fe{69~C=�4i �e����q}����=W�z<�W(P\w��ԜN���JUJt�����8ɝ���4��jQ[��Ibi� $�m40�p�ˁ`/�g?��K�
�����$BT�n��{�f��ܤCW�jв���?�b�0��(7J_��sz���a�sڞ�R��� @�[��0��a2Ɠ%��l��0�m�0T G������;�QW'ؐ
yY���B�N���Iۡ��S�E��D^v�Y��� ?.癨��ܗ��g�,g��+/0]�� Q*�KJ��I�#j�qP�{�W;٩&Xn�y�YJ3m�`��ܩ&�mX*ʟy��jg������b���n�����D%;c='j�X �V"\ �v����U�Ye4�}���ݟ%.ϯlr��x "� '��8F�M�N���|�au��l S��|�,��� @���iq@@��ΰl��8; U��k֮���T�K3(oВ�yL@�j���Z�z�:�
ԦE�J���^:H}���8`蚉�d�����iS"̴��5�����l��d���Q�� ��6�T�{�5j���uG��~� �D����X�d��M1�X8w^ekv���@� &���uI�>��,g���xXڅ7���)ƞ�0(�I	�N�� �F%m����t<!��; ���/{�F?���ӷ9���K䙊�h;f�#<+@$��T��U�96Q@8�!��|�v�q�,�x����6@��|�L����8�U>�>{�E7���w�i:7t�+�Cq�Yb�P�P����"�F�&hWՙ�
�i��
	�^�R`
�0�zVE5�G\��> 8:�����n'W� �,=<v$��>-��z~��7�9�^��@5@#5 ��2u膁�;y�T�v� ����5�{.,!{286���X���L�1��}��.��9T�"������\:7�m�pn�ڶz�S@~�f�Mi��t<�՘vx�	Ɓ�ٙ����F��T�w�����.O Z'�v}C�f.D���A0K��|�=�%Q߇���2YM��P�|��J8t��n�k>�e#K']��l��+k/�@c<#�/����+�����Q�z�,�)�m2R��|<c��C�4�|V5(
H��/ez\p�~w��
���9�*�w(}�yn����|��3��\�!�ݒ,�� ���z�!r-���*Uf	���H�%BO�L�'O~���Zt6ڿڏ���uM�ks��ZԢǴFF��x��[ \H���庡@��k���x�zI����	�9H<�g �y�7j�M�廝\.�r@!���2�iu$�b� �jX�����7Kw\�k�� �~!��ʧ=X�,�� ��>q/'�9���VS%�Lw������w���r���@p����!(^��	�nk2 ̎EM�K��(~P�|Xor�.�W�f*ڎ\O0�m`�c,͌ŀ��ӖK&e��9C�Z�s�z�N�c�В�S��wg��ץ�ʒ��O3;��:w�<�ig>�,�sP?��S��t�S�p�R�Ńt�,���P�K<�CA���o�n�Dx�Y�n����{9��
��k�W�i�u�d����\K��6r<��X}ט��U����3[
\��9)FhƜm`f� ��Ya�xb5���d�_I�$ג]ad &�+3h�\��f_� �8�;��uH�����0�ܪT�n�+�s��y�&��u޸�W����Ru�;Ktl@�,��ؠ8�:���π�s2i)� �d0��zI�3]�M�v.�����K �dH�Lʙ����@K��)P�;ˠ� �N�N�jUd3m����6;�>�e˖��v@ۄ/������ �tl��*O�#�F��Mg�����m�����]%�묚e|L��'�c%���㐊��;t�����T����7�p������z��A��{����oK5^]�m�M0ϛoF&Sf��ߓ�K[��:����]���1��.'�uR�5.����-N���-�E
�\��"o3L��,�Y�3�eu*�+VGr~��蜨��N�m೽��WHCf��vl?�ޖ<{p�6�v�9�U���������-!p_�Zu�o��w�x'�o�I�}�ȑH��G������]��o߾��[n�吀p�P�,�8�H�ܢ���}�Kd�Uﭺ�}_-�4�	�󦤕U�Yb��lJ�M���dI�R���{e��kk6��,���f�v�'�Q$�+��;��(m���Ӵm�� ��4k�k�Ma�ҔJ���UD��c �*���RGq.i�]}�*P'�v�9�g�C:�%J�1�!�7��,��B;��s�b�\�b� ���w�y'�ǎ�=�����_P����X�=�#����;�%y��>���5N��&��6}�_��=��{���~繰j4A^�#����d�_��M�5���ZH�[/��@�1C8���ĵ}i)0 ��i��J� -Z%jFi�#�0��Ժ�ѥ��D����v����c�P���<�,�:��Cܲ��������w��Y"�� H �m�F�ڳ#���}��� ��$�������_x��{ｬ#�ڣ���zP;�5�5j��������������:g�ިQg)+��h�L�,�e���4�\;MмT��J��뚛 � ��/�W+.��h;r�Q�&���`"�����U$02��.  �j�"�^��m;�X�h�P�7���@C߸�RjK~w�OKD��*�"�m�n�a�Q�2>�*����3�;:�y��	�ߓ��v�~}��l��;R�IިV�/ilO���h���)zݢs6�32�{><�v>f�g�� �g��M�`f�����F?�!m�HK}n����Z �V�-��@���}Q�D��b�̒�� ���dG��h�i��o��Y�s�� -���dk��:T��-�Yj�(���6��vF��vOT����ݻC
�:� ������������7�����L���:�0P���h���)I�7���{���u��A�:ش�5T�]�_�g`�9��?{���I��$������?z^��<�:�@h����o�ә��ܖ}R��E�l� ���QgI���	��� �߿?�LH��-���Q�Z:�7�*i���B��C&NN��}�����vpqh��ӌK>5�.,1:��'�K��y��:/���Y�A�i�;$���{�����C�Ь`�i����]  �������G��Es�e����=zo��kuޠ�1@��Z8߃ߛ��(=W��_l�b���-�������7V�T�y�U�sV�ۯ{���j�pMFە�z�k4�/��[~�]~��O�A�T���^� !��3ɸ]�1X�3S�n��V�F��'��XB��E�<���,yfIС���U� ��ўU�V���w�ގ��1���Ԣo�>_���w���������X%{%���^P�O��Hz�
������&�o��L�b�);�4�	��@��&*_翣4Rq�f��n��=���A �M��mvA�Z \P��v�z��|r���J�����:Ԅލ��D�0ԗ��6�K���q8D���`���\ :�iϪP�;-U hV��V����֥�H� �Ν;;/���]�vW;�$�Z�_����K��H���hR�
��݌FBI���Ԑ�Q�(-8r���`4��������ý��9��<�{CN��w�Q%$<���1�/��K�|�=�(!�QS~�<��$�o�
j�D��V�1H�� �:�!��K�<�
���	�&i���\?)�ԛJ$im���{���%�z3���8��k��{>�S�5T0�k�9���`o��8�#L�]��n����.j3�Ԏ��i<"u7�����������m&��a�?�I9ĺ���4^�P�[��{�'gùRט>���p�B�5;j��%�J�@�]8A0I��X�Yb�;tCC�1�q�a�O���'��l���F:$*�e�:W���	��w	2���Us�:���wz0L���勏��V͌Y�����k��&\�%�n�n�3#3�ӽ\�!��2�@�2h�[�a�X����0��TƇ;��7�}R�/�^p2#�:�:�$�,��
A'S_zBt�	f�A�s˩�.B��R�m�������r�e����s׶�t��=
�=�0�9�eX��	䦦��$N~��^f��!��_����̐}㪾2��66�K~F]��%(�Iwm��xR_�P#FbDd��})"�ֲXZ��Q_�{�Xn��I�_|�r?2cg;`&����+	Y"#aݜ��7�q���ҙs��g��f� �7�vz��
�fQ��&�z�̓��sA�3�_|�
R�yt���B�(}���S�烍{`R���]B^���lo]*���CBh����Sp�fC�僓y^��ʲ�xO#2�3k���8ziC�0�k1��������H��.N� L���m����pP:y�ɴA>����×)$�w�v�:���&�AC[gI����s���q�2-Xi���P�H���<l�2���I����||z[b��8�\�2~� h��|�Ӿ{�o�p�y���9�zu9E9�������J�Ϭ`Ɍ�����#�V�l�'��Q��ާ�5`I0��)��՚s�]���(%Ps��SF�mr?[��4`��4;N�&f�b;}�[��-�]�|�i� �SQG$2"ޙ���kBNԮ�<�
#�
:o�μ��MS���\�u	|f��m��3E�"j�k�"�u�}����잡����u2�#Jz�q����C�݀�2k��U"Z��t}G�� 2,�4ri��c���@f|�E���������65�x�eu�c��Z�*;[}�~@�>b=��
����Ʌ?��t��G������o�Fˊ��j(bߨ�7ZF��M?,9:z��YkYz�~���ˮ�HA��A驹����޷U������-i��(���~5�e(�������^iе���'�ih^䥾�nro/���g��tk1��R&z�#�)<~f2NH��m�벮=��R+4;n�D��~���LO���q���:Զ��ZtSE�B��p�Z����.!�����u3T��Szv�x����8�2���Fh@�	}��\0�7��4�oWݮ���bP	Fv��W�T�NTw�ޯݯ6mlc�fF��3DS4b �&�	��{�A&8�S�M֡d	{��9֫��G������[�^����[M�����O��O�4J��u&_��6��+˩#�%����J�{�����l37�;dP����q�Nʔ?��e!���}Vp�L���0�!<EtW��Kz��5�u���U��?UL9����|��M��M4~^����m�ϙ�"aP�J�2��u"w	�|���V�A�º`��E�A�>�r�(�vRC@�2��n!������zuN�����5ac�l_~*7U?��_��8u��I,�1���t��GD�(�
R��i̎��D	j�6/�a�=s!fg�_ �<����4�2�s�^�:�M�|��˭�|J ���X�5�vd���e:S4&�����B<Qt.���A�g먻�"v�R�1m�qý�)�W��K�{�9×�>m���m_C��.Eq�s���[�&�>9��L��o�~��I�`���5�N��
ϚKl���S���©k�Ư���%�<hI9��l���}E����hL]��n)d���)�zǺ���8�Le(�܅��r<]��ɺ��P�N��VA��4��=Z�v^��˓9d����i��r�  �T�ښ��7��JE�ɼNc�F�&��j&��c���Lvg��	�k��C�,Gq�0�\�����v�y�m�%�7��s;��6�An=�⊚�0�w<�Y�tH&T���`ć4�$�ԙ}�@E��M���%=ƨƖ�V/��M�S���G).iye�ĭyNM��6,?q��6���+da���yĉ�(O,"�MW�	�(6���J����]�cK��Z�_O��Z�2�t�*2�V?,�A!~�*�H�� '�]=��Eb�eǊ@	�S��g�ͬ��
���&��~4OE	����A���Y�$�Kߊh��܂eI�h}p��e>����)*�ֲ��-�1�u�!����z:���(Yr����X�t(lh��)��<kn8M��#��P��b�ݠ�UO�4<�vdX����V�~�����6�Ŗ*sI5j��p���?S��?~���+Śѻmh��kI�]!:���6Dp��M���U ��<����#��f���e<.o�恮�6��m�O 6|O%��Yklp�����+m��' �!�x�z5�0�G����ۘ�I��YM�Ğ)��UG1�'D���K�b#�1������;U�k��ޏ-mW�5}� YPH�Ō�oW�VgT�1�Ũ��3���&{8�x���ڼ���^�,?\I33�kC՘#���M����Q[�2~I� 3����2F�����~�
�k�S���xoɽ�צ��N�J=r%c�1g^-ts�n���(<��}3B�>+\g����]��?��^�~��NS 2׭��8�P�Y������|r�*���9��^�N�ab����t'�m�G~4e�;�{)�ς���Z;�Հ��fR���s�k���!`=�^G0U�HP�l�7_��Q�!@�omA������%N9�VǨ���'����=N�A��%��=�����t!�k��E�en��ƝE����I<2z�I��>�x@T�Ӥ(�j!�\'���\�^� �2�vH{|&�#���V��ӌ� ���7-0rs�H/P�_r?�*9[gt�cyZ�W�Y5(� �$�}���]��RK�+IՈm�?�tA�A�;��Y�'�ͼ��d����F�8h���h��hIR��%�Cu�'f�����l�B��C�r(@�z���=�פtb���~����XU���E�z�;�p�yK�ޝ\�D�1���J�zx��rX�M;�>�woE#yuĢ���add �r�˃��Y�vޡ��ឞp�Fh:����ru�t�CjA#���;��.��oE���������L�$�l��j�~�m��)�"������#A
�_"!n�JQ���
�:��[�%}�(	/����b���|����O�~�g���F�`�Q/_�������a�-O�|���h�ԝ�<���:T�<Q�bW����d�mؘA�llk7�)@kN=�
X�M4X���E5�v�R�C��Mބ�jJ1WDRY�Ҳ?-lc��\�^�C�	��L2N|�O�eEuf��Ւ6+|���t˿�<*�mjH�za�x���og�@ę��L�ԯ��vpx�5�#��(��=go_6��"�XPtE�Jۀ%<�4�Z
�%���\�֮k����CQ��m70�0l�:аf-o*����`b-� �{lE�)��%�wmG�W�J9�-fBF��j�Й] m�!����N�	{AQ)F�O'�rq��t����P�ȝ|��8]@R2��N|�\##�X����J&���6|��o�'";7�Ŭ���I��c�I�O����Lm���k����R5*4���t��!a_�VS������5����i��ږ�����t ����A	z�*f�i��Ҍ�n�Z�s��v���'H�����������4�F4�)� ��~D�e���e�֠��B�΅6�]�>65SF�nd?9ξ���?�_h'%������dػ��ށ�aI(�s�c2�D�>��m�*l�FVIW��ƥI8N�(�<���Օ�+�P��j��N|�h��}ͯ�/���U����@l��T/���ٿ��^�ST�A��S#��L���nI���m[��	�b�)�����n.��懌��au��Hz�P���{��j��4q7s�c�w놯e���� �����;����^"P/C*t.�}�Ӟ�6�2�9	M"�{��<�zu�&o��I������e2���������o�Kd��U�U0�[�yDX�xQy�q9c�"l�&W�ix�އ������絼}n�
<t�K��Zڭ˜�%�a�������%Sg��?έ%�`0��2�aF��C�m��b�%�b���Cg��H���<�K_�S��:�&1ڇ�s�-`*>�	B`��Eͅ7��f���خKs�����;h/8f���(����c<�&�M�)Y& n����J����PK   �cW�����  -�  /   images/6bda90e9-5ec7-4d98-9c70-49b6fbff5641.png�YS�&L�۶m۶m۶�c=cώm{Ƕm�<��3�EWG�UgFUdfT���$<��������
⿪�ߕSm-*�$-*J���hamg䕓�����t�{](�#�\6B%�K�$\`"j��E�MՎ!�M�*�@������d b�7���s���1��s�u��u��v�Օ �F�D:���k�>���Z��R�0FB>�qdx8�X���?g�ȳ}ս���w_t�P�4$�(�r��������Rr���8W�\:	4���x
�Lj,�@�>^�9��8_6j����^#�`�I�Tl=��ll��$���7� �}�x`Lf���CrZ/FԐWts�o���÷��$�l�`�Gh�F\E�I��ғp�\�
gh1`�?�9$��Y&���|�F�[O�Ī9d�4GN�eZט��SN�:�*��������0�щU��Q�Y�;�θUsr1����)��4:���8�>u�D�X��"k2sR��(5x���0��XxT�pϭ:nP��3��+W�K#���.���\mAo��(�«��0R�EC����I��9�A��:��PkӠ��1�K�Cg�1��P,�� ���v#8b��C1�*l�0��f�-I�7�;M+8�f��ͨ��X���1A��@􍠦���!g��@��D�������=qk�GQ�A���(�����1q�dP;聬��;a��!��Ċ ��R!�/�=���4Fj%RA��+���EM� �#W�J��ՠ��/
R��`���#}
�����%�2.�)��B֝���R���V��;��A9���[����N( �3)xR֠������$�]��j#�RģԦ첄t��SZ�iE��˃�~�i�v�r.������?�'�Ш�9�5Fz�n�x��%5#&�+#`ʗc�?�D�>x�ˎ��߃��a3��_���|�(f�ᾋ�x�u�h{S�n{��$t]d����Ὁp/^ R D �`!�������̚К����D��j$sr���|5#
!�n�h2�5����zb|"C��t�X�,K$_>i�-e>�.e_���ydc��d����{��j��4@�Z���z[ŧDN�CÂ�QmF�AS��O���LA���;yK�O�OO��j�*����v���q�zNeTe~�P��{��� N�����[3{�sLs O�����y�ӿ'����ʬ�:�(-4-�6.�ƃ{,ظX��۱�<v�>>��ψ8�l��a8�8q8���,��l�l���+"��V��:�-��E+spp��_���3^�V����;U���b���B�EM��!3������17����YyeyR�1;�=�r�ٙ3�F����-Ϡ���O�ϒ�r�Ep0p8��(����p�p�qO������>FrL�eX��7L?F&6(��+��Gԫl��;OI��S�t��#W��+9�y��_��v�fI&����PZ�ZѴo����2�yT��,N�i�7iV+w*W���M��'F�(v,R�#�9u)7�6�[�ծC�`�t�w�t����n����5����=���xn\�����=t.�N��ׇ�/����L��������֘�{��׺��O�ӏ^�o�h�X�@n�ϲ��8j�GCΚ&Dn��g�ul�ޔ�?V��\؟���>e7��G�����P�	8mq�r��)�����T(�(~��|_~G�怤����A@:�t�.�?t�o���_��ٛ�+#� ^H\Y��*X϶�2��+�Fs�@`����tg�pX۪��L���#�ǋ�"<G� ~0h�*�u�}���"�v3���寢�l�u���Ӽ���������uO�g=���|��C�ak�t2z�H�Ż�GQ����!Q{�D�ٻ��⇌"��~U���H��|�&�@�	�ͥgS��9)K�J epQ\E2�K�KK�օ֟�#���w��ؔÕlξ�'�SQ%�R$�.�Y�t�i+�밍�.gR�n���+ٗ������O��ji��m��΅�wf'�&�&7�.{�=�}��R�&�R��4�k/f���y��[���oW���门��>��"?HJH��{Znl��~�>��
�|��P�ǗU6/�.k�^U�M/SV<�v�mI=�z��R��CN�M<L|p��l5�w��Mv�ĴP{���HlQlR�AUX�;4��0�R�zV�U�xZ�R�������t�T�W�V	�b\߬�֗U���1z8��X~��M}t�jT�6�\��߁^�3��C� :�G^�?�F�vz��:Ɇ��˓�0=Gv�8f��s#����u��o��ǧ����*(-��7M=��֞V�"L������e�}���QV�P����Uz7����DzJv1C�k���r'r�{���a��7����1�>I�������@si��~j+��[��6}ކ�;�+ϩ�м�ֳ��^u9E_�{������{����������f������/?��9t�/�#�1A*_� C`�w���.����bOo�j���������l�r^*��[`��\��I�7㇡�A<�w��i��E]�����������ª��Jϲ_�o�aWkR}�-�NB �{��}?�JY�,s>�f��ś�O˳�]��)��)J�s� ����B�d�	L4�}UF	���At���x��d	��J�B��T��!����F��ۏ�ͼ���t~"����R���E�%J��v��Sq��? ��d� z٫��
4�'-&��ep��w�ї٢�99�ե;�A��C��f�\R ש�S�B�u���	k����m}��p��A2b�U��<�ɽ�{����͑ů@���W�M�	^�)� j��Կ���ӵ��K��`E���������{VK�.�CT����xq~>�@����(ʄe���D�$M�|�<�K����C�G���q����AXW�?�fQRR��˛!�7�ɲr��8��X��G���xn��|����zoQ�Z�����T�y2aٝ��G��TE�m<6h���d)�<� W��{��`X���Jq%���7,����5�KHH�,��)Ij����N5��mR-�<SiM���f52�:9�>-��3?�C���]S�X99��~oК��Y��{��g�H�|:�f�t��b�� r������r^�@������̠��p���O_������IuxyQ�F!X�q~���e��]I�|�m��nQa!xYCݭ3�UE�3K,���<Y��}}�
�J⟛A�a��0\�Q��a:�P7���;���[vz�݀�����+�O2�j�[Z�n5������{�(���
���Wqp�IɉZo�>��*�z��������+P�Uΐ����陈9l�7�@����#��;�ԥ@��0���n<��e�����pszH�ZJ{8(��k.�<D�N�s.��M�8����������NƘrR�R��k�R�i��{�ˡ�n�"��^Zb.����@���<�V����wo!%ٿ����V^���;i⍀�~Xe�|����u�1���Ns��#���Gn��G�<��x�2u�<�0*�;M��ѽ�Jw�T�AJY& 0�SN�Gqa���6��:� z���0��股5�,Y��Ṛbih+o��cS4qrRRZ�x{��j�x�oq4z<*���%��sԋT_<�I�kj�QUOx�Pw���ID�M5�4a�0A�!����y'*?� �ˉˠ6�Iw��Q��;D)Ɖ�ԕ��wGvqd�s�͸l�Wc͆���n���4�3Y�e|�p�M��T���G7]���[�-�VWW�����3�����_����'�ݢj$�q����(7�P�iW�?�` B��A:x�G����B�9��	r��LqR�I������ �����Ȟ˃��&�J����},�����z�'�v�qpp@|������{�@�gl\(+��}����Ou�w!�
 l���f�7�����5�-J��Y�9^����|�����6��$iM�i����yu8i�,,�YI�����Q�����y��p��K������&i����h�>�Hp^�X��!p�	�FP�1)yZ0j��
	D���y��pY�����`)�ϰ��r��ŵ5��3%\\^__\[�Z���������VҠb�l�6����ژ���A]575}t�^/K�!�����b��>����-�����V(�D޿��RT��1r��٨���}�H���n���A�L�"j��>>�^^\�E�ճ9�\�;��{����3pr��?��;�� �����4�45ء�������«K8��h)�7��]��L���צH3���
ZxcvZ��  �
6��&���_��'��1ˇ,8Cq�-�����/�H/�{&�寑����}��ux`F:z��WD|�%� e�T�h���W�uj��ɭɐ��7��pX�7��fiT���W����ϕ�G���U�>���d��� ���t�Ɵ%.?'/M��4�k�F;��Ŕ�MO���:�v�x�X3Z.W61����\��B��I_J�_A������sUT[����!���+/mf��kJm�w�0Q�.�T���b��s�մ\yoa���@$��b��#c��j��+']F7uZ�ta/L5Ҙ}U�V7��c��ۘ��2�`��#�i��J��M�Ɛ2++3G�q5��n��캸�ad8�G84k��)o�QA�"-��l���&����8�ү���'`uxZR���`&�ҙiʱdy��Nu"I&O=��<�̇8��gtj�i��]��}�% �T�+�p�vg�נ���@�9����o.�Q�����7I�sq�vA��@��ҟ�R��it�`�%Ԅ��AU"�LҒ�]��.}��4䉓�2����n�1��nV���h�/��M�����1�� �m3� z;�f������ʬd��a���:��<�N4)-)*�;L�v�XQ�Nt���_[Q1���U�CcI��ȴ��١�,�}����3ptFL	9�hv�ܜ;sqyt�#�W�F�J���G�Hq�����Ƨ�ch5a�����X�T)���^�c����f���d0 ��a���CRA��i�
Y�N~WȝB!�n�l1�c��ܡ	�X`����9�������#���u����`GJ>$�2@���30T�֮x�w{�ld�����{��k�M������\��@�]�x�3���g܏|&����Ii����[̦Z�wq�{���uu�������)����/=���H�h���>���[M�A8U8e�9/�'s�i?("��)ֶ�N�4���^>���6�Ϫ���Ϊ���ɪ;[�%��h}��Nz+��P��$s�/�r��eѐ�Y-bL�3���0�6'c186�~�*�zV"8�d��_�/�P���k��J�n3���k�����M��.΀�M��5��zA�={���A���$�I�6U �F��}��|p�gQ~=�L���=���ѳv&�P9: ����=-��@(��Y#)a�}�w���A��O�9T��_����F��:Io�X!��;{�lYʷ����rVs��,;�jk�DK������	��u��i�Y�\=�U93�@+GG�>����9� �������kw���xF3�������p$�H��]�>*m�d������nu�e���J���$�s��[���1X���ԛ���*���=����.Ȟ���NQ4!L4l�+?��R�g�Ŵ���{�}kEUm9Y@���Ɍ{��zj��E��G��v��J+�7�����B��Øm��s+M�YQ�sr����qH�.^ܗ�����k싍Т����״q�w�+q�l��r��Y�[UQ�	F�)i�dp��%x���v|!���Ra�X���f�v���F�L�v�û�%M�{E31��<Jx8�u'=*��+����21�2����a�I �&� �fkg�a��?�߁&�[������>�9�8O��Ǯ��$�j��CZIk儧�a���P�[:z��ư8�WE;�<��IpF3I��R���\펺,���I�s���󶯯
�m�������C	��C�)�/�HB���8�����	N�&*sp��Q:$�����[s(
us�Mb�(�Ww�����2S%�~�)Ǭ��T)�2ZP� �.�#�<���/>�:F����(z�\uZ�ܴ$�=���?m��|ZT���.�Nq^�`�O���,Ɖ�U����U)8
���q�/TBp������Kr�`$�^]��F���hʯ�|'��r�����`h����܎����6^�S��Ǯ��n��'��Y�c�ۮ>g�
}�v�1�>� ]gt��s2q8��5J��{m��?w�m ^�)n@��r3n�é�3c#�>�q���(c�꩚�T���}��o'����gikml�O� �Y�*��j�~��t�[WI \%�x؇sȏ��Ϗ[s�%�b�ݢw���"[d�ƞ���m�k�{�v��)�ٽ�����׾m]klz�7��I��:Wy�_�t܉��@6��I��e�?�W����{���ՙ�"8�5���.�������L=����x&|���Ӛ<.��ۿ(�<2�q�{�Q���Yx��j,� fW?h�t�,Kx�i�x�m�|�m�,�|2������Y���T�/�.�^�{�ul��ܚ�����>j����y?}Չt���ش��(?JQ�ǯ��E�����n�Ѩ�����ւ���{<��ԵkG8~��v��ͽv(
G�/�<:��)[��8^Q�V��N�tqy0��i�P�ՄeL�'���N���h��x�nnV&�j�@�i�|��b�m�2�7S.f¶6H/�j���������L��y;D�qQM��ܡ�R6���ԗ�o�}����u<n�����u�1W�6�+����@�B��ۏ繠��y�B��w.2?��8t%d�d��Cⴘ��pߦZ��K��r,�r�l\,;X�9�3������0���	Ws��?ؼ����.�$9&�^f߃��ae��#�����;� Gs���NBH�ꉯ�
��n��j&�T� :U�l\n��eۣJ�����Ou=0���<�t���R$߫�HP>���$���c�����������0�T��e�i��.�$�
������8�p�s� ,*9�2`s=!�H��S����1�է�vH�է����&��2�kܳ�h�t,�-4��G�X�CiO;n����j�wVLx��0����5��r���X
��(7�tYD┪*9���vں��e�Zw�<�4߻���ߞM|�+�R�F+P5�����ۮ2-���p��5��{��/�O��Ȥ
[	c}WUZ��-=>:e�U���j�]8�fy.����3�����MȜʸg��}�b�`u���tH:�;��j6zӝY8c>�7�^?��|������ ��ق���f풙�����y���\��j���v�mǬ����o���"���ͺeK��zIz�ykU��yN
�u�1`��<g���]�i��e�[�LUB�)21a�z�0%/�t�H%�� d�!�ߔ���/�5��!F�#���'jPQ<*ê��0 �� #(M�N�T�_��T�6֓xY�}�}�����a&���N��L��d��d��o���"u������,�ՠ�E��jܞ-Z*�������m���=y�@�q��HQ��w���MW��M�H��0�B�\7O�H��ٴ���*�v��L�$ٟ�u�� Fx�v��%�֦��n�U��:�+�s�77Vr��
�%~%���z� �'��y����+��R�+F�/';����xum�6��I��������fy]g�>�S(f""+�k���E�}���x�2k��c�/�v�ky�P�(8o$�r�K���q������J�x�:����/�9mO�^'&���2N+�;�I%��J�("g�@�G��6��@HV�����l-U��u���f�Xe�!��S2����E�O#�r]��5��3�1:���,-��;fD�[�!��
R����D��<��>iovG�����U�Gm�|}g��kI���*�Y�W!#�p/��8��r����a��蔵P��D�>��L�'�ubu7���y�ڧv�:VB>$	��r]g�o�4��M-��1������o�3-���C�s<>�>xdY �+���=5��^������K��{y�b�� ��u#ʷ�
��f����Kr����e��F�˜4�a&�
&���괗�i܍x
!�E��q�I{\m���󽒉����u�@��F����Ex�֗O]�.Zz���.�S�ćV=I�!�(vL`�pEa�Ed9�v{(V%4��(M��-<�ң-�U:�	I��0<�-m��؃n y�WϷݟy���xJ3qT�Ҕ�gq�����XOG;�{���i����J�~�̇L\Vժ��s�R�2��Z��˙��6��?�l'�rw�1�B5-8{5�"J.�����G�0��ӣ����`U�{�����݊�溉͍�ע]<w�͏����Q+����[�5.ɓlI��8�y��;��A���`3�5Vƭ��/��/���X��ì1�-�����$$Q�&�d)hi���n�E(ޓR?�X��x���q22U��p��>o�'O��*��� O��s[�ZM��OZ0�ǏTLQ�!�<S{�a�".��2�I7���$O��_,���ݗn�Lm��4x��A1��O|��i%*S�63���؃jezs��P�(-aK�2	U��8�rQ�0,��˿o��|m�𯼈%|��=�e`Ԃm�b�	T�ޚ�[-�]�JK���.��f}�.�E�GLu�R
�A���a�(��,Q��/���(����"SB�`���Ip�K�89�X�'w���V�����l��VAl��e�
O0 �aZHTR��[U����'
�`��`�{�8�]��˙�F�+o~��x�?+���S�oʎNY�T�t�m��#��ot�`�I����V�e>��(���c�qx\Y�G	>?C������@�r�>\+sZY>&)}nG��|N�#+�����o�Zs����~�zR�2�K
�J��"��xI�\ �ϣ���5�����l�$w�m�4a����ߥ�!Ⰽ�[5v�k�'�Jt%8O�@�5�$/_~=���i�tO��]�9�Hj{�̖��_��v�;2��w�c_�f���r��f7�B�R�N�7����I�5�`��c�QM���S�� �l,�#8c��	��"]H@���OO�^����2���\�"�@,
k:�2����@qFu�_�k1[%���Eꏅn�ON�l�0a� �/|7Y[�~ K��� g��Mgk:F�g�q@i�Q��b��$y�xk���~�-�l�g�<����Y'���R���{ڹ�+�.��c��&�a3�詩9,���usw'D��y"���im|�y�0��<sGZB��4��r�hla�׀�$��<7�s�P)ߴo�F��_�츼�ɽ@�xZ�Qҽ�����t��G ���Ev���t +F���X2��W��M�gbVGN�����%������"\il*c;j��	�Q��c=�jԢwSIKM����Q�ӳG�1�l��k�	D��a�D�(�������)T�P�A���b\SW���zm/����#�jUa�����s�gX��Wǣ�LQyx�fK�U�JP��� ���)��kc��N^=�/������\���S�b9��|�I�����+z������F�Z������������,�<��p�������a�����όu����>3���H�qi�������ؙ�� �'- ��ƶS���;
{Ǔ	[k"Q�ux�)\�>m���ۣ�ƿd=��ͪ�l��P�7���g�B�=�֞7<�6{�`c7�]il���RO����h}h���9k���	 ��qD/sC�U̂ןE�q��T֐`�{5ň� Ke��j�fi�P �)�w0p\R��yI)�}��i(��Y>���8E���a^��,�`�R�A�P&�bq���i�_b=J>=BV�uA�����l[l;��\}�h�&G�7�2�9]�U�*}nߢ�Y�@bd~�D{����'ە��rө�'9Z��`���]V���5�6MӼT���-W��M�տO	2������p
|@f����~8f���>bOm�[���#��|��M�'9J"�PB%�pPd8Ub:�CȝV~?E�"&���ְ�٠Э�1�� Lr`ߋ�sߙ��T����s�l	P7��)�ǀ�cD�x��	���'�fd&7u�.��2����q��յ�6}f�QP��tq_P]�`�L���+�#�L<20����7+�ݿ}aG<jW��J	k!^�Q��ؘ�Xs��ge������ݡ������w��إ�G�����"3iSo�k	�C�n���S��Z\�0�u4th2�xV]{���P�b�5T��A0[����]����eHJ�_=�0Bs��=F�x�]v���[j�c�ha5���3��X��|e��^$�^hn~j�z�*G�Ň+C�@GA�~��h�$�~��3�SBs�kg1a�Ј��uT,��9��mX�n��ƅ��\�������*#��c�d���ۻ�J�	稚�%����=����6(��y2ةc5y*���j�X����,�	��-��t�j��+9<����m2�螵l���3�C��S{#��~���|V	}�m���V����Wx��l'�P��Hz�$�8hK�h���Mޯ^x�M�x_���rRV�k��gr�o6l���RA��B���9w�r�/�znx�����Dn�����7�휼F��6^��5�	Y�.E�׉��6����l�i�!�3iKtUjFܝH�Po�1��[�#�V.�t�a��w��hT���Wa�1/�>�r�/Td�գ��Q��q��	wձ��X�yV��>��%��HQO����ȸ<;���� �dHrK�Ѣ5M�F_�7���nwܾUT��՚.��/���M4�T�:���c�����%D�0C���?�B��UX�j
#����x9��ː9AY'#��/@ٓz�7�wi`08�33�E�p��-ZN���3����k�5��O6��?f����h�Q9@_��+�������'�]KG�+�I9U��Ԩ}MFN����Z�W�i
ƴ��E6h�נ3��_Q�< K�JL+Q����0�6�����#i�C_U(�^I���}�	�Ҩy�7����)H���$1hXs�h���b��qz{V\:�P��
���(�Q��ޠ�5�qjb~�R{Y�^����l�{�88�|I�{�%�'��!�3TIR��`�O�"$�K�ă}����m����{���8���j��hS��L�s��;#����A��;�Yz�콇w���y���V^&�0���є�=��{����%G�p-e(M�;ܾ~�Y�=�ωUð,J�+��R�����Io4=�'i�8�(Y���p@G��J��7�;����0'{���5�Wv)X�6��2s��ȇ1��@*��稵qt~��
���_��&\j6w;B��c>���8��3����AS�o*.����P@��lHC;�#iƤNp��YR�H�=��i����q�d��yp�h�QM����j�d^!*�ϑ�}�K(��S͛?w�|��a�~�'�G(��U&4�d��'y��rĥ��S�h�雝1j���a*�3����xxH�B�����5<d�����Q�[P3J��b�t~��'��\�5��ʘ�d�	FJpp,J&����.�Eg-U��"#���+�̃����S�{?\����/uu�'����|�$*;h	��V5�k��v[��4�w���&d��A��A�u?���޻���H�
;�e�6��y]����ؒ�g^���r%�}+�fv��߮|{���ƾ�q���	��@w��G�q������wΘ��`�Y6ƆdH��4�[ ��#�F�H0����»wG�4�B��&,F�rST�s.�i���.fy��z��J����8Zc����� K�2H񫡬���C��	��>�u��+��o��o6X��W�*+�B���in��������,�������ll�L�	�N?5;k{y�ø��ʅ�-�#�/+�Z޴���3��)=����n(�&d㱠@k�©ȵ���e�i��^o��hօ�؞)����Y��67��S����1`�HuW�?�r�u�}���`z�7�X�Uf .#q\/+,���p��+�z׎ !�_B��P:Fm47[����(��W���֏Z�����j5�/
�.��YL @F�PfB�%����ى
���T0��`5y�D]e	����cO���_��J��٫�x,`��	E���^�<��:��ѕ�Q����\����B�,���ŀ�m'K>�g<�~�o�wnn�~���X�x��0*��c�*�2�VD,IT��+˱nt2K侜��ٮ�-U˔��ƯF�0�&�"���X������qa`\�Ee z���)�AH��Y�MB�*r�.��=�f^#�>��i>��P~��ĕϹ7��_)�Y�?o��k
u��H�LNF�,V��%5U��n�6�!�T�Y����"O���6���`�\�2n�}$�2N�����c�ll~��sA������Iv�Jl�����l��:t���Ľ�X��BcR��c�d�2�ѝmX�C����_��`L�[0zM'0	w�@�����~�n���2YM�H�S�.������nt���9�G��	;���'8�h,8���ʊ�����J���`�K�E6f�|� Y�tz5nu�w�|7Ȁ������)LCe�[w\RO5���i��b�tAO�Zs*�1��\��~GI\�>φ2O�,t�2��+��k�LS㫄�,�w�z1±we=�/Kr� p�\)������AL'i���ە��2wAOͿeսˢo�`Y�����㝀Gj@8P'�~٫,����6DJ�����F7�å�NJ�g�XA\L�4����&�iv��rb����Ѓ"�����^��&ϊ[����jeb"%�ĔI�R�����oC$�d�1z�}SIOK�n�fXv�$$G�~~�>Rb�&'c��b�>��s"����-����$���i�e>H�~�в���z��H%��<�nv ���HN6�|��6��ߦ���H�\׵24�����JB�I�+��j-/���d��K��9�+	�J����Q��ضX�7���I\�.��<9�ܶԩ�%tm�����I����4�tur���8HҲ����T�uG8���[�ʾ(�Ȏk"��/a�oY�H���_D��ė��yɆ�^�co'mG&´fI�1O�B��m�HX[s^�I	g�GA�҄�WpD�k��mt��pc>������ǋ�S{&Ez��/f˛*;�vR�Li'8���Y���ŧ���u=��j+_�|8��I����6l���/J}G�B�|_.)�4���V���k��8��;�m��$�l��|(��yn'�� �4M���A�f��ה=^��L3�����93�;lo낿�?^;L�Q	�4ZL�K>IBO'KUp�5��]��}�=�]�)vI�����8�%V�KE)�HN��5�0r}^������;������������$F$4�$"@��hy?�����a�=��{Gń�a¡��%�ԓ���p?���C�M��$DB4H��~Ga"���:��a�{�v�V��(��օ.܈b�J��y���A�[�p�N�3�G�]�j#�ל�k_վ*"���42 �ͅ��v�Ȭ��!��&kbË]�Пk������2v�nIr� �N���%�����0���t�$�ϫR!\[����a[����)�A~꘱��[X#ǖ��Θ�)��Ŏe~�l���?WM��7ܢf�n�dx��� g��
���;#�g����zo]fu�Q��^�����%L�܅�)<?�Nǹ�ت�䆺��9�����-���fh]�Nu꜄�����*p�gi)���
��z��H���������pˡEta���c՟o&�&v�l��'ՊƎv�������g<u���vy愙`"nw��}��T&��ڢ�L�a5���N�3�F�{�j�́J��o;|�\�̿6����?�|��_E��6a�e$id0��˦�A��+�c'��O7�p��*'0z�e8��v��V�ڇN��1d9yn:t�EX*�[(?_�oT�oB})����TU�bZ�[���:"ꎘ�/ �h����\!��D��(�7ь��V0ѩ!�e�s�d�5����V��GCB��a^��\K�y�I��"��,@�(xP�
���;	k@��O@;�4�3���0�#t���@�*���Y#R��`'���'G+�D��N����J9S�/uRab���:��1��.,a�q'H�l_�pv���0���4���n�RQj�*ߣ.n6����6�a�Ɏ��] o&����l5�h�������PN�\g����Q}�/'��l�%�����Z����M�<�ʖ�MxԈ�~����b���(�r>D�V�ĸA�G]�-Xƞ3�����*�D�� b�yG��|@��@�yVA&_��[�tr/�(�hvd']�<�:)���4mt������c�=K"�����ʮЖS-:�f1�t�JCr�6}_�uێo-�Վ�
s�����}�����?��'��	xǽ���CƑ]QZ�"���/��I,'�,�k+�c�n ��F3e����A�х�+����gX���-���`WP���5i�A����C����頢Yu�ݼ ~�i%:� �O�>̧U,��F��F���9��2&ඍ��	�q�8�]��{�I�[��Ԥ�"*[q'B�\�Q#�I�08u� ��v�{�����;A����L���{3+_K� ���O7���N"��l]�y����7����14m�+�6�WܖL0/�S�UY�Ae��X3]t��D���C��8�]�<��e"�ƽ��ӷ�p3����n��s��I��
�ku�]�(�/b��(���������K�}"b����T��y���u�o�6�����Ҋ�-��*�Y:툨���=W���;Qz��2r���px�{h�sv�o�o�e(�$�v�-�xN�D9@��ָ��Q=�g�F�EJ�g:	������h�X��
\U]Ƙ���^IT2v؇ۓ�a	�X�����H�-W����V_���U �9�� �[���i�� ��RYU��u�)o������E��l�5���e>:%41�sO1�i9�b0���4 �,�����f��_�t�� ]�Z��{ ��77����Q�%�L"�ʖɅ���ӫ������%�ɤ֪::�w#��Y�'�3�7�x��8Rvn;��)Φ�˝{��U���Z�xu�5�_�J�1��)9�	�b�ޟ�Ȳ�k���m���Q��"�B�P�h>�9��L�J_ #� Eav*��Qh���7895U�����7&F�c*�2�&M�}\Q��(��n#U��\z 5w�
�0m����&�C��5���*B݌BQ��_��ĥ�62|��g�K���Q��Yƀ{���:ݹ���Bv�ؒ݊�C���ZYG�v��o�&����5�fj:2F�w{�*k>�Os2���Z_��w�UO��a�E�����p��5�61��|ܙY��a����a����k�v�b�����?���B/!��3\�xaW�?����?�@0֏��4���p&H��p��/65���@�$���V���a�b �0ӻN�w��D#��D�%NVd�0�m��m�#i�}�[�{�})�� <i [���i�c�5 ��~y�u7���}���0w���_���3�C��m����!\_M2D�'*�X�<?�N��b,�,t�$"0F!��z&-H'��ֵ��PO���9h?<^@��<P���Ս����l�=7Ñ�z`���g�|�B_�$�F�w�8���5ͽn���C��DӃw��9�����Yq .$��M�(��Gl�p���D��%m`�)+~dW�y�߶���yN�(�����u.��MR� U�b�¶lLf5y���蘍�z��K�#$����h=$�(����oþm��T�7��������ȧ�kyv�=�k#�E1�JI�)+8Tn]mm �� @�15��ӿ��0�
�Z)�(B�gՏ|�p��U�v=(��_t����Q�V췵yŠJ��t�\2O;=���g�]���-#��jvV��4����hM)�R+KD�[�:����g�Fi��v�l�W�D�u�޼'�'�2*����Xץ�/�@x*X������:�Lɸ!F� �O���J��~�FeijM��y�p���%^#�2w��ڊԭ��j(�4{h?�R�E�kj .�{���3O��^~�u�\�q]R��=����]����.s��Ls�������;��� �ˮ����@Ye!���k��&	���(�`�b6��Ⱥ�*��N�K��T�W�"E��Ql�����6\�"\�u�a8i�GJ���XcZ�P�I�]h�j\d|FVv��d�d���5Q��+{��c=��q��	���G�A�	I��6�~���ʿ�-�\�d��dF7���t�-��Ïq=����/�r6�r�� ��ɢ���ʢ�(�L-~���݈1#��˹�In������۱K��|�l��]�g�p��q4����Y�@K�:�n��vpg�{��s�}�:�;���������N����'gY@`J)�j5���59���t����ހ�w���^��$�E(lOf{lV��c�XG�Yq1c8psV�@YS9�^�^һg�\s�2$����x�Mv�5?��.YO"�@|n�Ob�4�ȉJx��Z�o��iW��A?e�ZV��!Ƈ�$�˧�a�����di����o�ƲdU�S�a��{�p��T?�!����c􌨰���=�0�B��r��1�c_r���;n�:­����U���2B��]�\�lk+>1Nz��F�̡+2�k�f�{#��ݴ��N���eܸ���`D��d��wy����a� �u5*��e|������K	���!�N���\���K��������u��[�K4�����de�_�N�xj��W��?P�+�k4�ؙM�B�4�����\\��6$���&�o�2�U2�R���
��UW^E�����]R\e�t�׾�)��@��_�ڝv��$��t�zD������@�0ڥKK
�E��uv7�B��m�ö@�ܜ�3��y�]#���O��"�5�l�����$�AX�Ȩ��������:s2\-
�m��ɍ�����qƹ�SN!�����'���/}�gc}��CO��QM544�,a�P�'�Pl���l#B6ȑ�_��'�WX,_'��&J�L'��^�W�%�'b9�G3A��f�ģ�Hⰼd�n*�`�@:T����5{�"ɇ&�������fP�1t� ���~����UK}����/����_:݊�~��zđ��H U.����*��\V�g$y�u�Q��ܯs=8;�g(a����\7rh��wC;ŵ6�G�[�-�]a	���0�H�j&J[��T�O?A�����o�(��>�jI�������g���:�u���s"-�I����֬���M����b�;�-��K���ݳ��/� �*1�sg�Nd|Q�|@�d��tU�X��_I���Kz�'>������a�l���4�̍���f�h��{/�s��鱢x¬G����m��99�q��uNkU�f'35�ư�lVʍ7�@��G"4݀'�C4*D#f����bw�f`	���E��ķ^v��u�����;�z:���FBW'}4� ��J�Cpa/'П�e�+�����4d��͟�������C��xc�;����)k`3[|V��5YЯ#��i�����6���)&�%�͚�r���5b�T]&���5w���ʧy�����V(��)��\���Pvڼ5S����@D1�X�d¾E�K-&R7�Q�AOl/K�cb���oz��cAQFp��Wl��V���f*�������EM�Zi���hii���h�|����H=6b綾�v��{�{ݞ�m�ڣu�B�p)']c������������xx0�_e�Pb�S�y|^�[L���PH���t���d�^���q���N5B)~i))`���������We�8��M��,����[mk�r��{�j�]�Mc�f�t��0}.u,�]���h^n�աP�G4���(a%���0�����ڍ��_Ǣ=��r0�y��M��sr)����~ j3Z����K�z��?���YJ��I�%[^:M\��ǡ�@�P)�~�5х	Dw�$BI��)�><N���i����W��}�+E��N��]�����a:Y?ML3�y%\[�Mk���VF�e�;�8d�:V�0d`�� j$��y���ZPrȑ�p�v$���~S�(}���0ޚ�s�=�a4��J�4w�������b�P�����0K+��I޳�pg�y�9W��TfV�y%��Z�J�0Y�q��!^8���e,ſl���F�T�QT@�ބ�(�w
����ɕ�B$�sYl@��jA��x��`z�]��` r:M�_�U�K'����GH��B��8\��;�녂��Q��W��`����nh� t�Yg�iB�U����pɠQ��ekpk3��<�Sc,�x���%����(ߧ���Dog4x�bܢ8�|����I�7�%�~^�Bn���@=kSPl�+�D��(׆LUPc�݅�u��#]D��&����?�
����6c��#�'.�(&���K�Ԣ�RM�S�餐�������Ƃ���H,T�T���:����{,//����,��_)�����=L�)rs�K��)�ϸ-�2@C�u����2�1[�QB�^��.$x��H  �c�5NY�m�B��S��;�W��t��k��T�˟�(w��"��Y�/��=��#�U|>B�R}A��a�V)e'	�'`�[�q�\8Np�UG�x!B��r�@1	��gB����0�S|���ס￪C�!	���f�j!������~���qn�왐��e1����6-~�{���n��;R/�T�9RF�l��ӵI��y�V�Z8:]���b=>r�����҃q�g���{��߿2
�X�XƀALg`�
p���j!>��Ѯ��D슁]tC�M]i���'��:����ͮ�&�7!������)��n��KJ� �ȳ� �f7P�9�8���G����X�8�z���(b�YB�N�gP��;o�i�TփԊ:"�\s'-�Yt��1�ܬ�Ӭ�/&JM$��+Rϲ,R�U���>�i�c�4-�yz~
[��^�b�-��&��Y����/��Ns/���PSb.�l�J3�M�+=�`E�t�b� �#��lI�l�QkC�!6���~{.Y�L���ù���U�U}��߿
�gKTI��I��1|�\��Iq�бW\y���q�@I�I�0�g�����L�� <��dy�����+t����t����}���0�k���n#�h3i�6j�+� � :r9i�.B�@W��%F�%��	� ��ɲV�.��FX;"M���5�!W;s��U�9GB���[o�SO��3��I�կ���9+�~�!�L�Tr��$�ݭ��j�g��B)����N0��3���)��/����$��t�6]Y	!���A������9s4����ֶ�����Hd�� �҂��|�[X�"g=_	�a�/����
�݉*Kh��L����ٳ@�^��v��4n�G�B��������!��AaP�6� q t�������8qRDK������N���&�i�˳��������������C͝��EcEIz�y\w�W���	�p]�Ly�v�� �Hx1�*#A��$�����i�5��_��׆j��gAe�@���Pʫ:����&kJ@5��޳:�NrZ4�{�gݷO8�����K�j��vwsi��.��»٨Aܬ�hAP�W�պ�{����&�=dH5���7V�-��-r߼XK�\"J&lΓ����W}y�U}��������8����X7���0��,���hX�0����ܝlw⷏"v�̝���������NdP���QQ���U�F@���"h�x<Y�I�A���#^X�$�b#�BB��(�!��U4l� ��~*����Su�`��NKhDx�0�yE\k�ˊ𝺨�3���.�+�$?��@U|���4Y!���7
ܹ���c-�=�#�<�Tb���k��NC(�3��۫�QM�W���8.���f!��c̘Qtr��n���O�����XU�Qnjf��O�я~d���(5���F| b��uz��ij��U��hk�pj
�-�!���y�D�z�.Z�/�°�����pt�L���^��ۛ�����k}!�����C���Ȍe��t�\Dӈ�4�b�� ��G��͌�H�{%�9� ]� ����S#�J��R���f��1�y�p�	�3PP��'?9�͝;�`�����Ƽ��Ƒ����(�~5���s�	M��e"��"�� ������Eܰ�#m���g_��歷�u��Y�-��d��I�^~�E�)d�u͂��S�h"܊y7z����&t�R�����{�]��������O�9j���B�4zo^.�s�����x�����Y���qǦe�Hn�_j�!�\퉍in��+-�UE��EK�Ǝ�!��6w�N�D���m&p��]>������s��M0,�� �̠�{X�˴�/�	��qe����������IR�[G�M;�=�?����;�O;��"-���H
���P�v���F�Ϛ=�����#���(sv��$�,�1:=�r������������^L�z�lZ��7��2Ո�d�AZ��=�G�ODU�~��¢�i�K���+u���df�a��E)��K���5�)��&8?���F(�8E�1������ͬ�-��Ӧ�iS��I��jM�Ƨ�z�����t�n���w�XR�1[D$Zz�e�`B���US�'[w�bC\�j��3ڕ���9|ʌ�Qk��E�q���$o��`�׷ɪ�R����W��Hx��`��ᐬ�P��x=/"݆���%P���Y�Pus�!�{s�;��oә9�p`��z�s(�
ج��\@�Q�້r1z^����*�ɟU��$_��)�_�[���q�w����1�W��'�oe�pEи�(� ^=("�H�����y��Y٧b7�Nϫ@Xo1aKܞ�-e.���*a����6B���NR;��o� �ؤ¬z4����~��;�Z��g?�����뮻��C�11�,��u�I<,Z��8	����k��A��Ç�5�rԚ��ͯ/t^x���"�-�dS���FۨѼ���kaa�+AZv��j�ժ^����@��*�Z�N"��5)�b��e�b�{������]zɟl<]}�|��˷NC�ۍ���S���>IJ�YZ�� b>=�z��a|�c��}�=���[oqẺ$]I�,�a�� ���k���"dEI���Y��7���ŤH�o�bn��1�^}�^s�wO�f�ٳ���~�)�p�97��A6����2f���Y��1�n�ȑ6s���SO=��z+ҹR,)������[�k=���X_���[��=�i��@R����Z�~K;B>��k���!q�7H>����߽��[��+�q��ƩL��j�>�ݒR�x����r��Wire��˪��cVX���3����s?�Gѧn(e�=�RZ�����.\�������8CY������:w��GY����� �.������Q���@Ծ����"��n,!�Y��z�֕�T��WGq���®�ۍn��1��'�?��������\XV&,Y����4���$��XVz��k��#��,�#��k��"mn�������p���Z8���~��S��o�\?���Ua��Q�	n�s���/�*]XU㻻|� Y2php�)�UTE%,/�^%������x�ew�Yg�,OY�J§�z+௴y4Q\3�D�[k����2�yԈ��7^v?:���ӏ�[n�\GX&Rm�O����>���~��-⺡�"��5�!ȦЉei��<�p%�Qz������Y�E��ds�I�?�<}���* �B.��Y3�?���7�_��m�$E,����y�Ү9�"ף�̿��f��{�0ɮx� �s��pϸ9����:�'���pg��c,�]��慬�C`�ʪ,2GK��<Kc��2�/~6���O�������}���M@����B)A:��������p��T���+).3�����)�`�О6j���b,G�	�H8B!&��,�
���T1c5�ʉ����C3�A�4�� z�e�P��(�@W�k[Z���A0R�Њ��'�2ބ��"�<�Y8ې:^H��X�֛�ГS�=����v��nVMV���>r���LK�xkF-�{-����35��b?�^�?ސ��0�Q'�x������Gm�"]Ħ�W�n���'��n��:��Ь�=�t5�a�܈(�b�p����8�K�)�n�]�$)�X���V�o�/�N��o����b�0vO��t��?oq�ßp'�sCEf�?���� N�����E�z��ղ�t��xw�W ���hG�kc ��V,����W_5��ᯪ�6VM'�	W�}����p�;fCV㵂˧8�L�S4���%�9m;�����Z]���w��ƛm#v�9����PF���M�!;~j\�Zֳ���N�@2���Ku�3�ֳ~r�'JQ�:t��U'��&�	��M��"��6���D} ����+I���F�Z�bkk}�T.Yw,:(��~ȼys΂e���� -����vh��E������+܋/<�~����"~4��zZ{�?�7�j���&0�={b��	�~���--8kE�>3���na�N8�$�?
XP���5�h�c)�>��qz]1�B��x�+����Z��2|V���(�@Xo4���Hf̘鮻�:��
H�~K }����ݸ�B�Ɍ)5I��.Whj!Df�����mu���[o�6t�{����v�l�b�M.�����lg��z��!#��"�����Qt-*���SB%�ij&LZ>5kw��8��4D@QQ��:m:�i# &���6o��Z�&�ѥ)�*(nT���Wq��#v]�U��)՗Fa�.�]���u9���a��,�w�ɖh����D,>(B�����Y@�*�a�����T�/g��Mn��w���*�`2R��=�/Ƚ�Q1������Gү�"��s3��J&5��,��6e�T�%O�z�ۃPa_b��N���Q�Zٳ��~{qM������t0d��wtD�x��� ��ZP�̡
��W�H
���|>��?�����XJAQ6�OZ�Pu+����i���zҹL"8������d�ZH�w��'��~f�J���so�����:t,�W����zi�(�v�R��6?WD�\�Y����oM�ť��/[jZپ�3<�X�b����E�h�c�����{kk5��}_
�AY2Ѓ�dp~:k����erS�m�V*����\#�b4vYQ�,Ngg�h67CUMt���j0T���~|RQda<��Gq�毈�)BҠ�M�9��a���� o0�*��짞�}w��7'3LA��� [[�࿼R����n���I���>�c���!�� L*Ҋ�I�qa�a-��R̢�asj$�Z�N�4�R�����k�q>4[�{�(lk�6��^q������x�2Y=1>)rX�8����3�A �Hc���͚]�r�IO�>T�Y��d-ƁЮ�3��������+���65@�jr7E��k׵jsĊv�`y'뼺�(�i��Mk"�k��/��T��>Y��ge��iR�G�GvH1B_��
L�x\-	���H�Uz�W�-�A��w$� 2J9� c|C���C��5a����~��?��8�s�����g��HC���6�`UI��?W3�3Q��|z���8�B�	g1m�ұPq��XC
����{����.�wV]�u���/6.���O�(,�~�zF�
��jݸMF��y��ӟ/T��^��C��h�XG�����ش�q(sc`�bQ�(��<�Q�Id��״ �&T��PB�q��S�Z�S���/"��}��̘�Ek� k���>KF
$7KL@9�cg�����v^�nW��<y��!�`�D�D}"ʘ����Z��)J�fs\�iX"�����]������*��L��v�c_s��q�̙k�����O�=�T��2A���uN��)�(j�PSH�[v�l�a&A��ڥc�����4:���"����K ��@W��r�R?����Z�ڊ��T�5��� ��ѡ:N�P�-C����F�y5j�Sm��3I��:�t�{My�a�������P����$���+����XJ��\�s%b ,���_5��7Z�Wo�
�^�P���r;�8Ң!�^����T=��W41�[����=Y��Z�r��Q΁�E�	'~ǽ?i�{��Ϙy0�[�]\^9(J��y�3��}Ҹ��udݪY���;�K�ձdQo�?�}ĈJ��C4ޮ�,D����#1n0)S�� =8�a�� x�M�3�cTI�h�n%�����_���]?�J�b���;z[�W.@r�g��ꫭ�kP�w*�j��-N~�w�4l��jCtb��R/�I�Q(C��o(���3�Ёl*m$��[m��K�;}���%e�U�+	�k�L^�%��A*�+Z��Za��"6�A"���]�7�Œ��Tde_��]Z=1*jjw� 뽊-�k�bδ ���?�!�Oo�|��_ oɀ@b٢
��̍�9��.k�����矇/?��k�X蜪��-����RbdOP�~��GA<DmbV�� �X"�8����L!���[g2ʣNP��V{���0V������~��
�ɵY�泄�����c�r���{�i�e�UV��>��'c�5M+�3��Fa�H�Tǒ�\Y�nYLj�F!�:b�0F�� �U��k���O�6�^��(��������i�f�\���_7�Fd���������@��ޛ�u܉�7��-�:^�ɫWı0
���J�fqЖ�nb�٠.,J�V4n&Ż�qJ2Ɔ��"̝��b�f�� ]�UW]����#�^JW
-��u�<IqQ�;yT�y�e�1v�VW
Q�D�\,.Z�0�U=C]�A��3&=Y�^�AAm����S�L|�ID(���{}�{��6�T4^/�p���v��Τ9��\�������^<�IjZQRĚ.m��toN�7�H��x$P�D	����	R�.PaDj��o�!~�mwX��c�񸪍?���������ϻ?;��`����ϸQ*���&�`UNi����J��OfI$�눗�Y�V��M`+-�1" �z֥<��bۗ���v�"�~�qu"�V�@dٸ���~.�k�q��|���u���,QA�Ε��|X�"h�R �|��l�� t�t[o�W�E6�%K�Q>��"sE�>hb[R��qױ��6_!�,��%�R.?	�[__Y�5�%��|�f	����W��S���ON����z�h�ŋ����F��v��ñ����dġ�0 UAPKa�igR���	h����&qa	��'��N��g��-��nl�A`V�6%���{U8߇�}ёjY�m�L�d� (���黇ӲC;$.��#c���x�6UGp	e6u�n�n�(��U�`��mm��$������?]�G�5�����������ڀ�gU���:����8�p��ƻ4O=�n��������`Y*��^���e1]؏O��m
������S�����c�e�����du];l���qǭ����ݷN8�����v��eV��v�����X��J�۵�gˎċ�&��eqg̚�`��F��K�?�ݶ;�B[n���@� �`
��&���E(�l��a�"9��P��"��0vk���VG�\Y
o,�f�C�z��W8�*Hn�bk�#п�i�K��yXe}4F�b5
RO��.�&4����%��/��7�~������BI	�w[|�e{eqTeo���lh�v�e���{��H(��s����!=�l�4�BY����i	j$8�l��0�nc�j��R�eb�)�ҷ�W���{��g���rI+�-\Lk�zq~����3)4��Vᓩ8qe,�v�a���B�Y��˸v %��&�
�:Q���P$@�e�m:���o�ߧ����"��C��"���W������	$�ѐ��MP�\U��n�R{H//���Ґ�jB_�������o�;j� S;�z�u�ȗ�
D��.ǒ���ğ%>a�\
IGP�t�D�N�˛���j�$a��rۺ�Yc̦�Qb�rX`F}nEi.-�Y�o.8�m�%s-����R��j�fM&�zZ8&����8�jy��0ZD��T��1bz[��SB���̪�rA����%�CQ{�,|�˖DN���$��W���@��������DG�d�w��������q����ݐ��/iUwL�������uTZ=D˃bJ� �A�;Wc�K�|� :��O����w�{z"m(�'��_�op��ʴmu���֥Oܓ�a��b�ѯ:ڻ�`��|kYs(;	��B�T�j�<�kE�B�Hm��r���h���a?LV/�^M�~���_SW5�z��O4/����1�nG��N:�]ݕ(��6�X0^��y��]�Nj��ڠ5�	9��=��b K��a���A6�����a��$du5�O�_HPREf�s?�b�>�լ�:D��h���y�(oUqx���Ĭ�Cݷ�}"E)��N6��M���R����&����wߙ���A%�ϻ���2X��rp���0S����=XX���8����oD.c��h�,�G����i�q�s.��@�w��~�QǸ��}LP����+��6��Le�/"���u0�ئ ;u���A��[��F��/#�6��{��kt- �N�F ��ڭ� 4�j7�t�e��?�|�|��>�H�Q�}�"j!�_/����;�����#(7����2xj7����7�'^��Ȥ,b{0����W��\����JI�P�q�����>���_,��;��g�?��/ę�$���1�� �e �nZ�琖b�)�:2�>�h�.�^/C����۸���X�1���~�FcaH#W��=ߧ��X%�(��.�v_������y��~��C��S��F�gc$�{!�s���Wvw�B�޷}����^��
������=A��E�,#�ݎ�Q��s`�ܾ{���ݓ�J���5��oE�c��;hh��$F]�2^�B��VЯ�L��<���s��m�w����p;��������<Їe���"ReW(+��x�7Yh/[����V=�"��M�͡��ou�����/�M��Q��T�%%hSc��=���=�܋�F+�:F�C���<���f\W-�k���"�!B����t���D��2��J�v�F���:���]|���o�3���'�pw��6w��?ucF��F��[#��3�ޭ�%dy�-����.X�T�2F+ZXᛄ봛�Z�~V�Xq���o�{�},��ю�A�����|�X�]��FLQ<7�3����,���*bU(f*vʤ� Wt�-7w/�����OJ��D�Xv6�z(�/+gI�gi��
��2����e��`D��ƿdC~A��p�ZZ>���8��V[��hFQ�s]ɆVb�3?��/l��Ρ�L�����MM�
�?���6�5ױ��:�Bl�c0&�1��`v�b{� �P�7�r���/�u�}�Wu��٩3HSFؙo������c��o��)��/�I*��gi�_��.l��Z})e�2����]S쒗W`;.$�\�6&'χ�&��ŝ~��V[n�b��!�Je��g���P���]1���5�!�	 �q�w �f��FP�ea;�� J�2�	%������F�/�^y�c�V���
���!:��\v���=�ԃ+@i/��'�LqԂ�-��^��������\�T�&) �������b�?�b��ֵ�I��M_��0w���3qrWg�H)���s%����1�m6a��j��.[�"�*��xU�5v6���
�"u"�>�*�>�=�HR�{��j'C��2q�+��+|����6�*�	`1�*�XK1J�,�������L&nQ���̃}�ڿ�W�ݝ{�ٖ�j��&7)��x�Q]���^��� �qJۊ�B� d�B��p9cF�+.��\%�����o�f�M�+�;V�y��cK}�,��/�@(L:I	7h�/Q�]|�!r��'J[��B6>���x���)7�$F�3�p����@��@�fS�B�s��mV^�<�USp��\��|�
âe�n�56v���许`9Z,���+���I_n����!��r��Զ�aW�p9�Zk���-W�&z�5����<Jkq�;��cݠ�ÓВ��건x�@na-��{���S���-4�M��������=�¬��|���,7������/�]���T��΂�KiH/�y6�����"Ga���Y��G�]�����lW3h�}��%ngR�?�q�&^&��ܭJaV&˳���`CPڟ�_>)�N4��/Ăv��i�R�kh�pO�*)�ޟ�n��f�L/d\�xw�gZ�B�0d��~����D���W�W$_��Tq;��`�g�UTT�q�tr�r�|����?���������`WU		ȅ ��s3ϱe�P L��eh���!;��o1���z���P=A���S�@P�����ٛ"&2���߱���|0:$�U=(��N8��x),� =y4mu�Ȧ"i5����|��?��`�;��c����K2�ef�>�FҰY�1)BoH\u��JRՊmB������5���9�!n��^{�	���3��zt�^К껩��i�����
%��լUjZI�O�r���m,� >�L5(�W�O��~�O�z�5J�t���{�?
Q���I��������I������;�2��zG� o��!���t�S�=j� ,���;l0��,u�<c��m��Q���N�l��k�I�,��6+jdTY��!Ns�1"�\\T��s�}���A�D63��z*�*����\c,�͸PE�ƨ�a�����Ĵ�C\���{+(K)� # 4<H(dA!$�X�f�pjց �ĕe��N?��T�,��f�I0�5@a��j(�Ib�i#m���u����oK�:��{�����/ةE��Q��E�퀯x\ǚ[�v�"��Y/�6Q$)IPHBB�6���lW^קW�������z��Ǉ�,Q����
V�١�������}L4�,ϣ��<h+�@#Vq�/Da��&���{ZCS�QHEY�RL�d��G�]w��m��w�y���t0M�"��e	�1hXj'�'zT�T�������C���BI�|=g��_y�|R��Q$ �������u>ɵ,�܈9s����+�%}�Pz�g����/ɵ���kg�!�Yᩘ�2`@�{��ܿ��m��9�����)�D4,E��F� �9{�\���]��!l*���A
<�\AY,���P)��&5��&0*#=r�L�jkk����AF��@�����&��=������hO?0����L��S(}[S_aL�<��6�$����gX�+A#?y��]|���d%(����de�{A�j7k��F�[n���;�����9��2gM�/ fV0h|9�2���P )ݪ�Ŋ�х�|�u.�1�]~��~�	��H1�x�����;�*��$�qs�. -��b�Wz��Ī��/��3l�&��Ġ"�_?W��n(X3�@��w��
�/���;��#�'��,Tc�k�绅��q����E��y�7���g��qr/����2tS�C�����MeKw����E�6�A󻺛Q�����kǦ���zq��o|e1|����.�?�c�h?[�4M}}<��)��S�XUZ'���>��/�H��{��[,!�	��7�][gf��Hgi��K���p��OqC�U�2UV��0WQ�o`? ��$�P���F������|H��2��g1.�̌jb ��ɜ�r�g��������Z*T�*rKTǨ��0h��RX��T\�E~1P��ΩieT�:9�y���}P�6�P�`�#H,7$� �{:����;�`l*r���F6c���k���?�M���h$���^�+V�gy��xߥ� ���)���&V��n{��_}����/���Ajjja�����Rx�
`���fm��ک����j;8lImHZko�.޺���(�<�'�^�g�r� ����UaP�l��&�grS�G�����H!:J#S�q$���	����V� 1�{�b<EqB!�~�L�����F��$>h�D@
��[��"��)Yc�,J'=�T��x������|���  �od,2wli֖�o�=�zE�xnY���3BW��
n`Qn<.�:�X,�-�O�̟�G�5���;nw;�z����\
&�����ߐF>�!�j� ���/�]��B)��u�'�y����r|���k���;�~��l��V�\#>4Pn�9	�/�1�N��k3?�j�N
�$T���ܝuHhn�r��	��k�����cU�!�9;;s2����6��}n
���,CP��Y��)Ll&P�6�`5�H.2�Έ␤z��O�J<��7~�!�b�2`A�?%����ZW��)'@���Pf&�{R
Y�� 0�cy`�H�R ,*���`,���Ϙ�KH]�};�v�n�_+>�^�����{� }1�t4��1��ÈH(�!0�S�1�hb�B+׮�k�^TtHX��?���.m�m��Y�@,`�͋|�����#�4�b�K�����J ead�4�X.���jQ����EW�+`,�D[�n2���r/�Ճ�d]55:McA�3��",wX����IbB~�u\�&ʼX����A'4'x����(��4+Fm���0�`��#fؖ]&$�)@�����%c/�DhZ�\�ʀ��uO<� SyǺ}���U�`5�����đ~u��SJVA>�<�&��e���"CY 3�*]]T�[z�ov�<l��3o��W�믿���B3��=|�w,��&�F�/��)��R��x���k(~/�]�_Ԝ��>+��v�o7�� ( X�J����Q�4���/�v�QG��n��L�Wf����rk��wPj\���<�#�^���5-�,
O�=�����s��]c�$ٜ��Ҁ�@�N�Az�\J�M�R�#)z�#���}��ڗ��`LH�|���6���$�i��xW��(L4�	w��i��>��>(B��H�3�}���ؾܥ�.j�h��M~�G�Y�fN�7�t�;!&ZP.j(Tѵ�vv� �D���Q�jT� ��o�T �,����r��ͨ4c#�%�^�d�,Bi)��)^�`i�<B,�c�<fKZ�m��&a�:��E���/F�H{)�̠���t���~H�91"����#��e����q�r�-�ٛt�YY[�5e�����;�TJ!���knϽv'������&�B�m�:D_�nȭ,"Y�ħ����1 �WH�lJ�<¸�*�*˖�Wl]���j�0�]��V��:�,�j4��H3�Jϣ,%���b������`<�3��&�/� x��Q�f�W��J��a4JA����q���s���w�s���%�F59��y�z$UPMa��y��� �B�y�1b�á��.���n�mv���^�(Ë1��R�����Z�Zn�n��)���e�h��-�Q,�[��B����^/��.���0A*��\�ad~\�����%r@eK�<�J��ҵR[K/[�q5����ʢx0'7�x��dŲȎ��ah>�XBX�:F�v�{�T�qZ��ҕZ�q��4����hQ�rC�uCY1R�"�m*I`��%:���e����w3��C�ܞ���'�F���(���>w�5U��V&OR���CO<��Y�E�&��7x�, @����3f���|��|w��O�v4��n��^��N�iC	�_��|8�r���T�� ����Ag��M�6���mk�%)�R�P�����uR�"Ǩ�FSʜ{@��,H6#I6�,tD��״���^E�c��Z�l��ho�Ӓ��ˮ�ߒ�[3]�2�r��'�{r9�B^A��|+�j"��o���<n�xR�I�HU����g�l��4ܵp��od�9��7q�'� 8��~�~S�NF#��_q������E��E�b���%�}��XsmX���V�яXﷰ�eVl�;�AFMa�#� %�Ҍ&%ɄŤ���vݕ{���K8,h��(ؔ!R*������1�� ���w7\w���75v{��H��H'7@���v���q���7O�_�T�����ˍ� ��Pʲ��Vןj5bH!�I1s�U˟z�IX͸O��S��G�ʤ:N��b��O@iX|8�����:�Ni�	�*��r���[�k�5黋1g�d�bi�1�.	�c8�"K�u��3�l4�I1��-�v�Ϡ!�G,8�j[��ԍ⮼2��|6��|�>�u>�|%��]���V���6b ��.>�/!Lb1
�
3���߈�������0x�����l��y��oa|���W	�v|�p	��p��K��pa��?!��C�p⩤a��I�`3 g�{{�GL�ڑqv��2ޢ��8�������;�U��TL�mr�8(�n���܄V��1����#9�	_��fh�><y;v�0���B	}�]��Sl!�ȫb�TǤ��d~Yv-|������AsY��BK��ȩ��������:���i��	�`��C`GoVX//����ӊe-��6�0��s5Yn�͇�c�>�������n�Gﻱ�����r�Fpy+m�0�Tc3����mX���˷Q�/�OM�m����(D��oi︀���=ˊ^�Z!,�܀���"�1��L�������JK�	���b�bkK����[�G~�?�0����WF戺���o:~���v���si�k����e-�8�Ƃ�4��Ȁ��V�G���s'���|�]��K)2���:-�KJ����;jl]x0Q5Yb�pg��x3,��Z�=.���&��
s��ς���G� �Z&oe2C�3�����9th��ʘ���W�c��#�:Ziz�@�JF����b��O� a�����QL� ��--c�T�ia�Ai��İ�݄-ƻ?�n�м{.�L4Wr�����qCIAοa���	��DI��v�(nX:��q0�|����x������+K2Gk�XV�hg�Cn�u`��-�}�H�6�.�ܴ0*� *�����n��}��'�g���>t8~6B�2<���l���	��9�>e�X�O�B�"�L}ʊ������m�Ŧ�sς��G̋)��4��e��}�w�q;�Ut��e+.*�-��I� �^�Q������6�&{S�oY_�X
;�����{ 4j}�/t���,���1 �0k����P>��?@%�>fTV"o����u��鸞t�ˀ7s����2ml�{��)��Ig����cʂ�ẓz4�� 	�UE9�Sw�h���R��0dL*a�?F��ۻ�7`_�Z�/��������>�D�O��������.�[��n`UUŰ2�F�b�@o*\W����m���`�����eA��@֥(���g�p)6���:W3��2K7�x���޻(�n���ueЦ�w�X?�����{���n`��nUs��U4���x����Qw�J�W����&6��w��W�0�j��-�G��#O?�d��t췯��(ȖՓe�E���i�S�|M���U����Q?K&���3��� ������O�2�S�7����MYXL�K������?X�G��C}fl�Z9�n����{���)����`d�4��9Eu�2��+��E���Y� |R�$����?Xu������������?IF:$��1�� *B��Z2�b��ugX��;o��y�mm���;mo��q��:S�%��&�,$�W�u�>�*,*{���ڏv�FHͩ�iT��0)C>m
���8ؾ����ψ�w����X���NR��$�XI���=\a�x�-�#�>���������kgwƏNmA�&ݬ�x���X%'�r��1���Ms�� ��9p�JQ�A 6[ &�A���J$���o�����W�#�#��8�u.��Yz`	������ПpE��f��ȃ��@(Zݨ�C*���n��B�>d�?�o� ��eɾ	�j'�M����7\���w��3�A�z�Y�J� z�ҥ�r����'�	̄Gᔹ�$f�Rj��樂4���bv�.�Ӯ����'�Y�~����-��a�b ��:��9�r4B��ʛ��U�sz�O]׺�I��\�+;P q�i\�u�݄�:��m�/�V����X���d�����
SW@$�@��d C���8�zK�L�Q'#ac��fX�����ܮ��j�D%�a$v�`a�g�=�~��˦,}�Ѻޕ���r�F�)i���k$�l�v���\��V )0`$�>olÊK[�ܧ8�yM\޳���g���t��X�y�U���
�^�"h\���D�u�4��CbA���������,v�u�B]�`6����L)8/�M�b>�Z�`6�di�.��.��M���=�Н���n�A�hzSA/*�lZ���⬕�2��nRI���G_�K(�i���NO��*�f�,�����y4�|�Q��w?��C`�!���L�4��4% N���{�I��X�q�yt*�^Z���6��)	"������	>���)������x��}<����n��֛���x�xɱ(����2Ų(%�Y����I�Λ?�z/��XRy|�yi�����ɇ�hI�%WK�Pt&aI��d��FZUqA3|g�.�Ui�IJ��I�X�j��}����c�Z��!�SA��q��8�}:�&̜M�Ҕ-�$wG#u��ϧ_���Otg����_����~P�Q��-Jks�g�u�z�_F�IJ(#a��	���A%w�����ß\���~o����@#�z��LY�;2\{3,0���!���*a�ϦL��6t��cݯ����j��7��Է�N�)`��1'+���/�ނ��b�9g��E�M�������С���^DP���md�b2N�j����V����kғ��J��AYf�#��nJq�b�<
�;Q$A��q�[A���i�aBG��f��n����a&=#s>Ei��,X��I�	��E�� E?��nbQ�%�6�b�V���̸��UTu��R� D����2)-YgRO�WH�g���2<��T0A��C�yӻls�u(��3A7|��jd�kh�C[�'Ť�I��r�{���ݵ�W��r�� ��.�e��".��y�oS>��fΘ�a��Z3���S@P� �GC��Jb'����L;�=3=cޗPW�׋���dr/���|�?�Л"U���I�.q��w����dt)�FN�(�g�n�ճ0�կ��QY)�%ER�H!yo��KA��т�H �L�U�����[m��p�?�Ũ��R_�4>���@o���?zB��6a��_8�K�����:Dazw��"�2<f�,�i�.w7��
�	�g��h�������� `�$�p|��X�-��T��.�����3dq5�x���.�i�E��;�j�e��Gg��&�=��Ӱ�d�U1&�5405!�$I	��?��z�m2n�uN>���������-��wic���5~���)����Ea�v�#ع�䦐��}���?�2�9��+���;��.뼠�\���������2E�t.{�30����q6�|2sj�T�A��;�y_7٠�(�è�Mׯ{�H92b(��Or1ľ��ݺS�O����K������c�߅�xPݔ!iU�a�u�{�]���g̏t�{��[��*RBa��y�w�[K/��f�1F.�zX�DM�0�>W����5nނZ��L`� <(>.4D�_rsm�s��Z��3ϳ�gr����fj�'����W�r?�ᷓs=���f��yW쳴��Ej����r�]28�s�Z#��_��lKI�\��x������<�=����T; ^�[�-�������T�KV�mҖ,���]�%2d~�W�H������o�jH�#E WsN?��L�i �X�44~A?kzv]m�PEz�S6�3��_���}A�~0߉icy4�(���茆1��ĥ>+�E�Ol��L�R�&�`�BR�%��Ϋ�+V�������f�_ݍ��J�����U�Z�C�os��>���y�J$<�G͈�G�d��D�G�jW��γBnH���J�P�Մ�N���2c����Oq�I �$*�b��O��}:���j3ǧ�s.��1�]�K{���AY�i��OQTV:<#�������{��8�Pw����c��`���j n�����G��v ���؛���au�����yʸм$��6pY���֌�S�W*�S�4"�o ��R�b!H�l�i����E��u�n<?��|F�z�� ���wrn�؈��λ�u�5�������Y7{.P�)hG��$����t]�fӜ�[��H�.ÿ:�U�S#V����D$@��˺-^T�u�Q��'�l�(ru���E�������wr�����U�	�|���}���N�\d`��g���ޫ���d�JZ�t1x�ø��Qb-L���-(�8�B�u���ē���}�w�y?#�\�!��l��2�d!�@��n�x8Zz�㏱3���+���:Y��Y�-)�:jޜ�cG��Z�l��`��؏8!���&WVܻe��-d�A�1�L����`��&q����2�&��<�D�O/�`:�b�E��*�'�	+�IU�$��g�ƫ��vx�bR�;�Bs*�����{�����w���(V+��`7B��c�C8(�h/$��V� t��p��d�3�[4��w�G��j#� �h�㔔�X%m"���.;|�����L��F��/#�L��x�d*=*�d{�	6!�m������Ox��c&Hs.����u���^���ϧ8��{��Pp�j��76��#���X_���0#��m]�kma"����c����C���A�^�~��,v�?p/�}��_D�`#�\Q�Ƒ(�0��0���[��w�k�ɜ����L�������@`G!����٪4v�&:-X�U�W�]M�2�fՍT�!�KB��B�y�� bK���~�,����?�)|QA��o�p��5d�dUh�c���	+
r�Gz�
����B�b̾ѡ��&L��m�I���^�Fn�6}G�n��1P��B#�������UFK�|k9!�ߟ7��^����%R�}k��U7)�� -wV?��6�s��vv�^z�!&�I).�D�D��s�
ʲ�
Cf+�z�o=�x,��h����Du O=���s���mI�	T�X���H�@x��\F1MK3B#dvH�#P�^D�&���n֬iHʰ��V����j����VY����V"�Y��?�X���h�$,u�	�
t������{�v��?�9���ΣZӕ�/�+�F�U���&����͘e×
�ͺ�qƙ��od|��F��T�>J�*�m����h#1!�ʠ@��3�L�:%o��_��oy�]z5�K%��U��_[�^q����$4}JJ�+FR���A5��üF
{2�D���ıV.�R��{�bg�w�����а�v�t�2o�T_�Dh�k-�q>��.+�� 	�ܕ6�z�Nr�ʱ0��,9ܘj���8�?R�x�aǲ(:������/�X�1�x�[� �Z���z�-k�*��V�����nQ3 kB���S�g�n��{�*'8����W�8i�<7ѧ2e�L7r�x�D�n�M6uGq�e��*%���Pԍt2-R&ѪJ�Ȃ5����7�xr��=t���ۤC����W��x��%��d=G�~ba��>	��BV��h�I�H|���b��`}�,--�-.�Y��?�8�Xa�������.{nw8�S #+�΋�N7�zL�;�
W/�w؊���{���LY ���v҃��@ a���ڇ=Q�l��X*�����INaz�ݘ�ܱǝĜ�m�B������	�b��[�n���.0����b�b�3��5��>��͘9Ý�ӟ �����7�%���I8�#z&�!�w�3�
����I8T�N9���޾�ڣ�(�n�	�Eh�1�XS�2��$�}�i\�RC7��*�X�W�|M�Է!��k��^�
c��YRaD�n�Ĉ>`�/��Eͣ�xq-=6ðvX����;����_Æ�\�d��W�X#�!�������S������<��c)�C� ���X�t��+�Y�5;+ ����#�=L��B�p�-�]�����w6���U	�6K��l	�n���f���oOv���,7d�H�ˉ�u��%`��"�&�eӗ�c�]�S��ޒl�LR�XU)j1)UӦOuÆ1��0d��=�������FL��\[���Y�p1g��9�v���n{�C�osm4υ5&���\}$~*X�+!-�S@�3>�t��s��\C�"wԱ�2�����28��9����	Ȗ��8��&�XD��k�[��,��O�B�Fg(6����;�WV�ؚ� hFa�0����dff��|u�5
���,Ʈ�Ivf+��Z]s��Y�9B�=j�y�lW��M�m8nI1c�j�����!�+������Iqubl�mbeXR ��#Ⱦ\��6�����]wƙ���?�]���ٳ !k�(��ٍM���ۡ����%(�:|�@s��A��)��b�QF�1AÌ�u�^|��t
S�n���w�Q�7l�Z�vT��9��-M�iZ�-"��Fd1�b)����VʢxF0�<��a�|�Q��@dq���qW��R�̳���l��:�"�k��lf�fgt&9��Eff�k#�V�IߺHI��Z!P\��)�m��ͥ��<���US�,V�d�+��XB��';�9�����%��^�6�G+��n�9�e���ou/����)'�eq����?�bN7��ʌ	�}4=d��9AC??;C�}�R��?g��Lq�U��D�����;��߷��4�t+;kV`��D-+�ӿ<˿��e���W��%����TR�.���7�~�qYV7��^���n�}q���q�ͫ{��u�MK�HqT�7$3Mr��oIQ����q����xz|?~�t���p�Y�St�tG�V
�q��
����Fkj�G&�/=��Z�c/s�_Ƿ(�w_�����u��sqfFƣ�#���wl����ss��YVKa Vf��9��#�V����YV$�jtk�����f�D��#�~�z�w�ݷ�+����L/�Hn8�~D�L����zL���Xa��4(����X��܁�0��s1~��q�%
[I1q0@	���️>�ȝ}���^��Bh��[���䙒��jo��~�f��h��T���J�`�7
С{��W���TEۺ���W�vƨW�o~�$�iه�/�E
�u�d��f�M�����ē��&}�68��X%�k�8���Hʅx����z�@*\Hr���R�l�,^�E��GM��� ʚ�g��GL/_T��f�|�DG'2�*�Ŀ�|e2c��c�6���� p?d��@x,͛_��RB�����^Ћ=*�A�]r��-�7^�}�~����)M�q��"��P1�͢s[ZfYFH<���
j
�#���l8���|� �����b�x�ן��s+��BT�pa��l��vM	�\	�/�ǏV6alu�#���߻�x�t��gV������k .�L�L���x�}<e&�(��`O1𧮭�
�vz�P�^��}hm?����}��ܿ�u���IGC B\�&T6�!��6�/�&Z:i������9��o�=������P*�~�@K1$$Y�U�zh#I皆��5\ڭ��=�0�Q��u�Kv�V&��}W���ꞯRa�Dte���F�ې�5[�mR�����!����by!���D��|�hL��&果g������Ů����E��&�b����2��H�,+���D1:�>�p����1��4f�&�����L�/�o=xpJۙ�)d��A무�;v)s[Z<ί�++~ztFIuY*�F��C���50�Pܚ��Ƶ-d\�8¬HȺ*U�K�\�C�T�=S+k���a�F�͸3�ȋH�*������ZEH�(qB:�$J>qc�Y�\�^����W7p�(w��璘)"j�,��i���'ˤ�p�ϧ�!����䱤�dX�bR��-��������\��qU���}�
��vw�6���wGO`�V�n�W# p�pr��F;�"�M�b����ɚ�j��ߢ�y|`���}ÍB%��+�<*���8z���Y���&MiFV���촃W�����(���4��%(-^_)�� ��5�Nc,��|
�Pк�
�dO}�R�r��U+�@�R�WMX�r�4I`�~�U(� ��bB�c�Ÿb�.w��\ϟ�?�� W�O�7[n�Ă4�%�m"'� {k����*��>A�����}�e��=��h������H.�&B�@��e-(�1�$d��������͹��Y_�,.��,��˲���q5��rq|��E`b;�M*-S�_l���0�ͥ\r׀��7qO>���e�}��'���v����N��Lm�W�+��gf�K���B������*rfgkJq�{��g�ig�n���U���� �;:�[�)�oa��u��yu[�Wx7z{���{<�d��R۵��a���2�fjΫ%]h�FYG]�׷����Rx�#T��g��c����V�tc�� b��2�tjB�������2(HF��;���q1�0�m:������c�����w��3}o���S�M��S������~w��ƯT�ey�}�
�V� -�]мƇ#` ���)��!&�����iv#iesH�T�W߈vpM*���a�o�����x,H���^tC��s�w������b�%� �4^e@ ��n��M1d�X��8`� (�*ݯ�w·O���Ĳ`z̚E\T��y,<,X@j$A�X_��$��8W%+���DA�J̾Oi��1~=.T�e�����y��D��m����b�����vQ�2�����ӹR��/�؍5�}�Ѯ���
����`�r���7GV:�H�/��i�N���랖F��!�Pֿ�]����M6�ȿ��SO=���A��V�GiyY�e�%GFqyp�O��fL�ڈ纬�=^�+�0�����4�3ͫ�H�)��^!���`W�.i)[n�Ȍ�oJ�jG�>}�q��kB$y���=�=���~Y�w��?s�?����)
I7$}#apW3fΥ�	�ޖ[��w1��C�~�ACh���6����t��r2WAY<b u��n��Ǹ��?�?_�G ���+���=4[����q4�crzX�A!�����{(K��o*#6d)4�@ĕ�g��\�!��v����;L��ӧZU��%Ul���o��?>�Ɗq�-Z�2ISk�T{;�7ݑ8�2�6��qtbe���mc�EU���-�ֽ�m�̝?���-e=�p��[���|j6C�;��V�J7>و���Xo���
�˯�����KQ}c���$&���ħ����%@��o��ky�\�^*���,�K�ڛ�;－�d�M7�Ԉ�5:���H�E�"���s���������a}$�L��(Y!M�ta�\ª�~���nۭ�p���������믵Z��8ڣ�%��]ՙ��o
'֙"H�� *��f^K�Z��H�̐yk�M���_�<�����ۚ�y�~|�,�1:p`��m���G�����K�O~|�b5t- ��5�%�iaS!���ZZ�,F��N��:�M!�Bs�ƎG���2���"2�E��>�.����_��~��( صN��4^]ir0tL�G��E�yo���f�_wN�/��-#��\2��Ohm��5�#��z�{�gm4�XF`��[3#"�����JJ��\�mx�����޳������]ɯ���;m��o�=]]=7��s��L���àX�ޫy�F{���B%+"�]w���y�ql
Ҷ]��h�};�)�v4c�`��i(wC��Q1�T�}9k��PWH0�E���K|�^��Y>��g�u���k�{�r.�7�¨R NY�K.�؆K��'?6�3l�����,2p�ط.暄��h�++ԨB�(Tb$�H�9�s���L*	�; ��Y�9li�������d
�?w��͑�����dv1x��;;�\Qq�u6��W2���4/������=Yڽq�U1��]�U�}M��^+�n<^ss����Յ��g�},0���O���н���|�A{R�X`�<u+��zhR2�E
̭�����gW>���r�����_���$ �%F��6�B�@�y�,8�ǂ���t���sx��e�+�����G��Rn�,��2��%6����W�%kem$z�{��OY?ί�[ܱE`�4�.���縨`4Ph[)��)��.�.���5cRVA�?���w.)�S~A��ɻ�?��o�Ź��3>�>�VQ6��x���M_e�5��z$��u-�+vU�-#�h�����9e���s��Ak�)�}O=����^��� W�����w��^}�Uw�]w���3! @c��c]��p�Ԣ,AT9w�AyD��n��kq!7�	Z�[K�B&h��'�KK������v�0�� �C9�� ���ʁkTF)d#��s����
�V�WrM��ykl�`��;j��F�kۧ�x�خ;n���u;��Ǿ�����X����5�u`-5���>}6QKe�ҥ�K�J`�$�Eդ�O����^�I�[iY��~�]��?lԝ�r�򡉍v4���=4j��ߧ%z�a�W�N[;�����p�l:#i�:��娌��2�i��x��˻�m�zDmk{(�nBa�\��A�4r�z�QHksm��d��%��-��o�ۧz񕧢���1Sp�yb�<L՝w��n��u�GH,��>��r�*�ԍ[�Юk�fDw� �	S�ЊO���a����;��H@@IDH!}�Jn��:
�gY�t�z-T�����0�*b}������C}c����)�?��q{�Î[0�H��e-k�q�X�����uZmL^���S��C֤��`2�������,s�{�J�9,9��D�Z���]ZVT�HV ���{l
#&��54����;����R=K�.Y"����uT1�����A���`�������}6�2<�>�5k�e���4e����V�O�"hW��jB#Gq����o����*�6��D4H=�n/>�����j>���V�B��駳��=!�Xw�1'��}��gn츱 Zmx�2�r,��;I.$_�z�&+P�#x�� �J՗WFO�Pe.V����/>{��n�m6q��7if! �^!H1G2Բ%!Ի����̡(K�4c�S�(���c��=�H8�_���l�l64��F�]2�"�ca�K���[��0�D)��;�0?��qnj�pb�6�9���]���&�5��%�'A������YY�Teedq�1��v�d߸�%����̕\'Y�Fg ��]w��F��F`�\�VC�U���}Q	�L�g}�bܸ��ȲI�h���{�Lr���������O8+�Z���%7O��,�ʃ�e�7�ZY3�*���XQQ嚱��(H��fƀ ����݋/?�0�� �؎k�v�R�-"v)+F���-cL9��7ޘ�y4�Kx�=@~�]p�M��Au�}F�Λ�$$�3e�1��W��0�&��ԇ1��x��'2�����i����Q��l���uSend!<7ë�S����;'�o	�_K��	j���81D5�[J���N�lX��M�Y���r�qCrkP��b��ݵ��Q�5�7Ȉ�⛞V��c4`\ȂRCI��5��W�tO?�H�*w܉���¬�%[���@)\V�̦�B�9�fi2���êeB)��h�v��չ��u+�zϹ����7n43)�1�U��Ω�H�4J����o����H�WWt���I+_�|�n���{�"&d�z�[UYzY��U%%_���ׁ u�m�Ͱ.'�~�5Ԃ }idMda�+�"$GdۀS���쏵�d�-�AJֿ�!�0UUU���˟|�ݸQ��w���P�x#5�y(>|)h�vI �*)�Re����t�
�D���� �H:�H,Ұ:t�����.��fw�q'�-����)�,�Z�����K+E#�g�m�2����'�%S�6���P4	9Fo�5�;mn��&�C=��Q�c��A���f�d�Pr�5r��g�ݿn���ʄG?�ۙ���.i�?Ҫ���֝ad��{g��j$;� :�HN�ŀd���Ў���Y��6y�~s�v�|p��A�)��va5Wa-q1^�3�=����X�T���������1�3��N�A˦kTG7���(��@��	 ?���Fi�8�)���i���]l�?���O>��&K�3��������O�RO����q�����w�o��	��"Z nv7��kȓ���ut�:pm�MYļ��G�`y�wZ�Y0�)���ZjB� ����,���*��!���V`�vg��0 ����2�m�g�iMr~q�T�X�c�,��!=�M7]��^#T3�̇|X��jGAȱp���|WZ�T0nM�LW���y.��<��c�D*y���	Ū���&NI��2��ѱ[� Asayd���j�~����?�Sܦ��5fL�*+�0+��+���I�&ӯ=E�+�������xE�Ґ�����{�m��6��cq�fϲA��e�"�c��@[��M�8��(�4�]Av�]&*����v뿄�f8T"���I9��+26���ن�p�'���p3,[˿5*�W��g�_}�F���!�L�1���"w��2�����{<N��n�& �Y����6x�3�7����@#�Z�o�R���N�k��1�g�z�$�ؽ��tWg�2wr�>��w�w��]xQ2�Z��_�%[W��uѨp]���"�1��*eJK��w�<y����]����n��6����Vk{8��c-]����F4e�+��tVfB��ѿ#u�#$
8rӮ���Hlf0MC�L7�,Lt�ݼw��翈Vq ���2d�4h�p�B�O�'riP�u��7y�gT���ExG���Н�O밬MDd�0�b�Ai�)h*0�D��C�@"+E](���^��H�;���)��i��f�-cF��,� =kga�����0�*C�� ^�ũ��Smm>#J���Od9>�=��	j���o}�2cǓ!\���ȍ7�6����C7�M�P�T,��������O\����+Q2��ޤ���H~���)�)P�ҟ颛�Ir`I��z��U�J&��y��]�C����j��Ed���%�Un��FЪ�9?�c�C"T��*(X<�FG'�ap�7��N5��~$��0I�%�q�6���-p�m���.S�Nu����	��ܳ�ˀQW�¬Ba4Rw�S I�������ޯ��;1�$<�+��B���:@wwџSai�+�����;�`������@�'�)z15�W3ҿ:�|k+�+,�0PH+^�|ʲ	;�����Tp�v.뗧��T�"!ðB6wS�QA�f-��j.��`�$.S�"��Eذw�}���ܡ�v�g`��6�x�Ś	O�F�iLD��КF�#�zuS�]�-A���L�IA��S6�Q�������Y ��R�Ko�k�0�M.#��:>���6�sҭ$�����ses�)�H*]u��v�i *˳>%NDW��'=?���-(�y����VȾJ�[e��L��,��H<�#;�~<Ơ4��S�eaVv�U�Q�~9-���*�����0�OG@U�S�4.Qv��3z!�%���*���>���n74�~t2�4��A�h���Y���N��@O7H` :���o4�1J�N1���s��Pd�$�=��g���H��W!��S�ud����b�x�Q}��擌�I�,�Z�ðovc����C-�#d�eц$�hcI��eS
O�R����TYI�5�.P��Z����u�T�Lˊ�#U(�H�m�{ KF���Y��{�S�����:Կ�5kqyGR(�f��X
C��Z��D�Q�[;n�����6���B�c8��
�%s$���1C�q���y	q�"艨�/^HO=m�r���Fo��?n�}�w=��Ճ���q4 �{��@�A^�-�:�Q��hR��w�a�mK�h3�:��e���3��(���c���!N�J���!̜,J�U�b�$&�߿c��9=�Y�Y?i�S�I�kmDҡḡ��z_.//)|���+Í��۳���V��HM�P�K�:1w��"�<!(���w��t�y�.�}��(�4�U�Va���!�������I���{|[T�7�'ő�/���U��40��g�d���Fy{|��L\�n8�m�Vk�{����Mp-��o��;��"�t�£����qb�,�hP3k
@/�-@�@�lUz���Ԕ���a�9Y��=ȍ���'��_38��oJM��F\֍[ŕ*��'�٠ǂFP��$�\ݠ�U�U�dL�{�=2rY�S�&L_B\h��E������8?��u����W �+������(M-
3#���I�'!7mW~7��j�J�?E�*�}��z�lJ#��/_K���SϨx��:��s7|�>p���d�U}=S���|�!n�}�v�=��;�C�����eם�Z�I:QY6q����Ko�X�i�f�TL/��j#���A�:d�*+��C�?��U�7pS�s�@�x�YҜ,ZkS�;�Q��X��J :d�ixmVok�'�}�}n�e��=�
��<���w���nc��tb]��j�(��������,�|��"6�a(̦(��Ɩd.I>��.���mI�c�&����d�K���m���Y��	�_����[VQ]�*|��$i�zhz 3^s���?��~�5n�曻�^~l֦V̃��Gg��5k6��\5YV�O���ZHN�p�-���rS7~�Q�N���b��XZ�}6��6q-k��������2�J�|�S�&�b�,�&�o�P�����A�w��Y��뗮�Xc)=��I��^P����ܐ:�RG�Xg�ѹ���+%)��Hq&  [L�ߕ 8�*�t��]C��䖬���At��x���JyϚ����yxٽ��R�b�om�����be�l�0.Pm�BXm�X��K.��i��\�d�ZܓO>sd3���ۙ$\M�"�각ʺ�����`�y���\2�c�\s�����f
�^&�A��|P	8�)�P�d3��21��� �k�\��m��~a�R׼te� kP���v-���(������ɞ��X�+����u	��vX/
�x���x��b�h��[*�Ǝ;��
l$~����ӯ�2V�0^ �)���N�}B�L=����@E߇�ue}�QI��)�~V젱�>�~��UW�ͬ�Yg��~���������L3+!�H�I*XJaZ�����=J8 ��w�y�x�����Π�1�����\P;�U����	bSVZ��7a�7f��a�ܢō���~��3�&Ѱu�%� L}I Ͷ\
}�E���ϧ����U{ '3m��
�W�}�Ua���@��̖!Ã[Z���{"�l���Z��w95�\�������S�(�U�?���N�щ�(*Q�gg�+�܁P:��t
��_��@� $ˣj}UU.�������-�M�HC�Y�\4�q���n���5��[d�1o��F��5
Z��� ��/~�3���t��ܖ�r���P\�K)���u3�SP���S�`���o��,V�;��_c�������ŅT���,�u���I �oI��azP8m\kS �� �������{��1�E� 
���d�׷�(A?w��;����d��$ٚͪF����d_Ri�y��o?��u�R��y���JLp-���X��̌��lx���b�-�Q	�AÄ�'!.�-��i��Qyb��K���N/@�4KFJ'���B}{5���L8�^w������B7b4ݣPڒȔ[D��B�m���A#Ա%ţܜ�����3����L��`ͱ$ao��������6OA�d�D�x\j1,!k��Z�1������x}�W�Taz'���˨DhG�؋*����øI%L�����4�j)ʲy�]����z���@|���:k$u6������
��M�E�w��Zv�ݜJ��NlUF�.f����.*��C�/��
�=cGA���K׀�'�0y9K�;O�ea��b��{����w��0�u�g� ��w�i��B���Î�ª�3fS���1w�������o��{��h������]X�J�j�� �$��F�ے��R���F���L�G���/�\����
��>wÕ��]ezZ����3P�7P����.g�����ߥɪ�#*��M͆(NB+��&o-�,��?�D�t ��"�;��I��6;�68z-���cqff�>g"�q7��PWw�|�#��_J�:���c���h��~+q%��/wLidU�E[�����;Ĉѕ� ���0��J!�2ixf^<��Z��_�
� lF�Ag�#��H��p��B��������;�Rp͊!{MuQ�� 蓬���'�|b4(K�u�Ϻ=AԌ���\�>��%��X��D���yMI��H�2	G�&Kc+��^$�R&��r�'�ƚ3Jt�ʌ�@�(c�Ҹ����B��}2�D)r;� �_�Y�-[=@f?����zyЃ�K1���t�1B:���k8�t�4W].Uj�A�=	)M�D���2�K�Vc�O!�e�c��[����E��!&0_�O��.��ϰzn�f�dbu+Z[�J�F�3S��K�G��0�G�����1~w5ͤ���T��Y����0o����P��]Z\����/!���#�0bCR�O����sɖ�ə�ԅҠ� k3?"��Vd��+T�	�jE)巿��n�)Ppn��`z`X2�����_Vx/))D@�;�;��N2_��W���vБ66�݁��υC�@�H4 ��;���P%�Y�Y�Phߵ���^����W]y)�ҍ��<�M5Әo2b�������j�Sߐ���KI1���iϐ�����Ա��Bƿ"\$a�����ÁY��c��l�T�*1bi�1��'�,�Pm_��8eY��>r�@���lwE��N�i��3��K���gY����e���b`�@L���B�%$�ؔg�m��ɄXP`O	y�h�C`/m����ه�\���XO�1Y=Um�%z]����{�0t��K�uG}�;�Գ��<O��@�01���<�=#3Ƶ����S��S����\b�U]F(=�!''�m�`��W@W�/��b�i��$��(1
(Lp*ϫ�,:%
gw���tS��Q6ͫ]x N��C~i�m2M�N+�ja-��F��'�|�8�_y��*E��fO�W1~=�g\Q8�4�3#��T�g�kkj��=D���4����H'Ϸk���h�92s�gn��!nҤ�H.�aC��������,k��?��L;F�A�qy���̣�k��*���Q(�.�Gqj:Nĭzw�r]�P��c��ހ���ۛ#O�1�@[H�6��0=��:����"�W�K�V��~&�����2�#����qU�,�7єd��6�� �"\�DB��b�S�a9h1,	�� nZ~qS�#����,&�řk��Ձz	��8�+�`R5s�&H3���_ǒu�1p&�_TS'2��Ƙv�I�L$�81/3��.��1���כ���2�B��jqq�]�ĸڠ��
?�TL㹍���,�9Tqa�[�;��j~s^&��Q%����I�5���f�e�ħ0R��<#��=ٛ�2{�|kChj��|�����k������%�L�!v��cQJTtxFc�r�h�H�C�_����F����-�ƵԆ[�xr�9��&M�d��rx�� ��t�}��昱ӊҌ�ۅ����A���*�L�����םƌw���55���*�wA~�O�?&z��w������b�,�Ɋu���"�}$+`_vEH4T�!=$�H+��?���;����P��To��'w��{�ncƖJ{���:?�߫&RTTl�Z�/�Ũ]����Ӱ�n��qn˭�r�����w�������i�
��O��8�0���%��u��?�i􆑎.p��t3�p���(M�y��g�uGy��r
bEl��ݰ�a��X����זf5ud��m�
�_���$�2��i-~�+BYi�#��B������;�.��(P>l��dH��_��� ��5�
��\� �B�z�>��gaVg	��qtiރ���{���HrZ2�m��'(a��R�vs!ܲ.���L����(���¢P�����9rs��8����G��ᮾ�Z��~e�Ԋ���	������IEE��Y�i_���k�+{�������ku>��=�!��7�I*��q�[����ߋ���aw<��;:b� �[z�p]r��:3zKv������+��_�K]�M+/�b8�S �8���C��R�)��۽��[nP�(�[qM�!�Ӄ���*�R^�1�_c���SW'��6p���&��v��z��@�:X�:�^�Ġ��S�eo�R�\�k\��!'̥��]�����Ƀn���f� 4�!
*��"�)��xނ�p���U�uY��u.q��l���R����P�buaק�����鏙�Y�.a�F��_���	+��X�p�65��\�"�,4&�cǎw���7߃�`������@dZ.��\MM��AYL�L�Υ��^�/���W����U�m>�ٞȂ��νP��)x����ٽ�[a����[�1��� ~�U�9�ޤ��y��E-�+kO����8�4�0�d��p�(\F��{qߙ�;�x�����
��y�\��!L�c�P���֣�������1�=�܋fmƌ�.n��եxsS�B6��BY�3�.)eY�{��U���^��SI�����Y7{����ctWg8��l9荺@!�H!Pl�ʳ-K���VoQ?}Hd�� @KA=٭"��r�3���^x��Mq~��_�m��WWZQ�`�P[�Z;Z��m��S��)�����SO7�,&ȩ;�F}4~a��i�\�Z�Z}��𛾴.���	�!�腊���+~���]�I|��#�/$ x99��S���kw�W��b�L��ޤfU��A���/8��D�$>��D�c���M�M��k���f����� Τ]n�A��P��TSݯ/�%q���X�=�Pۉ�..(�z��X�2i�n���Ƭ��|�oZ���8�	d�%~َz�`��R��7,
���#�H�Ih� 5���O,�O�'n�q�Ѷ�bg.����d�Gzȍ?�v�R�Wh4I��Uk/�n����B�	nn{W�����T��:H�W��,��7��M�M���� �Ca�P�뷁�H�*+S�o�?����k�.�;K�݊��t�L��F�#n���<*������>mΤ���u6u��Ït�lhm(��l٫�����]S��:ܰ���h]�:{2H1�i���dgkq�񧊞D"��
�^+���g����q�La��zc��]	��"���}SG��5�0�}��n��5k�{�{!�hr%�ER�(��
���$?�x=է�ʢ�~��_�h$����F���<�#@�'�k|E�������Qz�y�Zq�Л�G,��V����.�u�h�� 7��Z:�z ��M�D�ѣ���	��@O�)�4���2�#u��
|m�_%2j9������z��e�`z�v�b�{ӧ�ճ�ǿa,�f!(;�?1�d-9��gY.a��+ �s�K��gYbeLB*�
�Y�|'+#�2ٯ�� ��)�7��_4�yy0��5f
������u5X�"Y����JK��\��x0��=�(I�^��۠�_��O�"�P�kūzr��ҵ��B�|�&w�G��΃�㶚��r�����޷�
|m�_�p8Q��PhK,�FzlN�?k�����l�(�r�7�~+e�B(�2.5Tn�`��=��:��I��4�U(�̬��` �Rvv��Ņyo��KA`֓�[�g=]�y���@��?$q� ���,�C��5���kS{�
��U�W������W%c��Pp&�,R�<��2ga�.�8���&LM)�t<���v-nhjx}��FOJ)˪���k�0Z��4K����W�͜�����͘��wn({+\�*��O����O�}R�y�����RH��1�3�K��}^��D칤(�@�P]�Ĩ·23�^&��uY���z/�ڻd�[�h,!�s1%���ō���܏�a$?3��eY�����@����xdzGhx]lv�ٱ��}S�W}��>�_z�������)F2`
�7�p_QQ�U�5��5Y���Y�jQ��6^��7�\����w���3���j�����%]��^~h�<7�~����nK�rj1��M����i��Y�Y�aa��DR�]�H)�J։!�
�?����bz4{�~���Ν�@ư���0��AI�� ��b5H�V�-�*�,a_Tx%?��Kz�9Z���Sx��Y�U�'�0�����6^�iwgb1i�y�@u(t��1��W�&x�Ʒ(��YY|����%���}���9���u=o���_��¬�d�rM�D;� zlܧ��.͍G�j��х������ �J���<�Y��J"D�;�8���3hyX*������)�YC9�ʶ�f����,sB��`+>�~s�m*�|��&IEe��7�oi����`�5���`�ey�ʏ`�i\�S�^�F+�R�5Z����an{G��X"������1��)�=E==6�y%g��l�z�n��'M���) ������I������O)�:�\�l���da,�(�9�N�mȨUa`
�\�	XJ?��e�q� �iH��k<Oͤ��_'��U�@Jaփ��# :�O ��c�)*�0=pD;Xl�W���æy��I��x��H��r���ǦWo�����D;5Xt2���r�z�*�S���j�p��1�xٴ鰣�Mc\a`8�"t&]#�Mq������r�lz�r03�]?�&_`�>�;���k�LtRf=//CU5f���g��k�?An� ��>�Q�4���^��+��?��裨�?�F(�<2�T��z��+:]Ja6�B�vC�����b]f�ؑ�>�D����lK9S��F�{G�ҿ�Mʢ��d�A�lqˋ��gᒥF�m����iS
��z���X�&<>BYv��yw#���M���U�G@�o�N��k��g&a]&�ɒ���iR
�9,4�F)�tw���A�MKە�eGZ����v����tY~��w�&�T���=�e�����9��ޏH)��ڸgmZ|��H_���	��x,~@0��Q�˥ޛ�oI|���1/�Q?s-�f�Z�Dz�R��s�����|�N�.7MH�&��ᴞ��:[C�7�'�3&���M�6�x6X5ʐ����s�E����P�'2��\x�SE������a>�_��P���C�Y�Fj"���<o�DG�jS�����/ t3��!���^��]�_����S
��vZ��y��z\ɣ�l-�#q���7n\�M�~�Y߼�貿V��R���vC�A��')���t�8]��̣]�69�`#���%�f#��X�`SSS�x�P�����Tܲ�߳��V ��H�@jR+�Z��
l��HF4-�	aw    IEND�B`�PK   �cW�{0n_C N /   images/7ec862db-5bbc-4dbd-b9e6-0d0e46cb58fd.png��S\M�-<�>���.������4�,�ww:8	'����� ��U����U�?M�>��}��{��N�ꪯp0�1  �k�7    ւО#rĘ���o^� �c�{  -൬����,t��?Ӯ�ܝ���G�_�RL+��1��%�R���������#�+��q��i(�yp~`�-�@�u�������|�2�A)���}�ǲ_����/�E� ��H�� 0�N�E/->#B���Bec��Կ �!���׾ݺ�A��#�Z�V��2��*�&�i�'0��|Ʌ�[W
5����yF���t��������R� +u,�FS�o�	�|~��F_؟gX�^���������r1��Ke%!��_�mq����������8����3���B�P�/�?�EY-�USM���8�����3J�v�'	�g�#%�N�ǀ��'��<
\ L:�l#�ZM*�`pb	f���fyek�P�h�WsQ���5���\
$ �e1���V�������%�.��U���VC�U�%��b "�;�l����b��TﲰU�y�������`�Qb#L�����D�
����!7`q�4͞�$We���/�:��ػX8tX1V�K*G�2x��ǅ���b��s�NU�D�N`4�F��6Ə4_���O���-�n��[#�HQX(/$���Ϥ���� <�����>�"a����$h�g~�o�ѷOAd�g6�����A��`�ـ���89=Ɛ���C����)��R������
�K�v�CK���
�C����{�ɚ��G-��e�on�0��:>*|��y�m��̶�,�����FLN@H��� Ж� �P��[9�׍D�d�6;�Ca���mԝ�F�?��8�a����|t���*>'������2G���}��-�~������>������m����lD �s��m�9�~��f�w�NG���p��BR�h	���r.W���������3��᨝���/�Q<��>h{�n��w��E^��.�_�N��b8�uU��*���J�F�2wZ��@Ó�g$܉�.��~ME�"?e��
WGI͡H�Pf��o�l����YT2F���An��OQ
�]�<'l@t��<��g�����+�O�s�o��"K@���/!{&��'딼;d(y	��F�E0�;]&���DI使y#�?o�&|@��#�3}�K7Gᤙ�l\n�M�FX��v�*� �o��%���o�hw��ߣx��Mt��a	�u�X����u��� n���1��L�u-��lލy�嬸"�1k@آJ=�B��O��]���d��[��=��ݶ�QL��<�{�����{��)eJ���v���4ߜ��x�a�Z#��G�ҝC� ]聹o�b�����0�U<�����"���Iꆭ�aNA` �ZU@�o����b�w6_��������|_9����M�_�TxN/2U�4�*�� ���t�+��|- �lT\��:��
ф����
MsI�>x��D�>�3u��� �Y��2��Z������4nF.b�L�̂m�q�z�����N"q��,�Ԑs�r�]�-�'A�)7����4�r;1��J9u��@����2���/0�PYk�̻������o������=܀Ґ`��)r� �	�oR���J�����̦����a�
 Rrr$;�^e_��-������AX��v��ہ�&��_��±u�@�$`�W@8wqD��P@w������z%�}a6z����Xh)�ݳ����J��ƣ���DV;�4�J��#\L<Di�L4�j��ϕ�Eϵ��zs��x7���oo3/9{?"�_�>�WԁZ^���m��H����9U���<1Fލ��b��)k (�0��}0�tm /���Pp��0��s�/׷���v5V_�@o�%Esl���b�a�c���s���S���x�Ѡ�}�&�׷�����B��YD�b�6qي�+��G�q}Q3G�*�Zv�	e��]�����:�Tl�²�~3��Y�?�n���6O��4��g?�f:���V�G!K/���۲���YD2��E���ef&�9�X�0l!���*a�3��Ǥq1�m��9� G��p�6-tJ����_9�y,~.��S�~0�Iws3e�I/>@������1��]�[��z�t��0�������{�����H�j��Qbp`b��`�$	�zN}�T
W*�3��3���򜴺��it���G��z$u*�٭Xj:C�z�����Ǖ�J��]FYb�/sh�PGKԯ���V3���_7f��ޝ�&2U�	��N����:x����pҜ����I��? ;�_9 +�o��� ����H��㗿���
i��d%@k�a�o�C�M]������)�'?US������������\�gQ�O\y�/��ayܯxY}��t��e��=ۅ���-��<A{�[J��L"*���2��L.E'��f��w;V%HW�J$�N ~�� [���<[|���>��X�:��������-~�j������M51�_/U�M)m��TW��E�PϾ���/���J%�0�����Uh�F	�ZX2#�p������kpjz,ԟ^E���x�Y�v��Jf5K9^��_�yVU�to}��ԝQj�������r|�N�?��{X}h�N����-�������h���D��0<Gq_A=���KVQѼy��$���:�R���Y�����&[�8?��R/�˿�����W�d�����ζdd����gs��f�1��������0i��o�f3�XM+�n�Ջ�b���r�X����4����k%����LVH�	j���6��Z�^�%�KQ����*��t��(p�v�`��� �dg�8M�������n>B��H���yufK��J���=�D��P��Ul�S�S�p0y��9l�YRͻբO�.���� ٶavjb�����PG�/w��N��7�LoF�\�.�giV�>����-�G��{��1��w���7�7R����8P�bQ0���"�����OF��<m,[�?�,��T���9�Y��Z�I�k��'q1s����2I�U{9�.�&�@��HI*��r��E��v߱�a-��Vi���	uB�����q�7grQ�p���wK���G�Ѕ� ��ҧ2��&�۷��b	�l?/:�Id�/(�IX��>'�~	�ি��C^��Ap� jx�V��=`%K�?Г.?-=.����(t��D��݉��??%�b�O�"=��.~�z�wt��N!x�z�݀e����k����#\�:���Q��C��Ǉ���H s�#W��О�c/��h��8�Ǔ��kǋ��T�zA��k¥��t*�,������~I�Z�\Z�P��D S�~�Q�
ہ%�t1�3/�Gk"��FBK�27�	u	P���_�����u�7h�Z��]SQs2�H?k�	�,=r�]�]�Z�9+ɻ�qɃ��).
KO|�Lz�3����Ć��^?���~j[����G�ҢEZ㻠J�;���$���Q�>a@x�>a_���U�AU]��S����M�^-9	�w�1�0�.|]a�j��W�;���8�l�@[u�"e�8ˊ�'�H7����.ེ�������0���P����!��q.2�|D���ϰ�T%�?�=S~�_��{�
Ƹ]K?�_1���k�;Ƒ��� 6H��-�J��~�\�Zb�ab5sñ`�x��bQ6�tq��N	��<��3X���I�9ɓ	^�=�w<:�{�0f/ͲG��l�"Q����
]<�׽��o��
��`���8��(�+h���k�����
��ʏ�S�1fz�����M��x?��Nl�[s�Ql�x���H�ܱ("}X�#�ʕYx�R�p;�j�9�OPDxFL�aA�$�����C�#�&�,C?t�[--^uޮ�<|��� �0�j�uJ�	~fv�TKr:�],�x�fн����9;�w_ؠC��^jDbZ'L�Lm�%e(�j�09
��{�s����TOT��>̕�(�ѲQs�p�����[�mܡ��F��l�ɿ}V��G
x����x�]��wќ��a݋"<�W�k�%� F�7G{����#�:�_�N�l�bA�҉E�Y�k��]�5:��;��8��~��R%t��q������c�]��z�A��;���qdP��'=}��^1�V�KYT�S�Q~�E=�O�+�.�*�B�.eܭ�I�d9�H.�I��5(���q�X��9q��A�A!)RسT͓������EY��>n�Q#�.��U�.m��p����z�����4VU9s;z�p����ܰ�6�Fn,LT�Z�(2g��%�,������N�]^A��]����wl�X���I�����M��`�8��.F��ڳ�f!ˋ������q�,yH�TL�4�r��V�>�YguY�'�^$Ѿ���,P��;�gɠ�5.��fC��˒��U�����o����6P�)�#t!��:�x�����X4'��X����Ov�+�X`Ň���X�?��\Ŗ]ܸ���_����k���g��ZU�x�������h���L�A9P���2��g�{Q��t��ʟ;4�ߧ2�!�j�y�I�IƏ�ΐ<f'v��/�0�7}U�ր%5I�킵��Qo]��X�Al#�.��tM��/$�4��`K���y��?��;,��6��豔�t��u�H;|���3,6��R31��߿��ܣ��_pB=�u���5�{�2�0����� 0I�l��h�o�Q(�b -*@�)$
tP�F��n�aG�E}[��A�:W{�k� RV�����G�]��ԙ��?ޔT���M�}7׀��6��@^�Y�E&��8]�����,!KFǘ�,�>O��#(�S6w0�L!�d)�'�0ft���`�z>����Mrr�U�ߠ���\�`�V�a��T���@���0�@�|I�<�
���>���9�c������՛II�{zI[ަ�9�Y� l�gND���RGc
"���IM	 ��`�2�����'0���� ( ��5�2*�ج������(Ҝ�1�J=9�3U%Oa�W���<D2�%_�6?�ki��W�S�h)ߐ�f���5�����}����UT,���)K$�\ �6��_ � �쉻iH &`�i"���V��j��\flI�(M��J���J�����/��:h�k�gd�L���?PA���;�B�_���ټ`L�D*� O&x�΋�uiּ�1w���Ugmk�S.��7
;"�B���u�=�,��ܘ��c�p��=�g|��ʒ4I0��b��D� u{  P�x�#F�;7��d` \7��?1L\Z%B>�w�>ۨT�+���栿UMG��\/�8,��	0㙦{q�"�y�H0[�U]��@�ʧ�+f�N>��-e-ʄ?�5!N<CMN.Y\MG4#sAY�@��y�'��^T�a�p����E��g���>h;b���#�*�i�lӹr�y����\����A�N�2ϊbC=b!K�.�̔�7�� ��\"ѲK��O���g��{|� �P�H�J`��j,Y��2r��٢Mv��Je6%��q��nPAs�J��m>in��(I��	�X͂A�dFS:�:j�e��"�,�p��P��Zx�KYfsN���q���K�_}�:�����P�i~#BZ�+��)�%;�RjQ�oG�^T���Ơ���N�kIu��K�yh�^�?�
��S���:��=D���E�*(��J�ë7�ru��%� pF/W&z�x��6v��Ln6d�!�Y(V���9ˈ�զXGf���f�E����\�]���w�W�,�qm��������O�����=Ff�vՋ�-|�5���'���C��T�AɠR�H��X��v�	Et 1�T��Q�v�n�I��e�h�w��\j'Q(�8�K�H�*�8D ��I馓I�P�¬��*�$�����/�r�ۮ�4�&`}��b`��P>Y����E��o�G~����X��&���#��� 6���#�>������.0�?G��(Lu_X����y�w��q��ͦ`4X\$UQ)+NN���pti��<�CT��)#�5��F	�,^	��ZO��EGx����;��DD��ݜ��y��Y�k	���(J��f���� ��Fbw����]:�Ъ9^�zuFmG����i�fDFP�,Q��ڄZ���y�7*V��&ǭ����I�\����K�q`=�!���Ư�,y"��ڰ�b��>wh�#<�����1��b }���v낥om�i>0�q�������0"	�#@�2H�f@ L�-pͬ�!��*,II�s ���ۦxޜ#�9�D����cOL��ďN���ϯ�
�M$�W��a=*>��1�zݭUv�!�� 8TʖE1�����RY��%n1@��0�a�1���@D�]v���T�Î���|�!Ҩ��ۊ�-���JJ����S�Ow�A�G�� r�����s������Ř*۟��1sc��_�k�x��S%dA��s-�L�4� ��W��2����ց-o|��xS~�?��m������D(�Q�qחb|2`W��� ~�7�B���2�	�%���LU�l�SE>��3�9b���R�������:�Xnp1�����R�<Z��6�I����.���jqzL�q�)�����-@��Oz�a��/Ĝ��&k�S��U�|`w�W&�@�0��%
9V����踴�5��-�4 �����(�D��1T��O��
�%&O>(�+VuC��7~ó�
ݪ��\3�¸��E2�e�G����I$�x��¾��@8���GD��,�$6d����^J
�����[y�"�~���@��.����㣙���'ㄷ�ev��I��r5�8�{����ͽ}�P�GQ�%Э�.���
V"��I#ee�h����<��UR�������H���I��!=m�f�ZS�G����������:,�����"�&�%�L�Z���1��u��ѫM<D%WVH�8"o�r�C2�W���#��	�݂�
�X����/	��(^�y�m�G�e�+��]�J��lhP�)͇:�dҩ��%v�`��F����������Q�U���"��A�q	��΁��$꣖�~���j����V�p�N�����O��T��[3@�4]b���}���hzF�zK����$�r�#�)�i#k��f�����(:\�O^Xs��WXL=1��	o�Im���Mi�	{�m+�, )���n�Ȧ�H7$=��R�\��g*N\G[�1j{[�LG�u6b� �ܨ%$�#������ �I�	��Q�0�<V`@�Zoo)����~~[���Y�`bFz �`!�w~Ni(�-��{��Wj�o0�i![��
�&~l
���v��인_鉧�i�H�خ+��}��t�xͨe��\@/W�c�a�E&=��$Y����N�LQML�1��Ij�W2�I �ҷ��a<���ή�"��Z1֍��|pH ��[�4�ΕIc[M����U|�W�3�'�1�O�i���E���V�6d�7J����e�����`�onL�a�3����T!D��X��)2����:�1��啍GF��hⴛ�C��� �"%���}7��n����9�<[<���;��d�-z܏���ө��.�yEW�"�i���o-?)H��o�ޟ�a��x_�8��"T�#�DWu��|�׃�~L��0/���K��w�"<&�^����X##��EB[�vw��v���#��>^�W��(�3hح���P�j��	.�Hfؔ��
_0�!)�t�RWDU�[
��ccx��G���w�ZJA�+U�n|�J�d��E�F����E���)	����X��x7�[h,]�&�A5u�M4��!f�����[%���ڋ 3�<�s#�ǔ.�i�A�R�g�������%�|� T�Q��i�]��m�s�~+a��|N3��a�Mu�D+��?;d�3T[��r.���*W3�j�P�E��Fl��Z%�+es֯%��s�=V��>Ǖp:����$k\��������%㉋�Ѳ(y�3q8�P~��{�31ӌ%������i6��Y��*n>6��D�#`҈�DM3��#�f�℆C�i��D�1�y�?ȤZ��ɔI?�V������ذ��� h�$q�s�Ѵ�_6o�z�	��G�e�}�x�,�9Pl��3@lؑV�,C<�#Z$�{)+�\�=&���=��߯��K>5�����D��~��w��$-���dEM4��u��>0�ݿ�
�_h�6ǿ�\�>�pu��I�$�5|�*g�uo������|�đ7��Uڬ��(�_�G��eh�ߘ�2��J���d�vOd��H��4Ӑ����+�~g�.����QQ�f�Ădu�M�ޤ������|]��m41�\��`e��aEq�o�A7�Mi��ᅈ�deC&H�����|����n\�\|9���?�QppY�p����9��ũ��v_q���b}5	f�Y.��Η|Y��_jy�r��jx�"�`�8ax�ǝ��
�>���*¹�H`N�hv2IG�%�@H��u�B\C����O5s�x6�����X��ri\~2t��i�0U2�p�����V��(��$��pQz��u9�`��qe�fJ0!�f��Ai���k�0
��0��;+h:S�,���p�}$�F��E��u�P��\��4�=:��e9%��H{���^�f4b�K5K��!���l��T�g�r�	�GA�e�ex=�r�uO+��;g� g;�@���C��C:������	jn�a�'���M���H�CH�);F���� 	1@���1=�����1��Ձ�Y��~ G��l��ё`G/�'����w�b=-o{J
<��p+�ʙ+�{��*�����&Z񪗶�>�Rd?-����eu|᎘5���~V����4�Lq�wsMĦ�1�4�A��:5��,��X�t�%R��)�3���iݔ��m1B�wb��Ћ���&&8�Oa�S�P3[L���j(+X}M^�Z1�\��-��'���{O.E��bD���.˓��@`8-��F�hnlE0k�IG�n��V ῶ���X1\9����d1򄐫���^ɭ��j�p�,����;�rw�I��2�wl��/dB~�����:�i�K�Sd��'�"w�V�kN����wM�zsj�[+�7%�B8���֌1��U�	�{��+�S�1��L#�d����H!kc:wD��3�I0={��D�NByn)�Qa!�Ӄ
���V]U���m��J��2N�h�2�y{��l���(X)���m�7�6�}6���/��B~���6�i�:�A��.�b��=1�H�eP)�o�#�\zs����{G�� ��y��/��Д�{Zl�3���?r�#�I�m������SPW�؇v���RA��)wr���>�x�q�{h�}�o���\c
�6'���1�+)�l7�ĺ}��r�ۻ̼�fR6��b�B�7����BLN%��#l(
�@ӑL 㩢����#X'��J��P��3�ZZ�S�~����Ch�r�d*�:��I��&�Н?�i�_�!�
��I���"�ߙ�����T�|��1�:�֬a���r"AgZ�&V,#a�z�����������7m2}{{��oN�>��)����LXi����� ��4�^l+����ƋCi�䆄����	��j?�Ej��	���7�ڳg���gn�y�]�b��
��R8>��j�$���)']n�[P�0�'�-���k�Y��i�{���M�RMH���guF�O2��	F�T�tVfo�J����`�Х��oy�����قJط�	oC/���֠�m�#���9��a$��/_�%~��Gk\�S �� B�]6�y�}�����{o����t+��A��"��8��\�(�m�g3O_�'O�k�(��7�i&_��������.k�:�3��6���:�[3�K+�8˚�D�����G����q���(����|��8vaq�U��yD�l� ;�g������Ą�`֐%ٹ!����[_s��b�������Y�%����T�ⰹE4��ᕝ����ی��v)����9��&��:�5T�#
x]�\ȡ��Do��5?pV# �QH7�o�����q2��(��'��~�B��7�����a���l�]���9��b��t
��1 yP�b���G+jj�YA�J���G��b0����-���s�h<����{��>b�*�0D2[�����}�C�궼y�U����b��8"�6�M-��C|i��AnTMɗ����:Wk�Ǯ�
^U�>��T��_h�ėN�NQ�m<�F��Z�pT�O?=��:����-�����!�ڏ�W7 �g�T5��ʶJ��o�qɯ�J�7À��qNƘ����/D���;�t�ށ����L�:����8D,v���%?��� i�T%-�2�~�F�� �g7'�<s�&K���S ti>U��u_d�-t���S��wU�m7l)�{��$�7%Eͤq;k�P־p"�ܱ�Ԃ�zZ�{?^������B6v���`�Zd��vd�P�pZm�Vᛊ1ѿ�4�ە�h��Q�nt�e�k��Q͠�[��D����0Wd r�-r<���j&�>td�ns�7�l�7�Dդ	G�ң����<�d6�X���z�F+����w#�;d�l���K�BZ�����U����4|��JMFƏY?��H�Q�]��0�#�B�G@��}��A���2&hڍ^]0'�b�KQ����Z��6˯=���d��=�P�Zn�M�YmK��P1��$eq����_�ht̟-G4�����<f��k��~�Y���%[��@H>��ˀ4��O9�.�<u��je��3"mx��&.{� �,�f��9�Xty��u���{ξ�&&w���L�Ogwvv�4���TϻORy?�>HIf�TrU�J ��l�ɹ��"������k-J��Rd/,�~�
�A`��Yh�:@�f]X�T��i�g)�sd�q��I!!�U�! <��=��"|�tu���~��g��b��Њ��R(
����n���ػ�藠�[v��X��3o��M엂��P���\� o��Ƴ�s��{O� s@�sv2�|J$a�S��q��yuEK"��m^|�h�����b�W��i��/g�O�;u�?U��מ[�&�����(y�?��`�Y�R�帲�s9��xq7j�ΡX���Y�-�oN�04�it��T�Ri���]��v�A��D�b�x�O���K��/���0�E�m�T��;�iwW�8~�"(q=����٬0����>;�:j{�S�\�@�Q9ݠ��|����9/�ee1��s���*G�H�a�2>#�$�pU�:B���G�OR��m`�t�+�x\�0�"�	�F#Н8��S��������On.��߿iZg ��^�Vȓ/J�S`�:�A��s�0�R!�(s	z��Ʈ�M��eC��wD� ������jp����Bc|��P�����������D���P��y%�G�g�%�z�5�ӗ���ʑ1s8����>+��m�������B�hP�{e��j[��Ӹ�D�K:o������\�=�^`N=���1��6�Ȝ�҅�O�:��y��k��~�;y�~X�����~�Vs(J�=]n��[�G7@������Ҥ�"拞 <�s{�v0�]sp��6��I�L����B�\H/	��!kf�NV��L��SJ��h�zF!�o�s+�Ja��u�`��Put�><\a.��A����"i�����.-���uc���ǳ�����S����Nh��6�?����;D,>� ~�U�q.�Ĥ� �à)����F�,�J@�bF�Ng�����_���Ë�ߔ���t��h����v��9���Rj.¹��	�zPGv�r)�;v/>�ҿ��+L�e ���3̓*���K����F�c$��F��o-6�B}�;�Z_�}��Rl��� p��D��n��v��`Kΰ�4�r��g-\��ռ���h����}k��J��jE�;�9l�h��=��l�[�h件�I�	���!���D�?bp)U��"J��v��yWs�)OLO����	�S�Ĉ�O*<
O��h�T����s��2;5�c�M�j� ��J<��ڱ�8����p΋5�qr?B�q΋��s35��}�e�t��+o��E�8��Y���q*�	A�o�0`ݻ�Z~7
�a�ņ�i�}��u%.O&b=6I����J�t!������-oy�����a�T�+�EDI�[�)5�sճ����1��w�BT���~8?���<�:�l���:L} l⻽���M��Y�[��r�C���q�$֡�[5���?���Ph=�'(c�|��J�r h���Q2�!2���ӡ� @�>�~*�[��c�6K���K_���[:MC��.�,V�c��×���	�2ãG�Dn`D橭ĂYZk��J��M:	�1 �Xf�	�3B�2T�x\��6y�;���p�K��3�tϚ�q�J@
�va;َo�b�ri���g$w�I
��� ���˸:DCf�4�oH0�J��ﮇֵ��)R�̉�u�7��(r�?��u>t��Qy��d4����V4���C�ׂ{f�}�̬�w������C��9<��=�5���g���5�~�	wC䞩����'K�
l���I-R�A�!k������KϘu�C�ٻ'���"�K\	����V���XA�"����<���*�O�9�����/%�5x�gw�&���n������_�r�'�.$BԹ&�5�߾;�����:<��z��i�]R}�!�(���
F��ݸ��n=��.0��1ܖ���7��F�[�,�EA�i��-(�*�
wx�R��7���K��km'��8ơ[g�о�ң!�ż��ҹO�1h��>+�&97D_��]:`��2nf���G�4�o�T�<�-�3��W��L7w�v�� C�#�ọ�b/�-#��\e��4��Y��ݓB��G.fɦG�F��p~�oSW�e_TcE	�-T��z�+�d��U�Ɂ׆9O+d6ʾt}����(��i��@`@���gM�X��0]����,X<3C�]����
Z*u5��L("Y%��§��4�)�1\�E s��y#��1�^)��/�͵c���{���&s).�����|2�E45���SB����S�`����)������*MdW�G�m����Y	u�I�fN�4�["}(yv�y��q����Vm~�c3�Ϩ�q���_����Z.�[{��ErR�ýj�I,���	dy��ަd�
I�W�C�6�,=��!����!�.*�~���2R ��E�����CH���u�׼i��%\`ߌ�����ܩ?cJ2Ʋ�ea�)|��oD*p���o9\U�-<V��m�ô֕�a���2�v��$��1�G9�f�B�P}e�"]��}���8�vX4"HX�Z���Jȃ�af����,�����6�V�8~�G�EP��arղ�WVyK,�il�dFW���=��?��'�n\���%�4>��i,3)"�S��}*�\�Tr�N2�<ָ��Υ���q��&
I���y}��/��Kf�uq
�|�c��@���z^����'���#�k�=�MK�f$�zi���M_��Z�ƴ����"�@ʦ��i��/�4�d�/�<���_dIkވv�T���pp�/��!N(��߭.�►{Α���3�۷;?�����`?	9~\�Yn��;�LM+#��P��g&�s4I�Z]/��t'�fwp"�:����v?!���W�h�W�_�
l���`�̽��W�㭆k^�J/��:��'H��������@.�>N<Ķ������g��k�����	��)�.,���x��?1M�9^��XU�#sD���G�/S��Ү�g��79%����w�i�@2+����.�j}M�;����&Q�4�z�j����2��Z�� 7���j��Gd$���@��q�<�ٜ�mqX�d'��IVY��� AF�q��r!��I\ݣ�K�v�C%]�q�O����Ƶ��O+9v��Ҁ�:��5
����8B����wYql?�p��;�,'��M7\r��2�[ ��#�&3k�<Lr09��������Jï��x���/�qeB~�͉��hT�SQ�wJ=�Z��rȢ(�bG}���Qmʦ�� Ea�	�2���2����G2�j������T��/����J��Cݏ��-�Y���{)/���ꝉ�fq��A�9Wb�v�����a���a.*`�m�'%��+t5��^�l.�/ޟ�&��F�`�8��t"#���}���������h��]\olS�(����P�?��?zt�j�� �Θ��Ln�y�t�����������b�:��(@Z�t��繓�GB��ᵳnu�ք>����X"Wdv:�6��w�I��s��H��F���&l�a1��Qy�V.���vm��<�����`�[>�z&#"%F~��GD@�=���F���EP����4K����<�*u)r7��-K����CB�F�,�]t�Z�RH1���:��w>\!Gt*)[���U�Ǳx���w!�v�?q�k8�(�ղ����|_zG�����dI��@�M�%�S1z�Ys�[s<�	����d8�n|mI�Dm��Ƒ"���`�Υ\A�����zK��#�̻��Zc�eD�@i�i5�􂰣�	���!C��N�E�b%�O'�5�b�k�$m"YK�]�+-l�S�5|n�����ij_?�&L�m>�-�h�
wT��,�L ���i �a�u-�x�c.`�^x_�$k ��7W���Ȱ����*n�[��P1N�}��9��Bc�$�N$^�o$XW�ݽ�ǵ�'�'+$Sn~*���,d<��X?���5, �;�`����]fW���^�KF��~�ttX��5�N�[|��i1~DI���/N4S�%������NC�g��L��߯	ר���к�ë3��6��~�j���q*_C�x��M�\qI��yy�]�4n�`A,yl��K钖O����T����  �0S#1-I����==����ޞr���;3R|���<>�3W�7�����j�1���ս�n�:�;K�̻!wU�65T.����f�lέI��w�'=������9ţ��'��!A�I�O[d2��T�4����m�xiv�V�$�D��Z-������ǧ.ѧ�4�����=N?�5Zz)X)�ji��9�L�T�j��{;�����mLr�טb��\����J�5�~n-�cn�
?����qO\T�|��y��������1��QL�٢7����#���
�>�,��\l��X��W^EmՁ��c3��"V�����MϿ�U�D�W�àkokz�
B�-{&z�3������>-�3�p�kP��Q�2��,��؞淵/�ZZL|�F�T���0���;�#d��d
ES�c��t�F��sv�I�l{�/?�ѪĘ�O0��-..��,��D��LB�N��复$9dj4�S@�풨ۯ�WO[MnM��q`���-S<��a��$�5�x.5w!l�����Ɍ�K���R�-q�Q�c�mDn�iP���l�n"(C�-��p6t?vܳ�����un��]/�GHT��_�� IẈ9�����hZ.��]�J)6PL��G���{5=��Z�C��A�;�e�EO1�S�dv�g�kB�w7J̨��|DɽKnc�6ǋ�j���/�±��l���]=���9.�nB:�
 �>o���N�!6�+�X��&lſ��=?xf�t;/��j)�!B��a}���ŧ׵�JgB�$N�T<�m͊M_���Xt)�����f\�a=���sЊU��QO��#������H�X�������WO�G;A{��(�_t}�
���A�/
�~���q�AV��z�"o[B�� �z��q	���~��kƊA��_�@RoFY}w��~4EUjq���w��D�<��m++|X^BJ�f�S�J��I�������5���������?�����O�����8P��K�i_��)��cn�V�����˳l�$q!1��8V�7�|�%��S�H��8I<�.>ũ��:���-7��ce�]ʈ�� ^@����w֮�t��!v��{�I+6��]c]3�zi&��4�'�*u���P��w\��#9?i�)ngۉ��S�z1i�d2`�X��2��"��*����G����U���x|*#MY���Z�u�̺o�]� B�5�E���綟y��������؊�g��9�L����	�,�[۝d>W0��L�n�m��X-�	M	��(&o\t�NH��!�0����_s�?v�֝M�3#U/�4���*[^�X�����( �Q�� ̈R�w4��M������1�Wu鲸rp�=�y��&���n|��&������|��9s߸��r�p�U��ج���:�OA3� �u�\��sƓ���4�,�� ZS�bH���#�P�.U�4V�Vue�L��7��9�|� j��@&����*غu�@�q���B�#�P\L�����]�Pq1�
̼B��\*��Y)��M��+u���A���(Q?�좊��� ����T*%?D�|�q�|.��Cpu�>P��RQ,�m��B��^{�z�cCk* Cb<ؼySy!�֖�w i���
/����o����ڌ��,?�<@m���hj��wGn޺}�o,�{A�㸶��\h��ٖ��o?q���&��2mʄ�C뒛�l�fƘ�:� 5)�k -A����9�����}�'�!\O�A� �����m��#����z�v����񮥾cV�`"��w}�uӘ1C_�����!V��~��կ���:��Gs-%�Pb+OZ�4�-$�J��E?���ڑ9�5q�F��n�P���C���
��q���������k�n�5Dn���,ńCY�Q� *+2rmjƊ�F]�S,C�k�R��+���]�����x�
ƏGaZ��B��_(�b�xH��&#�������R�B�R,R�ox=q��x�/E둴<���,ۖ"(�N�
�~��nF��8����=�j	��p
9سg�\/�V�38&��iz�}o�q��K'"��"�097�"���m7����`q�f�����_�|�k��Nڶ}�=��g�^�kvF ��'��F9��0�p}/׮q�[Y��6c��w�?��3��Z�1M��PST6���l��@�6P`���/�����Ӯ8��ͩ��5݆ ��H�e�0�j砊��X�O^i'Ɓ�7�(���|��~�H&�ǹ���������z��צ<��W�`OBձQ���,-����kL��󅛫��ȍ\�S��������-AEkD׊�����<n`��^ ��ڡ��gKk^��6?�
`]&��%	�r�L����檽�-�f���D�1P(��L��E��T&�!4K��n�3.!|}|<Z�T�yN�C.q��JIW��T³�P�8/�_4��k�ub�<n�(|K�����.�?عT��Ř���f)�b�Z��j�N~���0��~�mݳ䮻��	c�E{Z`�KϿrҒ%�glݶ{| 4@��ةt���@�r����B¶��u��\���*��x�I3���9Kf��,e���֓����f���@o�W�z�|���aC��;���'�[sg�`1̔
��A��Y-��� [BX6�O�O�]�XcB�Ê�f,���44���m{!��]ކY'��b�i���O���h?P���b5���8v���B$c�M���Q���ҙ�n-��f��z�������&�J�����C��P��d�4W.�-�?u���:���Ė�Q�H�\���
-)h1K$;�Y��e�ci�]W+H�ׇ5��B����|>'~G��q5�-lJ�
�q]�8�#H�7L�N��!CU}�(0�4��8ǽu�>�T�D�o�>���x^��=����<\7�P��
E@e:�s����7��Ү�[[�|��Y;w�9�uy��%R�����=�&a�}�h�.uu�:�ϵK�sUe&t
Y�q�Æ�=���?u�s+j��i�Y�j!�Qvz�Pv {2`!Dņ�p����ŵ۶����u[�a�t3���^��^}�AJ�=�
0(:v��n���?ũ.��w��D��������;�\v�q�&z�w�
V�G��r���+G�wi;�=}N׍�d9G�D�jz�4]��TTTHA$�H�۝�9䆎���\q��z=�nBQ��,������orh��dὢ�NY\T�&%H��󡚭�����J�����#�F-���k��������jk�ϑq/֕�\�G��5�|�
�;xneR�*���u ��T�U&-C���bI��R錴a�<Z�T`��e�HeL�j�q,��p� c]���*W����&:����9����ӹ���!���l?~䶵k�6���F��0*�|��Ftw
���uu�G\ջZ~ٖ	�[�B>+3hm��˺���'�0~᭷\�|mm����<����ͅ^��	���h�_�9#G{L�Ճ/}쉧_��e%&���xg`.`��2#E��)E���7��m.�Z��bm�{�e�аț����J�﹐ɤ�Ʀ�0�Jc�P^����Ջ�A�h�`�JEB����7t��j�	�����C*�!8k�pG$���:ot*G���-���*�C����7���ˌ(2إK�{�7vt��r�)= 3��q<-�
�B�

G���b�%�c�����A9J����*	5W*�K^�^T�*PX�.�((=r�����U�5P[[�D�̰�ρ��`��?�D��c$�P��q�(��*��(>J�g/\��~I%~�Zj�*)�u��09���"��T*��IBY�Z�/'E�������@�ܢRVJ�n�v@�����a(L�9�Ӵ��*�����S'Tϳ��e�X���?�����H����,z����oy���\�q�ى
��-�1:�6Hu��P�桥�D%�c�N?Sn�]�cx�8�0���*RI邐A� ��/�>GO�1K��G�v��c���B(<#R[[+E�
�U����Ew���T�z�:�����4ko��f����E�!��,3�إ�d2f(v��5�{!�VB���!���J�eЂ�c���4���M�3��8uJMW	K�;6�CZ��Àl���1<�_���1,�3C1��P�)�q		e��Ah��kvWm�q�	��SJ>����@�� "K\ �޽{�����ըZr��z��-�O�ʇ����x �|8�C�&�Q�,ޓ�, 6-�?�u��P  }�q�Y� ���f���g����.5����쑣�R {(fh�����5��e�v&�V��������]W�<=\�Mo��j�O�--����n��7o��!��&,E���ğ|��������J�e*xT��C:�'_�7	��!��y�l�ё��!�ǔ��M�Y@硅P�T%En��R��iZ�oI�X ��~9�B����o#e�)u��U#�U�&�q�kkm��7vyQaM� �s1d�5���klR�Ң˴�K]�C�>i��e�.�>���2�<���g��֩�V`]*�J-D���(b�
�ƎD�QQ"C��&Cn(,������Z�6t}�{Ǥַ�� ��Q�.�X�<���{ʳ��i.UB?x�^��c�]��]�[-������mA(<Al�0��{*Cyi:�]��25+
�)��ܝ�G� �_�&��p����یt��Ӹ�Y�_��7>󰙂׫ Z��Qz��!!�Ǔ�51r9�j�{W���?�)��NX2��D8x��BnL����B� �\%JEI� ���ﺊ-�9v����!��%��
^�4yM�≁l��7y�������'lU/��
!&]9����J`�����(��8���CX5�&[�+�� χ��ox��c����}2�c�PH�ZX�:Q�`숌ߊ���ԍJi*W�,e�^�>P�إE&2 -*h�y)7S��nˮ�x�����UҋEAQ4�[�d����h9�8��u��~��8,�6�b��n���pc�㝤�Oz�xG�k��/3�{)N�0��/^1��K!��!�>���]Z�&�?膥ֽ@1�²�H�r�Z�4n��_ �@�Y�7͠���n�������3˔CT(�&�B�dH@�	��w�?�'o��G*���1�����[����ڗ�Yw���?�jͦk-="`F�L���%����M`���@���تT�nU7������5(�a�����}d[Z�J�a������{�YV�Y���V��4 AQT@AQĀbg��q��}3�3�7���1����� �E	*Ar79t7�t���7��?�}Ͼ�Tuu�����^����{�����z׻ބ�T�dX4��ݳʤ�l�ȫ����O5X��׽�*�ɆP)�0TF4l<���ZX 2ɣh�t���B|&;I���� ੔�Ҟ��Pl�(
:�H�=b��g�B��	�z{�"�"c�߱������u�S�4%'׿��
)��~=������ڵk%$�g��[���O:K.m�a #�3"0�[�����>~ǁ�xZ(��$e�?�|�s�~Ԥ�Ѧ ��.h��1�+�g S�aB@5�+."�>�g��e��0����"O��=�6��$�Uw����������Ro�m��^W��-�&��4���E2�imih�h��Z�w��ϖ�$�Р25� D�4+bI]�~)��9�L/�r��+����8'��}�%4˶#+����m�F��)�%3�L<rFϬ6�["�n��t_��oHN�� fX6�_��=��j�@� �� s_:����B�7
1?��&:��~hs�[g��O��l&��ƍ��~�g�E3~�������iǃ�eQ�����-0y��>ސ;�x�U��ˮ~�?^v�Ņ�����,����J$;G�H� R3�lttt
��E��IBi�3:L$��0Ѿ�+�A�PHX$�4�f�y�4�
�4~l�Gڦ�n4#�!��f��!
�6	%)8�6ԙ dF��%�u�ӑ9�U/D�;c��
Tǁ�@Ϟ��E�D j�^OO��B1��M�� �q���rGE�ȫ�8P�L=��?�>i�}�8��A�l9`۱�ɞӂ��Aq�ϷPz������{��m���"ە�y�:�	�&��XY��?���?�z����nKwde����x#�̥��,��"�eX��N��
�#�J�c���5j "5|cj��͛P�i�%9LyѬ��)���']�u�e��N��"�WY5���.u�6�<�.���]��	�.̛6�`�8$>���w�m	q�֣C#<˞������֭['qU�� f�c>�k��Yg��[F�d���2c�c�\.&uѴ��4,��5^{�dB TY��+�f(��qKw����~Ձ��,�[��}��@h;7��W�,��Ͽ����ݶӪ���m�����&�y�(R�B6�!G�)C���F3{��������>ѽ�D���]F��1oL�~��#����5F�>�����x�A\L�M�Q7!ܑ֘ �6�&�d}14ֳic�{�u��T%�Su<��-�����-ظq���٧�i�g�\7�軔2�kƏ�s4�Q�� }�5eh�cb{l����=�;��EV��j��BK�?����?����}�9�,���A�g��x�	��ۂ;q|1���q���d�͗V�̑��w�|�v�G|Ux�`0!1��5R�G_a�"��w0��4���Kq��P��0r�C���D�7h��I���іZ���\`	'�I#d���NJ����&����kE+�l��3g��I2�5�l�$�rTg������]?�h��� 3&֯_�l]D_��d?$)KD&��ۚ���]�1$�\ђ&L�'@�Ǆ���?�{��R�n[� ��s�8
�7t�[��o���m9��Y�~����qg�xw�����K��;7~�w/�h����f
�D�<E�k�Z��b3�օ��d�����3VÍ��LE�2a�A(�}�?F�|�}Z}��"o
�2�x���@x�)91Rt���\'�rN�1ۮ!�N����2��=���`�E�@� H���?�A[��ћ�=��~2:12��V�D���ި���iܜ'�g�%J�y�`�F���2�q�x��]zJ�C'��d���;�-JEtw�1<����*���|�ʷ6�v˲H�5?�h4��$u�X�q�~㧟��#+.̶L���*Sc'�&��ˤ���fΜ%�	�6Zl<�����LD�lK,�K����w�\Ե�alR&��'�EF�?/z�Hm�)����|�i�iejt�L1Z�=io�������귲�p�D� >��0�>Fk�� �a�u��b޼�p3J�{�P��D�4�z $��ě����o��7�x]��}N D��a,uئ�L�ǀa#rK�3�"����1I[��ϡA�;?��@�b6�G�ĬMz~u-�(k�/}������:��|�b���gm��<IK��A�/_���_xi�y�U��,?������p�:��WM�x1�#eh���L��w7GV    IDAT�)	���Ɲ9�������V]�B��?�5��h��h������z�d�P�I�g[2㪫�[\�)��bL@�-��={Bh�FJ��_)̈́�k��2`h���"��1���7Z�F��8>����x2Ǝ�S�F �����H�`�@��:�^�tw69�&��j�OsOR�>��[qiݱK�������x��MO��钩��8ߢ����,��fS���+/[�z�9�U貝�������D���������s$<���8_�=�a>�N>u��;c�H������M:azH���X��5R�\ ���Zp۸�	������oR˩Z�Evƌ�ho�6�,x�Zwc ��9v�d3���M�mn=�iO[��`��6"h���14k �d�fr��$��vn��^�̀K�z�I���J0����;��o��Y��e�����[�	�&�WY_l���i��o�v���ø�n�B~���4�b&��:Z t�r�C|��iV�V|g8DK.h���af�qβ\�ҵҶք�9��i�$���Q�swM��UՋIS��YU���C�P���
}�g����y�)�
y�/�0خ��iߠaY�+ 3\���al޼Y.g4k�;������ ��JHcE��`�R��p�ڟ�Yt�=�i�8�5��n��m���	�^~}�m���������;kAN��d����LǱ8!��b�Y�Ko��Lm���ge֐=*P��?�\.Ձ3����=�>'C$���S�M�9�Bf�z̶��Hϛ�+�%?�����$�I͍�S�֘�=����hl��v�gi��+�C�F@m�I�cF�#�$YJ2Bf,�������ؕ;��c��T#¨���
Yq��Q���'���#��fYV���m���{�,6QO���@�7����߸�3k��+�Z:-'��	���K;r��З��v�C�����d�9`(����a*�+2,A��"Y2A��ٸH�	�bDݏ�d�m�M(È��
��"�n��hΜ9IQZ͸2%�� �~���D�hr�X@H�hzU�&Tj ��q�X���ܚ�f��X�W��&Tk���QxwOȺ��s�H������V �ݭ�dj��������eY=�^��=������������������Vn|��O'
���quU1DD��u]KBy����{�)�V�a��(V�U�`e��9��Ys�
���4���s7��5a��zN�J���M��G'�CBc�<S~�ր��76��hZ�h�ý<�0C�"�X$H����L��U�]ONh���f�� [BF'�aW��Lq5p��S_��������Ѳ��z��q{v4��$�O�>��_��Ǘ����/t�ι��	#��H�3vlo�I �4c!�͛«tJV�-�0�`���ZB�p���"���"[Ө6�Tpݵ�ޕN��:FG����g�93�؆Rt5)I1vH)�^{j�d��7hǀ��_�oƟ��5 �1G DA=�3�J��1^��퍭n�٪�P�`ݎf�F�� ����?���~p�Y��`Y���}��@h;������M����'/���������2fO�^�����ڪ���ڞ�@���i�%W2ƘB�EK��}�T��1om������	><וE�`�V�r�fP�C0d3�j�꡴킽i i�捭 ;
by�+�;}�$m�z�^|w�&�U�:h�����5��~���h�P#knW��� �th���rb����+����VH�0�}�ɘ���&&���J��Q��k����'?����<��&#4�A�g:��p�n���;�����_��;>YC~i��+i޲X�l���mfv�U��m�}$s���XL�\��QL����w��?C���q�Ɛ�=`����g�d��F��\-u�^��t�<z��L�%�X��e�)h�H�_fs�m������ӽi�m����o���ۙ'�ڵ�]eh�R���k��d�(�*�i���<L�x g���~Hv3��Ѭ�ĳN!���L6?�`���R�R�V�cWk�<��O_t�'.��ݲ4�����Z`W��}�!&��8n��s=g���/�l�f��^ޥ��`�d�I-���5��Y#�&��w�5&͞=[C;I��-v�c��@H���g$@�;W��������i�B������H�B�	���}����=�y��i�����)Ca�S?�a�	�R�o@��,&cW��a3�}�.��}=�'�荧�\F���@��j����_�`ťJkK�����W�r��;,���~h�u�[�	�&�(���Ŀ�����o���r�lx"�I%lO�2����n�Yb��Cq#!��P��#ϰ��orE�So�Q�z@hDu8K	>�N����������بN(��X�@�7����fLD��F�=�ȹ7�cBL�7f�2n�гax2���w��ϟ�������Z ���r�Ud3@��;<gV˯��k�_K��ڲ��D�B�S�{�
:�-�� �cZ������;��ř|�Q�:j�>��d�ˎּ�/��k
O!���P(E�Ɗ4��dV��nml���5�0BS�To}����m-Di@R��y���{V7_N�Zc̑{'(2"�)l�����>4Ƽylj��ٸq#�=E��m��f
��f���0Dg��F ���a� B�9;f�\\���Vp�����G�薿�_�bf�,+��{i�y*[�	�&���8�zp�ڳ����_Z��T ��]H�혽~/�.��^�g�$
s��0B"��A!���ٴ�X@����9��`�h[p%���dmؼj�����6�d�'��Q�z^jPG �{nTWat��l��i��!�ٌ�}�(��nHމ����V��p��*�����{��$�O ��M@Z�~։�1b)��J�j���"�j(��\ڸ���8���.{��r�����A�{B��+��|;��p�?��{t���g���#x��Ҳ	�ID���$�w���ݘF;ߔ
=,�lV����FH�����:��0�ש��EF����R�2�
!Nt�Z qi@���@X!��ZL��G�v���5[`�-0z�	������X���^��з�����)�Qz���`�c��_�XU+���dc��.����Qm�����kC�?��_��g�v�MM�}��KWн�S�8�}�=O��k����}|�l��}��а�LI	��H-Ѝ�KBc�d~��qBB����4��� b����~HI��I���k�@)F���P[�Y��J¡�:��M�N(�0��#�y�{v�YёwJ D�47���*ʹ�A$���6@j���ݴ^Ȍe���w��-���2��&@Jk�F��y�E�nI����t����}���t����ϯ�?۹߲�Ҟ݇ͻO4��xZo�e%�MX�����G[�����-bpĲ�$�)���4tC�2�@h����� Y�|�C��Qlu���2 �Ѷu�����I�yĴy"�N[Ȅ�����6����|E1l��2���[z��`k�l�q������7�x#5N]�Z�Zha?����K�>�-�.�ñE��R,�M�M#ؠ	BL��<K��(D���<�_u�)o���_z��2 �b|��Ҫ�iC��~���G�e�"��h�桓��[�&�N��k��W�[�?��w.�E�Sٝ�cS��s�UhG����*TԎ"M[}��=V&��4�h�7ޅ�[�l��JL&	CY��Q?3I��NPFS�64�M��xO��Y8�VU�iz^j��X@(%�3Az��P2u��H�M�����Ng}0��	�P��HS�Y����]f �IƟ�>k^���kɨ
|��+��:!�_�Ӧ׋�n�<[�},:!G�Y:��0�y��E�Õ���;2�tf�V�͊B�#�+��G�����������ZA!��B��U?�`�2��8����z�J&떳y`8 �[�af�7�Ѯ���;�	�&��G\)�cg���?���s����.,�G�����^ΪTCX�?�a;Rs�L�d&h���͑'�c�9���2e/����#��N��E��uK�d���'�^��d���M����#�5B����꟱ġI�&�he{�'Iŷխ�a7^��$8���LN�<,��B�U�R$J�Z�W$!�䴊c"�m����-`Z`�R��- 
�d��%��㿽��\^
 ���Hn�(��h��^�\�͑�z���1T���j�
r��֖lq�ܙ��9����+����:7�l�������7X(Ujg`��a�Zh��w����ۊ]�ms��޼x��6̞=�ͅs
�|���Pi���݋��|�{v�U�g��8n�-c�~���?���]�V6�o���Aj��g4���ӯ��2�hl�l0�&��$�N����D�Œ�o-�eo(u�o��Y�xٺ�Ζ m+@���~�h�x�jM�1�e��RK>Wg�\ە˲VW"����C�E+=1�7=;����M}_6�`�j�q��p�fΩB,�B��b鮮NtO�V�U���z�����#|H��a��v��,`�m?���T���A���ڒٜq���͛8��ږ��7k9n�Eh"a�-�j�FQ�A���_�<{��������n��Yo���'�pԫ�]X�X�l�����cf"��8�����;g_wn�q���o��r���bo��d�ص����6N���@=Uݨ���Ҹ
�Ӟ"�nI?�.��Ѓ$9,-�4�4���)��F_�]jgg�04�Ch�A5Rv-S-����"����D��n�&��i�*���e���>�l^�͔Li$��D|e̔B�����{���6@hWqH�m��	L�<�K�tww����L�8�.S'I�'��i�B�ZfȀ!���*�9��z}Rp5qÖ��R���L\)S��h���2��B����u,�(���;� ��:�[�����G���g�����;��d�&DM=��V�w���w�M��0m�@�˿w��^Z���[دZC.�o���HY!c�1�>�p㞌v�i���S�"�;���s%"2�}��^"��t����DK��r�$�S�5fjm�z;62	m
�XW��ݡ��q�Rq��g+#-��u���F_�]� F)�'ER�d E�0'qm�����>r� ����X�i �n���w��oz;�c��	��A��
����L��B����!�[��Z� b0+Z%Ƕ�9����x �*@�#ɂ�=����`�Xp�0�p��8��Њ����:�^:�c�8댷?�`��LXoY��m~���;������k�ql�{S�z̷������o�Tq��im���u $;e�U��r!��PF+��#�#�V1�ާ��[����
�Z�8�߆�2j=�������h���+TG�����t�����{��dYAP�ت2@B�r.��6ñB̘ގ��]��0�Za���p�*?\�n ȑݣ�[.i@���	����x
d�!C4��� �w�74�Y�F�j���7��^��ꆊ�&#T,�f�|7�
�g��w����drk���|6�J��>I��H���˺Z+��٥ M�51#N��8@�Wbǎ�8�������w�y��g�y��+7�C�6�v�Q�G����s4|V���ǑW����V<��m���C'�˥Z����D�P�x��Mf�6 �f~9u�X�Us���NH�-��13��2y���� J�����k�O$�f3QnO#d����g�9����.�,�h��3�~2/���.YjD:�V֮��/��G}A��v�b�ĺ2z��4Z!�F�eS	d's�4���[`�!�,�Ɉn�4�p�"��ZM�	g�⃙7߼���$�w�=����'Z@M~h��ՙ�	����;m>k�%�>�<�K�G�Ltc%-C�'ys&��P�[,�U��>3|�Z�#����8��cŽ�]{��������s�of��^��X�����4�o���u�Ǐ��h��q�]w?~�/n��i����`��`�XD|��H$@(Z1��#��@cK豋���1�h�^X˖������U�����5M>)���F��� ��
�tB4e����3�����&d������4u T1sZ���1��b���Z d\uz��]�s�L�oG�5�P��jd���P].��ki�Y�7��H*<��։�%��Qz�3 Z��K�N�F���f�HҴ�z-�խz������.	7��g]0%֟}l����1�G�w�����{ߜ7ݶ;2�mK@Ө0��Zs[{����[�ӏ(�5��Ce�J��l\�}B=��&�k)�ޭ���}���M��{G��1��L֤9jGZq�+�x�d�%z ���͛7I�>Cg��y��L�.�`��#S�[.�۶��f2�e�#�1M9�0�?!{���~�6�0k�15?�8b!�
��$�9
#��a����9����}�}'���eY�l��Lb����[�ûT���
f������N|z�����/tʹ�L�bײ]KR�c:G��Bz��LVv-�u�\�M��d!�����u�#��4Z� �p�G{{���+d��ҋt������f��~�R��@ �,
�B_De̟ӂ/~���%%r% ��
�A��+���ɲ[0\��yD�F����8�A��r����7��!^L�����U#�X��T�x�" �!
���Q�؇|�u��2�N�����VbZg��� pc8.�U�ժ�e8����R�c�/W_č)e���� ����d���i�$�� /��z�6^�N�2�����[ӑ%B�ѩQ�黎��c�Ԕ���#�F2l/��ހ�Qey�o��n���i��3�ݖܧ�o����/�~�?�k�,'D��Ɉ^�sT�f��ȯ³	`����^$̇����d�6�[�y��m�k:��zO)š����7H�ʄ���M�x��4�M���yb	�S8<�F͖eT�$�N�b���3�e\�R����g����~���O�U���`h����`��^�y�j�z��V`��?��z��^\}��M��[NvV6�o�0cۖ��IYV����D���/������B��B��hr/���E�P���."#�M�����ft*��>��1�ì,D�,F�F��lT¼99|���"/@ȧ21S���I��~��_`�l!v��Y�u��Q
���2�j_�:H�]�2o6�k�/$;��K@K^�`�e��9x����+�c�2F6ۂj5¦��Z��Wo�e�#�s��� ���g��WB�_�)� ���J�菎 ��hZ>�Dm2���&Ԓ �$�PO
HE6Pd�r5@�4��^HĳQ3N��_}��ʽ��i�s��3I����U�,.n�?��&�i�� e�h�l9� ��*8Ծ����	WrB�5�a��!�C	���^�?Ν	�!k�z����P�}�%,_�:���ps�Ģc��z�z[�pt8w��_�p�is�:����B��ǖ�יnz��10B۪����w��]x���eY�Z,�_w��
8�K7O�#-ǲ%��aΪU���ؓ����׮_?���33�L�m��n&�m�X��L�ճ\/ű#�l�Du�2l�Y�%wsq�zM���kutt�5)"�Ef���� ����s�[B\��5f�UC��_`�d!�[Y���e�p�Zd6���:Wg�T�@qDB�h���ru��4�2츄�~�\,=��N�3Q/ѢJXW�C���v[4Q���������Gf�1�z)��x�%�l ��v�\�@H���Q6�JeGR1����5J@����0�̓!���z�	0���e�F���Ʀ2Bj������
'�0}<wR��������6j+��ypiȪ.4`H۸����0
QH=����y�;�f+��)����R��q	��O����!d�:�nܒ6e�K:�$n�z���v�;d���{E8�Pۃ!2e���%l, Ľ��f%���F�r�p�V|It�K    IDAT�n9��'ݑ^�,�4X�3�-�w��	n����d� *���^�^�q��7�o��n��i�7ln,*ո�G��R%X<\�..�mqVN��u6"��֝]h����%��]]]�2z =�(F�,vS����uFhk@�aI.�1\���W���n�p��s	��.��	���B�h���!�G)�H�	��0B\\p����1�P_���X4?#��sIe����#���_���7߃��lk�r�(`9���(�Jj��z�c� 	#�7��	�5l�P���HC ����������J�I�~[�7$z�$$��!B<� �d$&�B�2��f�O�UB�50,�Gָ�
�ewA�L���ܿ��H~O0�0P����p�1|�@$`�[�]`s"LVp���^U,QA6Ȏ#d`���#�~WA��C�;�����w������K��t%�j]��l��Ɵu�L.�*�cb���1H����h�c��M :��	��j��U�2�˥ށ���S����������,ˢaS�3�-�Bظu�%���| W-��o 6�UO���[�x��ZN� %-L�P�U&A�do4	�z�\�3��C�Ӥ
5�N��Ic%�8R}ǞhGBc�B��Ƃ��˫��ݦ@�nAB	rH�&�6Bf����|{��g��LTF�r�H
̊tF� !'.ⓗ��C�t	S��!��� ��ƣ/���o��RV�PK�_Bd���tee��4�t�q�3Βzs��:1�z�(����t�g��:�ur|#l�<�,�#Bc�'!ǆ�1���Г�?�#�|�!4On?�K�'�K�H@��)5t�h��0�1����M�UC�jTݏ��u#�ָ~#4�Q܄ Y/�(��5D�"�^����ɰb�wEҷ	��)�b+�o~�v�]_B�x�UT��O?�-J/�i�;+߱7S��>dT�e�	1<����ޙ�M�w�b�$�>��˳�|�*Et��DC�=���Ǿ��K�?����k,�N]N�S컗n�}�o)����o����~���O*�vͭ���%:�d�?QV¬��2Sv�=D�K1S����f��_|N`j�%d�S�-@��?��y#4BR#����WBCe
�Z$d��rJ(mZAY(Z�7�����E?M�iȤ!�5�t�4���J>P�
�%�q	���8lI�pE\(u���B����kp�-��Vi�c���r��*cB�%�6󨆇���h|��D����4��	h��'�ta�xA@��� e�:�Қ	�%��]���K�$���7:-�-L4F�|�e���3|�1ݔ���5�k0K����(��V����J莀S��
�%	{z]-��|��E���zv���� ?t.>��S�������sP���y�d|�[wc��2|>C:s�>�Ƃ7���݄�vv���� T�ذa}1Hf(�;z��|o�����hm?l�w��F9�7Ϛ�z�_��~z���,���C6�FL�h6��� APX|�=��yݵ���o�r��i�^��^&[oZ�a���T_��w�>���m�;::�6F���:+�� G@��%�t D�����Bd���G	#D $)ʉ�����aCq."+�H�5� �͟�"63�	c�(,�����
b5���cV\��} ��!wbK����$�ǃϬ�u7ݏJ9Y��U�aDtͶ,M��E� !�H0<�@D2aD��@�T�{ec=i��ifZ��h�T��N�W@�aL=�hbU��Wt��sI�n��[�֐ЖIz&�m%@HLCC�+�`�<K��>%��T(O�j2�LXZ�%�������rJ����ՙ��|;��h�2N%,=|>r�)�R��$�e�c�)B����xs]Q��@��J	�HF�\ӀR#�7�]]C?��S���0��a#DsE j�<�	1���5��M���G��"IN`��J����1�ׯ �Fa�Կ����y��cٌN<���ps���@h��l�9�!�*��-w=��������G[vKgk�4{h�
��j-�������vqHh�h����:K�h�X��8Ho�Ŧ�w�[��ziհ�Ɔ�\��6�� �.o��Bؠ8��b(�:���$��ބߏ�iy�.~h�\<-G��YR2�| *�F��c	��+>S��{n���T��N+l� T���f=Tk:z���"�D�f6Q��i��CC\�4m[���C��՝�RA��/�Ŷ���@yjs$ȧl�,���1�4L���K�'��|��P���VM�p|&��\BƛIMA�������2�
�l/�^��2������K��IHL�Y�ա&�F}I�E1��<�Z��<P) ���c��������}�丰=�0���wn�o����}�7���d��}�0��5ƾ�(��^Λ�yQ2S� �6�b������n �w�؝�_�f�F>�I_�Q)�����8b��ł�����.��p'�S�t�q<��o������G�o�{k�����m�vr(WCds-����qZs��i�c����T�C1P��Y3gK�!S ���v��&� �� ��ϟ��E'�����E5v�Ҫ~��[Q�p����;�ڋY����ZY&��b��(��p�����1s��b?��
��ݎ��6twu�5Aq����>��T�c����bEʘ�?*e�Y�U!����Ѓ�D�B�����DD�x��U���_"�`!?a9|���}he ;#�Td�
��0D�XA��G-(����y���<�u����U�1á�
z{Q,�P�2� ��òX������Ԑ˺(���2LDW^eT�e�f�#�҉b); ��@\N����g�B{[;���ѳ��RC�Edsy]<=fk��\[���>AkF�~��kF P�4�����M����h-��<Ɇ���Go_?�(B�F��1�����"�-��*}ҒoC�ȚT� �0�i_QX�0"C˅:;ڥ��m9k`����� C�*,�}�CD�ag��|�����|�FP��G.Ƈ?�Gh��)��"�,��2p�n�o��������E���Z �ِ	�M���U<)�=[��&���_�zhՊ�ӳ����H]2��$���M��s|ڬu�s�	X�������ҪB���҅EM��7O�ȵK��o�m����G9�f���RML�N�Y�8����~�W]���+�k���8y���iA�\�]�X�$�$F���~��`k�3�7��3gI9������d�Mxc���y��6^\UN��j%t�<��̛3��\�ź��q�0�x�5���Ph�bp`2n��3;�`�,�p�1��ȡВ�WkH}$`��
֭߄G_�ͽ��(3<y��K0o�lxN�:�CZ��3�I����t��e�,=��bū�gf"
������ ��
}����ͷ
 j��sp-Ã�p���_;`�X�x!�̞���0I%q]fJe`h0@E������/㥗Wc���s*�S��8 �7-�7����%���n������x��`;��!�܄�f���O¡�̕葊���a��{��{�GF8��C�ߢh-�`[�����X��y�]�V�<��XgG3�wᤓ���wvx�dF�xn:C �z�M,_�2^}o��CG�l�t�*��\�˅|�<��Ǫ�Ba�Y��#���5�m�
ZĞ*�,��{�����\���6�!ݤ�EGu8f��Bk��:��3�p�!�${�
�+n� �K���/��+�C{�6���^]�:^~�u���Э�]ړ) $m�j���֡�(k�X��M)�A!��^���h�R;/��d�Gzᶒ�`#kN�Cl���7��a�4XGV��8��d��������ΓnN��Fx9�7��^�	��®e)�Jq�C���U�]��:�沅���	N(z��^y��i�)�h"�l�2v�)�u�8ﴴ�aڴ��N�͛2@�a���+��g�Fȶ�S�τ��spġ���0�g�j �q�3����dg��ނ\��?/����I�p���c�Z���CO�G��'����Z*Dh*N|�'&�� A�#�j۞8�R_��5����Y����}�>�,����/�%�80�y���֓����`��v�SC�%�1ˡHH'�$B��A`�a�����^�Pq�ݝ(U�hk��K_��9@P��c��5Xv�Cxu�:q�>��%8��C���ri��>�>T�t���=�ђSٍ �$������[���+�;�p�i�`���RS��6J�0�J��`��*׀_��o~�/����n��J�"��pӻg��Z%,\؁SN9��Y�O܌�X�N%`==u>_�1ĳϯĊ/a��UX�`.��0{�'�h�߃/% �8�ᵤj��q]�}K�1~两{���7j��۱~���یd@j�3љq�l����	-��X�~j��h�X�^�-1�h�g4+$&�u��x����2k�~�	���'bj`��Xո4����C��W_����ti-��1�B��M'��d��o�I��~�/���n/�1=�-��~ZnA�n[l�uª��u���_I	T�w���C�e@g�t	�4R��/6�����F?~FH�P%���J�"b�³���g.���Ub[��-��[{��{��ݿ�5��[qک'�')9�.�ʒ��K˩�@Ojm��l��^X)�.��S�T�hɑj'�QI�z3e�����p����� �A��=N�K)��'7���D�e��V�P�Ñ����z����EȺPO�E��N�_����R�-d&�%.�C�ѧ����o��|k^
���_|��F;H�4��f����ǟű�-���9	�:	�*#�e�f*~����q��hi)���W�5�(���F�����@@�	����:�g��-�k�� ��S;˸GF����]w?�ǟ|�KX8�T*������gc��;N��'-F{������m��R1�x��%`ձ	D��$���j��?<7ą����Bd�|p�Ed,�G��鰏�"b���61[Ր�'L�Wފ�^^�\~� ����@�����mLCE����! R�s�Q��M�ے��<^�%L�Xlю���[Fg�5�W�9��Bύ�f3�c_���x�)���jYv������	���P��9�߳�����G��cj�������%����y"0ld���S�����;(SkjڴYR\5] �0B�>��Jc�ؑ��U�nC�BƁ�;>�`_��Ǳh�'�-P4�B��W��O<�4���8�����%::הو#)����AX��4-�V���}�� �bX�RgC�K���QC=�B1;I��&�F���A  �m=�n��AR_�A.��C��{�>]�Z���ZcI�LV�&V�Ntb���ʢ��f�D�wۨ�9�cO�����
�J�k�_��� &��AY��g�R���V}|��"����d@!��❉�Sh���> ms��O��w��E]50p��q�M7��O�����[�@�aNal���\K���ed����� ?��m��K���h�l;D{���>�^,9 +�R������ر�^�����B��!�di���_xGu�G��a�ڣ�b4���qOX�l��K��l�Mjxe]���;Y�Np�
��'�b��}�bf��
����F�^�o‐�Kz�6��w�
�%���cR"�)��d��f�R��$m#�4G܄��e@�ͼ�h��`S�c�|xNEa����;�����G�
<giJe�Z`�+�n�P�4���G��?\�ɧ���A�0}^ُ-.l���"ȿg�4!+%�cƘ�Q�����}�:��1}:�Ҥϕ�7�3z�;��}k|�����c/�.᪟�&�1G�PY��'_�8��%��i��^F4\�<��8rz�)^��<#�%�_�"���$o��tS�#^*��ǹj��p�/hJN�Hd�a��-�$y]��e����G6,[KP� �'���ͷ܇M��(��p�����&l�_���p%�>Y(�<��d��ƬB�Ȑ����EC?�X�~�U���_�ul��_}E��Fd������9���G�̹���ȉF��AX��9z/�@5l�������o;Q�� (j���ko�Æ�c��m���,�n��@�w�hK$�^��b؎��H��F`�3=���P�0������ǽe��K�!��t�k"�IJ�ս�+� ���z��*��@����%4D@�',������%��[B @�M��!0��o*�R-B�f��n�˯n��u!��cfߑJd���D}8n	&{6m�"��lF�͖��<��x2�#�y���g�\��R�$�4;D�\���S����5�w��W��vT�����O��kW̟��oYVi�n{���ԍ�}�9'����q ��ş����8;vm��J�ɱ��9�r���PRs8��]MJ���������=3fΕ��$r���D��e��]fҾ�{���2<�(Yc
��J8<�0���p���Y\�d�SV�Ra�pO�� ��Z.��$;���{��5��$%% 4�D���da��5b�'��x5��\$����PA&�&B�n%n�����B��L̟�U8���V��nփC�F�����7(g��lCwwmu�\�i¾��3��̭s1\�pϯ��}���d���}�GP.������r�j5
+��B[Z(���y����Vޏw�u��l���k��ٚ�G{ f��5�R�2�j�C��MS�M-5I㮄�rdUj&X������6l�~>��c�w��VF[���
<+'�T�cdr�����
��J(�U�3mzf��4�X
�U��,�U���=W����:"2SJ0%u�n�%c/��~��B�8��A���w�`⇵�M�Պ�%��A�j�@cMu�����А��r�,���dsG@$�'PP?:<���b�%�-=�a_r�
C>�����Ϊ�G�سܕ;��'l14U|��}�CW���#o,X��흿��o�);~��o�l�8�;xx�{���+.��vJ9�34J�B*�1'�8�U�*�j�LY�/�{�i8�n��ӡ.�Ϙ9�\� db�{�X��6I� V3�2<e�+a�������
�U?��
���G���3�� K1wY}i,2>7#U�Q�c�Z�I(��|(���M�{4��s��FsWk�F d3�ƔJP��%7� q NN�]Y"����K�ɸbx$�~q�
<���(K�����:�uyh�,�\����y��><��
�Z�V�����l�����8��p�҅(�)�
q>�3e�p-�����nħ>�1t�3ӊ���?�4�����l�UJ�R�{�v�2DG��!B:�uףh-dqکKj�K����Fc��>C���v&�!��RhL���a�4�\K��V���n��n,^�������Zp|��<S���Y��~`Ŋ�|���ӇR�
/� 4�L���c�h�f���ɵ|X��EXs���͂�b�Ir�����˒vf�1		fQ)Ӿ@����y����_Ʋ�oA�F֐:+2lf�N��e&�"�a�|Ww�h������l��1:$o6B������Y���_`��79�bIͼ�'='ɸ�Zq�aq�I�v�W��:<<�,���5kG�19=��w���v[���_���x�͗f�]Kk��E�y�Om��P��72�(�b����Y IsA��:�O��|>�4]��g��V��`S�i)SӔEMB�bn'@��,M�����g�!YL�Me[x~e?~��NTj,{��<�v�/\���g`'����c�I?j\�%��Hy��x���v�:tOkǢ�sq�iG�5�z��ZML�r|q�f8�ƛ����c/�s=s�~X����� 7ٽGtK�m��\�o~�$�i(W��E�OZ���/�������%����B{��W��
��hA@�/��?����J���.T�U���Q+�A��z���c���2'�e��.����c�bƴnY�Ӣb    IDAT�dt1��W����P����0T�vŦ�
�o�f��^�Z��\�{�`a�:�x�4ܠ�����l:/'iyL�/���/����^#��=K��E�h��&�q������[��M\s��x׻߅��>Xܮ�Α�Ւ
�+�O�݅�^Y8
:����������������,�<}�l�@R���M�{�)��	�GX��<u�a2,�L\�-���|A����Ҟ����E�Y�6��\��0Ww�T] m6Xt���eD5Vdol	k�j �J��`K��cY�ұ�ɊŢ�C�ZE�hjШ��c_�#����Jq�D��$���ߕV����9C��?�����o���+�X�v�eY�)�6��KN��'�k��ǋ��������?D�C"�暭�Ҵ��,xZȱQٺKH�o��[imP:u�g�Y��b8G��IHL�L��S�lcށ�ߚl�h) :��R���R���d� �<��? �CfD��}��/����ߑ04�lREߓA���ga�*n��>��F/�*-WBe�0��ݘ7-G�2\�@�?��o�W�Ĳ����p	_��EX|@7K D��@��O��u7�~�G{ɒ0�8q���g���'w��C�n �d���Ͼԃ�o�_�Uh��x-(�h�Iz\ �JhoqλO��# �Q��"�1C&�ŗWb��N1F$``�ϰZ�UAA��i�_l��ؓO�'�cS�8aO�֍�!k������3O?F��r݌����OV�a��� <��
�{��*�e[���_�Kw�y��[��#�+0ִu����,Ϧ~��:��Bgg����Ƭ.�oi���w?��?�J�j�-�@�b�jy �]��C���@w�sj@4X¸UBZd�]}3�?�:�=v).�Щh��e\`��!��W�\~��xc� b��GD��ll�ڃ#�H�:��晾3ua�� �^rc�����-7[f����2�d�D#9�и��9��O���C7}��-K�Ȭ�����Hx�,��g�e��/x�O���+O˂_X��i�����M ���w9�������]����j�]/kK��T}*���}K�z <����(hLtc�Ŷ�'�ٳ��!k�5���~B������W�0�ֶ��E�w�'�[��~� 6l�m���Y��Ʉ���A�픣�?:m����|��I��X�q�������W?��d&B��&�`�]��F��g���{�ܼ��Q3C "�f������>��C�6�@�,�1\����xr�J��@-�/t��bX�!��l���8��Cp�Eo�"��u&b�z��1���B�E��K���.=��Q1w�w��!{vϽ�㉧V��S��&N��0�Ze |�T�~�!��d�,I�(���D�0N���q�m��ko��X���Q�?W`I{�K�pВ���犆���=I���I���իW����������04��Kkp͍`�@�lS�<Tjd3ҧLt���z�u����A�牗e�t�Q&)��v��p�/�1G��\r<�*Bx�Q��s���6���;�r�f8�,��"p�I��ۅ�x�� S�ҙ^i`�mi���26��/���Sҥ�,��C�q��n��+�~Ȕ���Eb�@H,24��@(���g.����w�	׵X֚���?��6��^���8�����ȍ7��1��8؇ck1�F�N�hEm.|jҥ�t�D������]�i.١�F�Ph�gj���T�x�ԫ��y=��6�Y	.|���_���7߅�}e�w�Bq������gY0XV�U�>}1����_�a�!"��$գ������Z���3;�<K&R	RM��!�A_�W�p7jA��Q��`eQP�­��]x�d!q��hCJ�SEkוq��C%ȠgQu!�t�H��E@��h]�>�����:��j�R�H2��ZB.�C���a�.1,��T��	 �����+00TD����C9&0�,@yD��;�D�~ځ	ۗ����W���#�t��x��פ-��v!�A��ޚ�kUQ�n���<o?m)\+�t���H�b*:s�Gܧ�}�T���y�c��}Ϣ�ɶ�V��Fdb�1�_�
츈3�v<�{�шj�3X��t����+V���Ò%�񑏞F�K��n���
�-\~�ݒJ6��)f��W�/3�̇����}���٪�e5�WY:`�6�&i6=�4��pf��uRў���j�m��86'r��>_8:�S�F�_ڼ�ܳO���?���f��-5�j~����㼵��c� 5B������^ui{׼��5j�d_�ex��j�4q�F(�%��00,O�^�C̜9[ҿM�j��mQO�zaC%�~x��)��wcp�"~5L��X���_EG[Ae3.8�L�v���P<K��/�w�6��-æM��ҧ/ ��T��[(�ĞXу�n���?bٍH�*���uȹ>.8�L�l��P_��OV$���z�M\{����UfA�L�X����MA��j>����Ӑ�ג�u'�?1��Yg��m�Y���[�WU˃|h��	?�	��C��&��
��7KL�>����q���Q�4BT���2��_�=��|�L�e.���@KU�B6B��	'�p.������OۊN"D��0t�*�����W,�+���yI�7EN��s��dS�DcNsgw�?w���$���R��e=)�z��7b��y����D��>�J�?��b9 .���~�O�A+��
�����R=`�3�@(}�-AI���7l*�V�G�@���a�Q#7�R�!Ɋ%x�PS��!c����xq\+mZ{��^��_��U˛~B�'4���i�I;K��=�����?��3�����.d#qJKܣ�!��-1����0�㙌Hz�_G	���, &�;�
5��Fh�y��P��>j�X��~|%���>8�(�h�����!��h.�v��֏��]��?y},��s�/(�r��o�q#zz6�`�8F�P����-O,�Ų��F-�"�3"���R 4���_��g;2eB���L6�J`�;~�~�8B��9X�+zMQ���l^��Q�{�Xvr����iK�84�1�5E��"C�4��g���g�܉�~�#���ޭU੫"mR-Q,��q�y���SK���T=��Q�7���(ŨE.\���ְ�<�E�8��l,�Ї� ��ȱ"ք���� !q����]�[ߏP,�q�U����U	o��l�����Ł�����Zu���hkQ�%�)��!C�1��ͫ1�\|�ӥ��U%�M2m0�����V��_eS��WS�T�V
��>9KH�'i6h�i��Qd��FdtNl�֋fH���}y�$s�&w�Ġa�FH�f�c��9O��?��m:���?����+��=aM��M�]�!�yrF�BKN�3�q�Y������Y�F�9V��+��~�rf��.6~�6�0��'l/kl�H��7'a������7���x���Ij����d�ƌX� !�1F#�ɏN�O=�7��z�Yڢ^6�����.�df��aG�8������BX�"/Ԁ%!fē�c��߽6���K���S��캻������_`�v�>� k��_�ӻ�WB�d�,D5񺡚���/��5�$�:j���f�'���\�Y�(W��z1�;���n�'�r�Ч3rV��,VP3IF���N��|~��gq�ͿB�k!��iA���m����|���? @譧,���u%������oW��;V&����pĴ/�̥������t̝U����vKX'q����C�,k��'����UX�S�P��s�xI8�i���D�X�eG�O���G�|�B��ۈ�^.�O(�m|�?���E�����f�D�� |�;w�W{�mi��|��Y�c2����|&���Q�&m�fx�99��h�����rX�-1e� ���[BF#DA<��p������᯿����[����`g&��w�h�&��������~�Ƌ��3)��!e�*6y!&/�Ak�Lq����oq�th��ݸF3C��k:;�d75�j��Yc���B#O=�?��>T�V�mS�3kEe�;���%Kү�jN=�`�w�1h�ŰD��rz.��|�����7��s�8Dh�e=�$[�̞~~?��n��u�d�i�
˘=-��_v>�Z��F�'�E����=�����G��IRƴ��m�~(H�K�ޑZZ�UxW��c-�aRdZ��1"$�Rb6��	��g0D�l����f[E3EmM�󐁇��|��p��%���Alg����ml������ڞa�h��+�-	$� ���3�x�,�3��N;��:r�f��(L�i���2'�f�Q��~JK�՛R�F���XFqT�����ߣ�e9�
˨�t-d6����Ƶ�5k.��h!.M"�b��C��������ܼ g�F�3�1/�B&���M�2�44B[]��������1�Bt1�c��͛1<LV����F�w?��A���(F(����"Hfx,(�EqhNw���/oἎ�X�!7?�n��ݳ㾡�	��qw=�R�;��~�@%{��m/��uN���'���>U���BZ����@�Ϸb��R��xq�JRQ%e�L#��/}t̬1��\�_�ˮ��a"� �.�C}JM=o�,�YW6�q�p�~��OB�^2	�	D%�Bk֬��?���X��� !��"�������މ ̉@���i���8d�,|�w�5K���I��,ʐO��)aXL2mFU��R��r�I!�Pu.��m�e��ԈH��E�$�]½�=���~��xy���s;���0�|���Q\��"N?�zyK�R��n�TW��<�,z�k����o }�r�~���a�~�aEp���j��G{A,�~6��U�p�m΅�h�D�RI}1�Fּ�
��̭ٲ$F����	�b�T*����`�<��������k��3������|�X�zb7���yR��+�͒N��z㿵 ���a�]����Alܸ!)L��5��Y�Q̹��K��} DF�a��ܘ���||���������,Km4��n�{�(��7�"�co�&�ȟ,���=���J��\�ũV�z��B[���d��LW2�&�2N��޲���֛HR|3�1c&
��춤���� ݯS����S��+^ǲ��J�&�c)���9`����k6`�:��O��AȰ��k2��Cxˑ���-n^���Ud
����1�=#VbES���C	���AӒuIe!Q�tZ�CpS.Ehi!�:Zd���E���G�����^ �gk��=�5ɝM5�1��?�^p
N;e�x@�o1��'�Gx����ب�.�~ u��o� �Z��31g�48qE2�ZN:a)Zr�B�?{�f�Y^��N���4����r� �s!j�C0���{�?����or/�.	�`Sl�\p�2�d�V�]�)���?�}�wΙ�Q�s��<s�>{�|�[�z�2`���ضI��\��k���w��/����;d���+�g��w0��ٸ���"�.�sur
$��{��������R�� ��(3L�9���:��j�xM���`Ϟ=	D�l<2{��q���I��с����iG�����?~���@hRc~�M�Y�$�KqS#q��ª]��?>��w�� D��o&����:�G��ԩ���櫹�S��I���p,���<�-1��,��4���>O���!5R{j��	��#@��6Y�T#4�+/���o�i뱤t"@���Ʒ�hN�F��#�N�\q�B��׀�zqLj��^�(����r�cN�I�K鼬y�M�kʈDu&�T�h���A��V�g��e���of�Nǜ�xp� ���@5�V�ߛz��1Rn$�,�n����w�|.�p�|	�(z	(��FF��~��uG�Ed��>N�^��Lٴ�z���l&�5/���ȇBq������\ /sW�\Ɵ5�̒{R�<�e���E��	4U�c�~����J����RJ�7�]�� s��G�-d�2�:�C@+�����w�y·	2��)f�w[��w�q6a�O4��+�41B|�����h��R�;��ӟ��/��rjk����ݓ�Oη��2�����q�g>���=�z�Q�.B����I���h��՞!�O�#�>B�4�f�R������GB+Wm T��� L۪�!M �HQ�@h�.@����k���K*+m����1���g����?���^���P�3A�h�A����.8�8�hΗ�%�t~��h���H��O�[:��[7�Ų����M�E���aW�8 t���"v�I��.���1r��ӏY�;�7�����%bmBĳ���6�%�<�x���eƌ�pO��P��i�Rn�뮻�ܑJcdD�?Y���������L��beuj5�"��<��R�H&N6H!5T
ؼel%V�j���b��ۮDZΙ.z�E�?���:��/܇M[FH��3�K�g�X7�����X��1n�I��!��A�R=��4S�yM���8�@H�P�F-��8!�Nmhv_�����/v�X�)?���@����
�B�v���ۿ��[(�F�n�;N��z088�L.�@��	����0���N8Ȅrg{wooo�j����32<G�ҩP�cv�-����� Df��e%�3t��-x��ԇp�%q�M� #���xҥ�����mwP#�Gde�U�׋2B��7������u�,%B�%���a<����,j�7�F�W��I�C�l�7��PZ이+ר�P�K��.^?t3�gtkH�t�Q>�s�/�#�DShfV:�A��T�U(`��%�]v� ���h�hreH���_Ų��_�R�o�VJYY���jZ��������bd��:#���A��������
^\�C#e�>���a�AlݶS�Km�n�XQ�
��G?��P�Ud�qP�%-Ǎ7^�B&	�%ps#r�t����݋Mۆ�Ҙ����T.l''��$bL��6��� T�����Yp
�t|'v��^ $�u�2Bls������?�����	�ϛ>��>��o8��i���8���Կ��m����?��z͹&��3�U���iV�T�-q��MzbY�l���4)��v�F��E�&�G�od⛚����z��Ȕ8��9� �8�$@T��"�|��`��PQtB@�w܃z@�k��tP��^���`Z'��/�;���:&O�,w���x���Hez�G,���~�bƙ��I�Dp鴇t�j��i����� B�RAg��?��;��h�ɜ�)-��j2������.�NZE�pZj�":
�,\����R�[q�4,_2]�E�/�D,=:�Tپ�c�wQ֨?�0���F��u�]�|�_{x D���Ŏ1������_<�d��v���[��a��-r�	�LF��ƒ�8�u�%@�S��Y�q$A5��.Y���~�Ԕ���^��N�[E����ߋ��F�<WI�njަGޫ�ێ�&
"�q^t�޽gg�� � �	�~z�� b�_\HT�6���k/�����֯���\�P��\�m tr��m%�c�
��u�}��w�vp�z�܀��3uZs�(���tzc��@h���|Xhٵ��ى��.iO�V{mQ���)��ݎ����aN�@�8�%A�CŸ��~�ː�!�0BᤁЯ�ۇ۾���"��YR�g�����3��f��]
zTc����p��������J@E�N�!���B.��3f���[آz��t6-�'� �Z�rV&�u��L|�r��$=�<_,ݑ?��kA dy���O�J撍L�-�3Ћ�sfÃ��6���{�b�l�]�Ҳ��k��0�*{�YT*�֩/A�u�$QI���Y�����)��GB"d��@��j5O�ƁQF�8p=�`*a�P���E��$��T	�SWl
�s�t���i�W�V�;���y�W��n1    IDATG�O��v�`��)��?����e�B��C��޺�����>	MAr�,��.J�Q�ٻK�P$� $[��u��>}bi���EQ5
k�ko������7^s{&cm���ֳm�&9�m����_v�U�����|���^�ȣO^���[��n�c���вU3?(y����T�ؑTw^"-
�9�M�>]�!�B�(o��z�+�0f�8y�F����>��7%i�l	gϳ�5Q��L��W%}>�(��` '�~�̟͜u��pF��)����%b�VN��&��>ť�t(���6�+/Y��o�R�������eK����}l߶|�MX�l�(CX�qI��X�9������mߺ�0��by��h:)aG������) @��&` �-������۾��� �[��fe�%K��y�>}f͘�\6���hQ������:��P��W^���6Ջ^)i>7�K��}p�ᇖ0"dF��*�9g&-���g!�R���s��h���#��VKr4;���h1�/��U⻴�h�(�u$d�؄@Pg��f\\w�r��
���lv/�UF�������a�ֽ(��r2p��ek^؈�R]�Ů )U�S:;r���@Ow�ٴx& �̅�=�Q3gt���{�&�.@��:�&4Fc��JFh��NA��lܢ
s����{,�:��L���@uz���"d���D@/ �t!���Q�krH< ��i�<�I���?��[����/��eY{��s�lۯ�s=�m#7���e2 ]�G���>u�<~Ŧu[W�ӹ�;=7�
��ͳcˉ��
�Ч�3��c�^�Rud�u;�^��~���kl���
9a�~ �i��l6���D;A�95V��	@݋eJKv�+};����9�:���9p��I�"z���5����?�$����q %|�#������R�R�B�L�x+Wm��}5Bi�Rx�cMc7>�M�J�~��+Iʜ�a�C-?U�3K�.l߾x�-X�Db�E��IS]�U��u_����o�dP�d�ݙ��3� �����W/Q�)��~��{-T���w?�G�<���C�Љ��3��C�В�LjΓ#9N��q��<,24� �0��ظ�Z:(s�i(��;/3�g�ŏ~�(��4���YT+E�;����ٍZe;Ģ*�[1����F�@�Ԩ"�� �G{eR\�aI�>���	�^���s���\�s<~S~bg\ �ɜA/�gYy��x�g঻8�)֐�vb���g�Ax�,*�*��:1{�t���E��L]%���)���juر�s����3��*H�%��m͓#��{O�'� �:Qc�H��e�uQ���QF�E�dX@]>	����٤3�xl�#��*�I�b<"��}�*2B���SE�s��d5���c9Y�f�,M�f�*�LL(p�p=���*]����>���W��gY�ș�η��3�����H�: ]��,z����{��X���Мb��[���������lGW9��a�͘�7xp������Z�ՠEN�� ����/���vRR��N1�ax!c7X*�����[/��1M��$/��]4(	K�/�+�`N>��7"�8-B*3' X@���T��b͆
�z��#�@(��+=�FbǕ$�	�zz�V��*�s��+Ҕ����,3�Y�<I� �x8�ju�K�~۷���?�,\���p�_C��X�>Q���
��;�����"��vk�W+Ⱥ4`,b��Yx߻^+�Cm�S��m�`���߅��~�1g`f��A�Ё�]V���R͓�p��IG;��9��^��K�m��as�w 9O�<�"��V,7'�F��(�gNò%�$�ª�9��EX�p�̆�D��d9(��G�j$� �c��U�V�yޅ!P ��1@H���&�pQ�בNe��ws)��j�����;�5;���f����w��0�9��EoO7z:�"�f���x��ߧІKnV��-�g��s(�.݇ԙ�(�Z<��f���u+'bs�HW�%a�D�h���z
>l�.�F���g�훚����2$�D,�5��L��}׉��ף2AM+ c��q6@-N�����?���現���c�m�xbC?�=I�jof��@�2e��f�{q_����R�Z80Rv{���lGw��pe����;w�]288X�m�a�϶m����Q�M˲��
8��.6�!:::���'?��@Hy��$�xY���]��bI�@�@$߶�f}_��Bq�-�H�Ee��1�6�
��*�"�J^%²g�&�sb3���n�
veqZ��V��D
5�����m{���ߊ.��(�K�=��+����$W���w��~1&������BG.��/���1�Gc
�[f,!q�U��Oo�ڵ[��v!��J�������-�4i�8�|!�i�f�C�\���~\u�E(�I]�PV��=�R�v}|3��	����7g�s�p�D�#p�BTÊ��d�a����2��ow"J���e��\I��@(
�ϻ�����]�v d��U$|ڷ� f�͐�d�����:.<�#�^X�;w��]|K T���={f͚%,E�� �y<4_�Et��ۃ|� e�b�,!��f����%�&_X2/���������<��W���b�K��|���A&׉z�"'��2q�p0g\�a�x�	R n�宒��(�b�(Yc��a�����B�zS%��uʅS-���k����O~䭷��,��ۯ�1mF�d���FR2cR���!]�1s�����׾��]�+W�u��:#�4a<��j-�G�Q2�3�ֶ̓�T3�!n��1��(����q��ڙ��u�R5���trT Ėq+*c`f'>��75!�: D�HJKc�}|�vB" G^\�~���
F_�A�٥���Ҙj�<��R~P��XT+�
��i��>sA1�j��S���_q^����0�R�rhRZ"���ǟx;v���p	�B��[��f��>���~�7��k^}q"}a�5@����C� �IKIn�΃*ahhC���R�7�E�ʒ������y9gn?r�zz:�<b��q�E+�e����G����ck^��O������#[�aC�ϛ#�#��}�X�|!�,���/\ $���(����[��D,+m�� �#�wp�U�wQäm�I�{la��͘�?�B!'�K�
�%k\ ��0����]��}��+X�~#b����^b&=�R�-����,fΘ���i`:	C�_|q/6lܢ��B׼�B�S�R�2����YT�1R)��ظu;^X�^�o��s0w�"����=������-���.*j�,N���?K�i���PY�O�2@�������y��䬙Ȣ��ZdNZ�KFX4�\:��պ���������^{����w
O;gݮ���Yw�&��;�j����M��ӭ����ev̴��R���͊Hu�~4)\��D-~E�����.�9�)搌����~R�� d4��!hP 4���V D�M���T!��I�<�������ڄj�,��Zɮ1�EDB,%��<���Æ@��K��m�5�<'9���~ƕ��/��}l۶�柃�~�5Z��/� �	Jr�{�Q���M�����gϭ>�ۿ�-�M���o�s���ԑմI����i�G�i:K��Р���VZ+�l�ɶp8�Cq�(��իpފeH�l	���� N��#m��"�Y�	{�lݱW��0͟w� �X�Hj~�BӵٍI���y�Pj����y���2BrF}�	��(}��.@!��"Ӗt�	��~Zxn��� �t:��HJ�c�NF.b�R9ā�!�H��.Hl:�ّG&�!�q���LA@`��2�~�Ya�x/�`9�t$�I��Y"��EFȒ�4�=���Ȥ�A�]��{�i�n���K���*K��-+��ԙ|��n|���5O#��8�����P�c�M?��p|�t�)j����Z>xp���޿��?���4�˲��a�~m��L_ſ6}���PX�f�����?n�]�J���z�^���z�+ͭ>���#��QpX(ƀ �:������D'b����1�\�P� �fiL���8���b͆*��MB�j1�}���-X0;�~��4�\�ƞ݉��| �(��8��c�vX֨J~VT�Fh	���i���L
�TB t�?���{��Y�?�V̘���ez@�NF���A9�@Zƣ0�m���?�r7���e_�[�7��:r�_+#�6YHΝ㉮��e>��S�Л�I�i/�!_�����3�p��+���~qI<{̮+:��7��"t��w�6lX�ёa��|���Jy�4)KI�-^ԗp~�{���<ne�{l�����+���	�&rp��.��}-��g����{����00���./��nK�>��	6�/���m�I&�dqbNI�( (�'��6|�����r���2���y.˕�ټ^�*a�r��y����n�T"� s,2�rBg��mȋ[Fΰ���j��~R����� �����K�c<��M4S<�Ϫ	�֘�ym�p�0(����o�⎏������u���=m tr�s�nm(�{vo}����/޼y�:z��j~l�[ߕ	"�1����=8�q����!�B������rgO�����0���K��Ur����k�b��A��9���e��(`͆�&�17B���fu�e�M�9$B:�<��n�~�OIiL!�x���Y��ʸ����}^��|�p��,T���CB���W��*���K��y�\8˲ΦJg߯KB�@N�4M��%�	��߻�2�Uc�����k�\ �s�ِI��
蒛e8���H�~����Lb"���%�J"D�ެ\���S+q�e�Jg�L��.D`#d|��]�k�n���:عs'�mۆ���X0�@��4u��s	���Ɯ\'}C	#��
� � Iט0)bi�c�"�Ii�BtЎ�:P�Q懓����a�&���9�9�[�X&a^/���D��N��s��,��f�;SYDv��EP#����ĳ��OJ�6::
���e���H�m���7![Hi����z�^;������߾����~��`P a��Z@����^�2�@�9�1�V�8xp?j�jb\ʲf"�?�LW���)I�M�+��:�?������W_<p�eY�ԃ�%�3m �8�G;�8��#\�������_�!��_�G�t�ā��jZ|"�L1M����W�COO�h����I0qC֖�3��<�$Գ�!���ZD�,�#T�� ��'�

(��NA4�R���P�P-a������ނ��8���	IK2�	ڇ����B;�d�eP��JYN?*%�PW^�7��bim�g�������E�m{D��?���w�1��Ȓ�	X�a��Vb�X+Z��!,/�j<���u�}�Q���B���+��V���d<��;�t2M��Ve�$F���D��6'x
�y	����<��p�EI��Ʉ5!��!�~	�v���[E`��v�u�a��ku,Y��\VX!v��!#�ha���눦� ![��c�=�r���)���ҘvbiI�g��h��)��>R��]�\`ճ��u�9V�y�-[�����=�$Z<���r?�O���Zv��z!��D��x����[Q�=�I�g��X��G��`H�JX��"2i5�`�z-��;$�K�m��	�_��ב !2I	"|L2��li�P��X $�[���b�F�\��� ���$e^�ar��:�RY����"j�y���	�!���-W^��?����F�'n�\��_'q�@�$�T�;Ȫ����o���߿�Nw_d9�,=Kr�m۵+g̫yY�����퐎0�ν��W�aw�4)��g*�f��'k
7O��p���;���X $��aU6��w��}��͍F�>���q\<���ۿ{�ez�puYEƫ��x���dB�X�����X%}�x� ���(�bx�,*� �.�F�2qsR�G%dR6�r	�_�o����Z&)UK�d�T�4�=��3wb߾aY��QK��׿��	�����"2N��T4b�D�n���u���Gd{pm)+�V�l���u��}�L� �(���I���}�f�Fy��58���ig���طo?���rt�*fR�}?����#5B{����������Nd;�����Y�4���j�-���Kz5�>	^��x=��#�/����h��L6�@�eU��9)ai�D���]�B1�D�x�7��c��شq��.6��<{`&�͝�Lf�E۬�$=��&�p���h]�q� l�1��[wah��0�D��Xl-�? �md����`@��VԄ���G���!��ͻ0R�P���"ӥe���a���B\�ժ�2bEڥ*T|���y�v�j���5�k�ۣ8��KZv=M`��)s,"?�Y'H��,�K�k%'�>���_�v鲾{-��?��]�cG�S{����� ٠p���������_D�i�:쎎^��E�쪑��C��ÒW���U�1�u��7]&>�L�'@��N��dZ�PS���P��L�S���/��3�7��0{vy]aS�� yQL-�W;𳇞B��U>;s�zu7��5�����# �A�dO=�?y�	�V���hl�NTY��lxi�OE/`!�]t���k�?];���M٥�2�;�G���WT���Sg�����p��KŵY���5�� 3\E�픀�#�߿�w셓��$j�u���҅s�xQ���wvvK"娖b(�Qs���f�	��A ������h	���M�]z�d��TQ��Z@=�lێM�w�v
ҭFS�j�&&�ߝ�Bb�ȒU����c���҉f�'06R�r`�<�"`�Q�u�l)���7!2^�,YB/��e�?�SX�9��b�����kw`����x����|!���}�>��]�r�3MT'�3-�B��X�	�۽cJ�*JUƩ�=J�P[Yv�Y�;���NG!��_�5�L�N�#E���w��w��87݉P���Z�IF(�N��;�ό��2��S^J�ǘ%�5�"�F&httD�f7���H�|�V�dd	�(�$/�+�
�wnz����������-�u��뤎@���Z#D����?�;�~��J�z.�ԑ���u���R��/)u%�G&C� ��/���DT͗a�ZY������ �� H�\-r|h�g�u���ӕ�x��μ�$G1��:�F��\��%�S.3@WjN�]��
Y�]��:����\�c�X������,�B����[�Zp<��(��;�2ӻ��̧��ӭҁ/�Q�f`LĎM�ץ�*�S�ɘ=�K�C�����}J�pϏP.V�k�~��q+��܋�z��r%Q^Jq�����s�!���XB6렫�B�
Yd3)	W�>�@L� шG�� �j�RQ�E��J�Z]V�V"d���B��ȉ� gp5���w�XD�TGGG��{
�=�t�������&i�A������ ����3F�J	��(ҙ�@`ioء���A�F�f]��z��t���9{���d�l��O�>��+�A�V���:��Q��z��Ύ�0�<���Z-����\��T��X.�X,�Z�IK�V�]�nZ��0o�v�E��/�h��.�������&��!���88\�E��?��Ͼ7Ӆ�#��E��Tш�N�cO���1���D�qJ����t������3 �V��'K�I�����6�c�~uvu	@�
��q=�l�`oW��?���n���Y��AG�����������8�S�\�����߽v��7�V�?���i|������$jR���)�z�vVP���;M܃M��9�V��Vc��X���l���X���)j+8����j���fD�����L|,2����J����Μ2>nJ�sBɂ�8��L
)��'B�9uaRN����3��$S]�s�4fP��f$<�-�Ԛp��eSR����3    IDAT�5��?����e	��yqAp3A�Yb24ٔL&q����^�X�HZ�WP8-���3�3�\�ۼ��<����>���1`�#�]�h.�������n2iW��&t�����iE-L9�V}���'�s�J��Y��YN�#�9��;7uU"��bTj�^��+���	(��8Խ�|�U�!�l�5��,��)t��*�8���4�I\�^<�*��p_�1��(K��|�$  b��;���x\�N��Ʀ+�l�x��hr�Z�U����u�8D"b�v�Z�k�����_D/���nƾ�E�1�o�҅�z��t��K�q���Mx�Fǰ��ƮC������%���,��O�D���8����O����?�\NN���P-�=]�rid߳�{�[���7\��i`��-���)�6:�:U6�q�#���������_�ʰ�ŕI:��H���F(T9�a��������X�U���������NDק]l8�A7��f٦�_>�$R�]$�
��Z�����d!���J�VgǔLE�n)N��(�e���!��r�` �S����R�������VͲXnN�N�j��'q������y�����@��z�F��D N�l bY�"���E$Ò�4Ѧ$9hry�)ӊ�����Kazw���ض�pdK�!�`*蕎�$�U��\Ջnǔc)�M	�!;Q��"�&0|�'ӳ��Auw��$�2�h4���&�DC��Mp!�YLO1e���P�e�0�Ô%`�m�_�:���-N�
bQQQ�Bq?�%����<p��~-���0J����+2=��v��A�G���	����5?'�	?q#&��/��f�sm9n ������n	��z �d�/�M�w���[��!#0& N�N��L�ة�B�ڞf<AY�y�D��9�|.�����l�+���10�~�����g����"&���땡��^u���7�9��,��~�u�F��^ŧj���=��,V���v�X��fr]v��.(�sPgC�g#O������ �VW�J�����Ihxݝ�$鴘�e1�<�e�Z襅>��$���������L�,����*S�FR(�*�\21�R����Ȏ$%���7#��Љ��k��Ղ*ҝ���W���=�k�:9���ʕ��s��w�`�@�<�ђ�zP�tk��!��%#a"$R��2�f����y�e£�	ˆ��L�ԣ��t�����)�d|�GV����2�Nlu�� ��l�-�8�k�Mr`��S�K��'�(,U0�ם���h�*і�%L�&�' B�#��Ĝc�Fk����lu�#H�V#E"�$�z8I�;��F:D�p��BEwv���V'���0��^I��.�u��hvdO~�
�$�Uh*5��@h��*�9��tQ���u�1q^��)|��H���:{a�&�$bÕk�)�n*�j�M� ��s�����1+g��8�*�nӱ]`�I�4�[�Kcdd���
 DAi���/�����;����Ҳ���>��o8�h�����8��=���3����<���7�vn�e�-�L*�z��b��ƅ��2B|�K���`ƌ�ˠ�CWX� �I5yh76Sv�4�]�S����E\Mz����XZJ :I%�OfNN8�T%d�l���>?��M'i�.д�NNH=]"(NLl!�MEt+)RV�T㲜�(�ذ�l	��3Ѫ�͟Q��x��J�"{D�Y�c�ǯ;�\p�iUeb�d̟�V@�aA���H���s2{^�"(�M��ɒ$�+�B��ލ>;���������B�'���R���\�
�ƍ�d�ԇ��<H�e��d�)i��m4�ACIY�4�k�(��0[�̈1�RF�*���\ԅ���F!A.�" �k��D�ȵoZ�5JD�PM�\1NT#?)1%��7�M�05t�R�<
p�%\���`�L��L�F�ꡮ�~Nr������.�N�s)f�����j-Ě֋�b#b#1\5Բ�����x ��`T��TO(�V0�P�Q��2�!��ɵ�d�ά���E}���@h[�����������f�ߒ����T�@���=�ێ�8�����W���p9��������V� �>p��Z[`��ͭ�T�B����	!�1k�l��)��<ԥ;&)��>h|��8�)�ա� e/SI�a���?�^#�N'b\�(|�(T�ɒ=�1ѳ�.0�-��AY�eN��I��zԽhG
i�uu��.���R�c�W}�]W�-�X�T)Z�P���
���m�>�7R�5��قcd�'bYҔ��h�v8I&�Ɉ�{g��y�1��Q�2!�����%-*d�I��CH6E�U��녥����shZ������k�0J:)�d�,u0���L�"�l,����K���DoDP�ϲ��8i9_2�"���$�]�.ϥ��L��ď��Eg��'Y�	iך6�9'㐈�%�C�*à��sB�(���Ҕ�x�J:���me��J�m !�"ZW$)]�2J4L�9��!�O��?��cO<�J>!�l�]MFQg�]-���ɇGG�ñ�y�n��Hږ��l��a��Fr��1��y��L��L9�d,����8����0��2kQ�)�}����+���?���������.���m tz���K��?�����/| ��W�+x��,R�HN	��a��9�pB# ��"!�\�fA6����S�Ĝ�s�}��{c�w��k��fbS�>q�V�������<�L�|o2I�0Uk<���E�L��hu��c���O��ҥZ��X� �a��%űR�!0�ޅ�
q9��|�?HJ9a^��BV���OѯG5#�� Vz�4˯��7�?[G�u�ui���yi,��^7&��L�cS�[Ʋ�CMO��>��k�4�c��4�5a�s�������:��s��o���#��P�	.Y�c��[��:�>����Y&&�"���$�,��*e	s�����Z�J����c�-��Z4�� C5�����@=ـ�.�~~�U����u��8�8�ɘ&���>e�ԔS�e�{z�<nj��Q�V�wϛ?��w�r�.�x��`g�U��f�y�ɹ"Ndڟ=%#���t�[���;�؅KB;㰛�+�z����՞�ƚ���]EQ0L����{qE��:v�|�L�S2��m�G���V�g㵢���੿;�D�Rr�.-k ��k�s\|��.�߱��!�y���E'eX�bK a�V2�Φ����/n���`;�sQc���N<v�^g��"uÖ `�Ϟ\s�\h��\�R3���M	�O�Q�J��R��J��ё!Tk�R�r�BC�>h�3���h�'6�rOq�Ò�a�dQ��/Ѽ�ět��l8�p�ciϊj��%׮oY�x������[���Y`w�ع9�O�9z��k���@�s�����������v����
�b�Y��I��=2j8�W��O�	�3g�K�Kk)������!s�n6h���؍�����$�&XmMM{�<Շ�!4�u4��f3"��$%&t�Qy_>����KHB$�1�<�i���� !ɴ��ITKHv�]�^6m ��S�:7����P�y��6�i����v.����P�A�yĿ)�Vwh�J�s#!PƘp�J%D�Z�n5C�
2.
���������N�h��WB�9dU�d�������8
Cߎ�!׮�����喛~��ªp�];��?��:9W��ܣ��N��q<��o���o�u߻,�s9���ri
G�)-p١tFH#3�mX��ԍ�l�,`��K7���.���C���ȡo�&�lrES��Դ��\�=FD�˿s��Ycǘ���*���������ڱĪ���,��/����E<D!?(Ŋ ���w`ǎ�թ���V�X���]Z��K2i����� ���������-)��Tcw#�	��"��'��\4��z*e��q�V���H0��� B����aJb�Մ�d��Ǳ�Y����q�.�N�="+�Ҙv ���3�kŴ�����>��W���׼��Ǻ<�0�N�?3�R��q?�����;�����7��+�u~lg� Jĕ�>��b��|R�j7tR���E%%;��T�f�o3��0A�_&;�����$5��㳟����ƒ�mS
�����3�ubZo�O�.�n8i�B����te3����<���KnTMHth�/Dm��=�KXlܸk�mA��-��KT�A|����Wr�?������E�ܹ;w�1=-&ҙ<ҙ����pA*�BͯH�H:%�F����2��ࠔ�|�a	�Do��`Rrk��8�i;d��x���A�c:<Ku����y����X6G���8�k�c�e�^ܓI{/^��k�z�o���srk2Z
���\uS�0'wL�Ci�T��L��'ֽ�o�����+#;��56����%�:2�G횒^"Y�qu��#6�帥e��G��k�5AP���6��.�ı9��B�H�uB<����R�]��W���|V����DB�/;������=���"a���U�:��B��.�̓�s�,̘1M��a'gI?+e!Ǖ�<Fw����m�.Ed����t�q%`{�jvpY�W�`9��a�#@C�ܵ�J�k-@Ȍ��#��!�e-?��f�����&�]	��.>F�qa�^���H���rΦ�.=���ů�/XSHa;�b�=�d_�ǿ�6:�1;+>�q~��W��_���u��z��Z�� i֎>��e��$1	bj'-��NJcf�����a��C�8�y�Z��wʳ�}i˅f���s��4�P���	!�f܃�`��M�9s�љ�
\'"�d�blb���t%6�������X���|O�dP�=A���x���ؽg?�̘13���ECL��weW�������'�j��(H��/�ö;�ّ��4&��9�ߊ�pL�g�\E�%DدW3Le��πn���N���[��uC3�Ǝ�8��A�%׎�]7:�Jٻ����^p����]zыK���P vik���]ўm�ι8�{Ǳ�(��O��S*��]���r��(둲�,�Z'���1�>/e1�T���10cf�0�cD�b8����!�p���&��m0t�k�h@��UfQ��<=|fL����s����~x���,a�Z�^��i�����	�ڌ�QO�~C��!s(v	�²%*�gV��¬��=k�\Gt$[F;�flq�kE=���H�x*+��K^��;waժ�ؽg�䱹�;L����d���^�?a+XW0#̤ �c��Z!��*�Y�) ����QQ-�z֮Y3�W-�?��f��/\�}`N�|�3�A����wC�4����GG�8��:��_��?}����� �c_JB&i@Ƕ걭��P�
����O��6(�5��V33�i���L�tO�w��q�1C�keW�z�N�GB<K��h1�K��s�����>�м���18�����0�vs��:@f�1,v��عk7/^*��t#o�.n��a�p��>�P��R�k#)�U�c9��۷��'����{��v�T��7���1 8'̐jV(�O��UGL,Us�E_�/���c"�d�+f��>_���^��[�cLVX.��|��|�w�/�z�d�G�v��p�~�@hj��ڻ8��V�������?�'��/��\�\�c�'���'��i�pSᡁim+Qlˇ@| ��ӏwr�,�lZĐ�ō.���K�K�+mj_�M�D��̣fP�	��#|x"7V�2B�Ǡ	����ӯ�b��j��MlB>��7ے�	>��!ho�F@�ѱD�8��˱�\�`ΜsT�,� �Hc�i�>�2���Y�M���,�UktU��v�ރ'�|;wJ��j� ��Q�ָ�,&�j�H��(��%D�8�@�<N�F�:���r$�if��,?�VA��s�|�����ܛœm�s�i��ԞaN�`�Ծ.���H�������ի7�^~v-�m���v�Z��sd�@(q� �I��ݒ�,�i��l�A��O�K�Uli��H�@��h�z�l�W��ԼT��66�����K(>�-UE��4#:�etvdq�yK��VJH1$�$�'��@���pCL���R��^jǣ��"G���պ0Dd�0�A���JR�q�1k�њ{f�B��}�(W*��� �y�v<��'Q,V4���a����B�2;��X){l�è͡��CF�O��\O���������1�s���=�4��,��Ր��1���׿���?�|-cY/�Ԯ����L���<��ؘ@_�{�7��_yg��\���f�)]�]��މ !�%40�7-%�B��x�eDZ��?�#In/���y�Uwvv�~V���vG��_Ň5�|r��<Ӊujwt,ů�PzF�+PJ�̚�c֬>�X���\F���'�����	�劑��6#tj��ܺ����K�V#�k��ø�/9d<���U�nZE�$������j.��d:��S���g�١�=V0v���E�v.����>s��8�"���I�Z�Ϸ�5��T O�}h���ʘ.(ˁ=�����W^�����[��Sy���>�#0�+���D{k�n�8NVp�g?�/��r�7�f����Ҭ��*��8¤v��Ā��ፐ�5ew��@kl=i�7!;��� �"�g�0��Uc��Zc_��S7�G��x����R�*m��ib֐�,,^4W�PT�S�bj2�2���u��6#t��c*�^��x$���$UK�t�i9�8',-��3ARnח���R�ҩ�w::P�}T�Uds�88Tƃ>�}���/��%�L����e2���D��K��@�X�h���Ui�gH0�=�W��3N����S���M�,��:�L)D�pɵK��_~���h���e�Nb�폜�h�34��k�;��/7��_����+/sӝ��I[�x��3y $n���E��4���}2$��!�� ����1��3�
MB�/�3�H�8x���%>2B]]]�0�ß�pJ_����	2S��0)�H���/G.��?&� q�NKa�G[K�;	[�R�
��E:�G���)2-
<��� DYz���`Jq�(��i^���4���6uv��b6�Di��=���=��r�Kȯ�J�|oo/R��Y��100}}�P r(��k�}bxd##�صs6oފZ�G.�!]i51o���_��$_�gmq��Z�b����O>��.�j�&9�g�c�������v#�V��%���o�{ӽ?}�-��[;�T��[)>�&�hͯyTBS'&|�e~&�	� m�6����T8�)��Q��xFh� !c������aN�f�#����I��c��Q�Kc�!��^r\'�ؗ.��$,�8 �lw�1��R��6@�wq$j��=�\%˨抩������XzI ��k�������� .X���\�T�J��y
�)�R�����l��h��EX�p�9�3�@���8�ึ�ͤCZ�-�ڵ�n�FKBl�������$�ȦS(��g��3�y�M_���t��r�E����,�I_g�1�wU�˝wW|�s_�i�杯��9�]��j��,��RhNk-��!�P���V[����pP��2�0C���z �a�z��wj۹��8ttt
���j�D��١�|�O��G�h��A���� �+Y�ƛ���ʡ��h�r�߷nQ
�y��E�CiW�a�]z詘N[�
b�'`9��i-q����V�'>�'r��Ϟ�PQ�?�#�g�a������)�����i�o��,�h����n*�z=�O<�u��i̶q٥�bٲe�L;�� ����O@���#�E��
V�~k�m��7��C:�<v���!@�ap�vܒQ� ��qߟ��O|e���-�����l��S�l:['���0텭�W}��_�sϽp}:�5�ݔ��[���j�)LI��<t�d������یe����,�Ny����    IDAT�a�][>)]�=O�bK�v}0�k
zuUJd:���.4�,���,]5��+�C�T����ý���:��%0඙�n���m�f���G̲��]�w�g�C�x(�=�B�ۤ1��"����J�l��v��N2Sb��d;�oB~>�=K��]�Y�`VXMR�Y�w��	��_��*;kBzoϫu�a#�lyּ��y<��#t���,�?��<�O��()�)j�� X?D.ۉr��t:�gW��/~�zѓ�^�����Me���ى��KZ�$t!@֔��R�,�E����V ��=����_}�����女m�����{O�<5����<C%`�ޝ�W~��>����_g�z�Q*�ʕ� ��X�g�|$�e����ֱ9�
0�>&`�e��J�)�� b�k�A���
�ɚ.ƌ{�R=A%�僧��/a���QS�M���[��ͶLk������* j��DԭN��q� L��Gֱo�y�=I>�	�(��5ܵ\�`�ipפ���q*O�Y�+l��J��y�����1kf��OdB�W{���^�b�+��;w��K/��8O
���L0�8|�@,�冨5�RY�DK�
rpp��{7mU͓��\�t�}�<��R���>Y��\���L�{���q5��⁎�u�_��?�ڼ�4٠�H�\K'��m t�#x�}>�c�L9P������<���J�x��ez����ض�l��'����S!}i��}�1����#5۵K�l�*�j�t���#�b����	�,5a�Wa��$C��3�Df,��/�%2v��dt�)�q@h���q�>Rć�vQ��T��Z5M����ӱ��a��(< ],�U�cŮ>ܙϔ�5}���]���,�����3��H�̜Ѹ����3{:�-�/ (��<j��Hhr#��ԉ��N��~hhH��]w��MCq�������lܟɗ���ℨ�5�r)��r�`n�㤰{�><��#)J��� 
pa��$,Քޓ��J[����;��-�ɢRa�+FGέVGv�z��o���7���2��6t�Wř�|��q?��J! e`уn|�=?~�e��oZa�ހ��v�pR�Z`�^�2�>ʆ��\�K�g6
�
�=��׵i��E�3�\��/l����ٕJL�Ƥ��	u����z�x���BdX�ܭ�������"� S�l��?�5ޓ��:1)���r�IZ�c*���!V.��es�F�,��؂L�ӴiӤN����t�$,�	0B�p5bu�6̐�<�}t���*^t�rdR�8M�|i|��E����Hi�"�������G��Bk6��1��g,�q�Ev��P�gc@�����QlظY���ta�|��҈�1JE���L��U�:"���ɢ�Ȥ�ߎc��_ڱ|����_|��=<�����l������CU`涝���7���C��x���E�3��Q��>����9A�k~�p4�39k��e����՗\r����l�����[F���t���u�R�(d)�dф,�`E��`�cl�het���=dYZ��Q!�8,���a��-��9�D7|���e���#��"дl��ʕl�zYJ����e;J�X�&3DF���Ψd&u6�8��It\��%a��q x%r������%<3� k@��Y����=�{��u�A �SWg�4���
�x%O|I�J��އ|�3�h�LN4�����{Fy�h��[�0��z�5�?�D`-�e.~�+r����+CQ�������������G�kY{,O����or#�B���̧u��V*��v���k_�8o���Ӈ�G��G�y�q=G��"?�͎�3g`�y�.߱`�9[gOOo�=���yݗ�������K�a�-�kHe<�&@Ȏ�R���"����@}(�B`��$_C��"3D�Yd�������c.�Ej2A� T��f�U�e�KeC�a�",m&uΟIl�㈋�1��/Y-�� �$} 3�K�t���/%���'G@�Cm��fsϙ��sg#����]��>�?��Ɍ�Ѵ�7v��������nI�~�!�C1�D�H�S0=}��\��o�A<�����i!��1�����%y�aH��1ȵ�l���#
*qT��=�{oy�]7�x���ƶo�d����6�:���	��X2�]!�Q��P-�r��� �R�����T����V-�
G�x�#�z������V�� ʸp�����u%�	���(�"g�G5=3��93v����!v�pP��#�U�EGCCk���"VI�k�XGG�j�5�n�l�p�e�t�%�tm�#��v��R5ڑ'w�u�lna��e���,)�\�5�Ȥ,Y<=�����k�	��������P+��F���ǲ�����L=�J�r�s}�m$ek)M�4���C�Zp�����{��-L�=׆�`�kT� 7a����	.$�S�Q5v,�n����K/���>v�]]��,�r�G���T�6�Jgc
�K�#b�$ɸ��K������8�z�ɵ���g��?�_Ĺ��e�G�biLه&#���/�$�١�H����"O��-��P�1�����i���9�����\Eևe:Cת��V�>�j���N��xĴ�Ji��G,�%�to,����h��mJ�ҤμB�S��Y���J�š��� �Y��% ��_�8##��G�μ���/Z!.tę]J������t-^�6X�@�ӟ=���v 
B�L�r�L
qH#FMFH|�o��WҰ��������K��䓟��w�NK?aY�������h��:�����hӮ�+��/?��}�vR=��N����4�|+j�l�5Bi��l�^�Ǝ��dz�DE�� �g���o��n۔�d(��@IǓ�3 �]��Q_�0�K�Ę���p?|q����f��������Ӫ��1���ưe����7��+I�]2I��߰>�h<g��ϕPV���e�s[;��b��*��=�0yd��W�%ϓ�K�Lw&�c^*�{��6oF("�Xn𝎫F���V����+���W%�&�������]��~�#|�]�.��(�}m]�����6�����+j��>.�ӿ��{7n9�bř��w[>�xtl&���ib��"�Q[��L;IF�P����E���}�N뀶�
�ݎ���?��C�D��h�m�(���X^E�`X"�������L����y�<ʓH��2�d0IL�����( ����i���@��8JsŝAgG���I�lZk6\c�Ϻ����g�������!�ߟ��i*Jƕ�;�6n�&��N�w�b���|2Q9�+| �tFLa�@�st!�4��ϥ�Ӻ�������e�� ��n�?[����g}���8��T�w�䉷~�_���Tv���κ�6�b	���dSh��R��M��1~M�Pv�.��6� 	*�o��Z� ������a~7����bgC� *�"(�f�Zw���ح	~�p\-I��������E�n1�U�k�!�C!�Gڣ>)�|.+`(�Yz��R)�V-cZo2e�Z���ĸ���>?��G��� �8�Pu�K�����~k7lu�N�=�N��XUj-�u��>a�Z��lڥ6(�U��qP޾pތG��?��s
��C��i�S:퍟���Љ�^��cF ��5�n����-V����;�Ȕ��YZm��W����B�I���2N��g< j 7� 4<��i���oY8� 2�����d����i�eUH��2m%nt��t�M<�H��itI D ��e0��=�]��t�;DDֈ�Llv=z"����8+���v�λ�M��35f�ت7vC.�b���=� �l�!�d~�{�m���ˤ%~õA�_G.ぽ����p>㭽��������'�t>/�6:S��}�	LA�h�ڛ=kG �c�`+n���[|���\�g^��M}M�&j��U-�W��_��cKj�;��Em��5f�7��cb0'*><2�V{�F�9��>E)��o�e3Ӂf%[�m�f)�9��uwwb`�}�=Hy�8�Q|�cDA8tX�P�d�L��׭w�^��ɏ@sI����vO�P���G��{��GWw�F�0�5�0R,"�Ɋ&����²�ȯ�j#C{�,�;��W����W?���p��Ҽ�&?�4ǣ}T'8l�z��}������}��ue"�KHۻ9	��F-���t���ph>s����n���l�UfH���ugƽ��d���!�0z���h�@���Lcy�~CD��5�l�`��2���M����,tw�!b;W��u�r�@X
`{1C_龛�&e��μ�Fh�'����6����o�j����ھc'V�|Z\���_ ^^��(��صk7v��-M�L*je?��ig�y�-y��7��#�W��L�-˪���j�i��>�O�������8�S#�%�7_y��_m|��t͊����Ň��%�P����u4�ʡ�N�Ƨ�U9����Z!�ov`��K�c�Ӹ�/������;��� ��eE�V���[���V��0kf�Ν�ޞNB���t�u�SaѧŅ�b�L���*S���Ǿ��ȴ?��	a�fHLȓ�(�&�?�0͐,pll޼ac`� �{z%��#uz��Ɔu�_|��խ]p��W����/�p��T'6��m�ė��z�O��� ����G��3~������;�:/��T��1��G�Q3{:��jq�m:#'�sD}�5�G�pϩ���M�9͏��'[[�2��#e�I�؉y�V�`��p��o��W��S�f�C����d��5ݴ�=��`��kE�?of���	��)F��+y����8j��|/�Md��?��ΰX��?������B)�qQ�]�I���a&�DF��VM DSS��ٖtV�K�����/]��W^{�N��jk�ޜ��K~�@�%�O�
+T�E�鯾}��k�d��s�tέ�!,�� �Ύb:�&B�|J�4�]Y��~>y�	3b�pS���> ��!�i�)�}�s�"r� �n�`��pБɖV/��>�
�-���:�22;APG.�ET�t�\�8w)
���b3���Hd�Z���o�x���N�����ǘ����R�$!�y�a�{+�eGUێV^s�������g�m-Љ�����m tv���fo�8�{�������������+uLs3y'v���;1\,
��P�b�՚�����5�ՕKIA(m�t��EK��vX�خ� ,!��`<?S���(t�iae4�R����i�76�`����"1����v4�q����;����s�kx� Q�@�U�XDYT��X�dG��^Ǚx�l������n����Nvf��zgSf6gR\�7ɶb[��%[�U�B��	vt�[���{��� ��} �{���[��W9�/�ouws���?�#E���*[���\���� ����������o,��1�-�|�I��0j�m�����o�޹��!���;��B�ً[j&RJ�F��O����|�яOMy�s�����7���.]B_5[�@^�
U*8������h�kG�హl������P��F�N�W%��E���BwW�o�����_BHw[�ή�
ؼ���}=]���K��Kj)�촐#��	B薺���Yf\����%�.nʽ09Cr��t�ҸA���ر��kWv�X1�K� ����뛾Rv��D��}�����y�R�w�N��r�̑�I��
jN�������u��S�tS��P֡�Z3�?��Pet�W��"�1jU�Iv.ך��름�-C��%u�x웎Fx%�Pl�W���Â'TB�� �y�v�m�:�B��u�=G����W{�$�e�]�q��X]��/w]{���s�^����;kV.�ڮ]���D�����)�Q��,S���K�꥗������K�;_�E��);�~ M��wMS�?`ː�z�(wX�0ն�e(�=�Jzc������2#��ˣͭ�wW�Y�<un��T�W.����.��������tӰ����1��B�݁q���}I�%���݂��Oa�Q���=�~jkɫf�I�$�^C	't���ԘEbTX(�B(���eH�꨻�/��L����*�P�����s+{;������В�_C�ąڷ�B(}{r��HJi�j�sv���կ~��_zcW�ع����f-'cX���_�
bd���凅�n%�����y5I�eͨ\�>�n}�k�Տ��ٱ�����:yj|{Gg�U�� J�������E��^蝸
!ĢF	����"��V������Cd
>qU*Ai��@V���D�q�XR�~����
!Cp/�l�ck疵7}{�[�!oӫB��ٛ=2���&�D��!"j.�~�����g��z�׶K�Y��A��FƴSSa�#&�H9�HBJJ߫DQ5���[���];��r�����M��o�5��/�곟�*�=D9������_�Yg�[BH}�U��:�E%�x(�=0�O�/��U�2~��h�գ���c�^lKh�:�'�^�V���¿��WV�R�_����V'd>g.�*���6~�!����9� ���^�b�l"���
�>x��m_컷�:{~����*ð;-+SC鄑4,��eE��Q�{\?PQI9�����@���ܽ��o_���Љ)"���O}������v�8�6+�LՁZ
�u���I�z���.������|�����-[6��]ەEH�;���Ks��b�8�1�$�t��R��n�`����p�=��Zu��ݻ6������\�i��)# !��Y*��@�Q�A�w��к_}m�Ё#kFGƺ���R�媵����\&_*s����X__��ƍoۼ�h_Of�!:OD�B_J��ʁ3�����702�ShZf�>��8'	���֕�F���]�5���,B�Q�QNa��ro�={���6�o�n��TԮo���>�z�묞�I� uE��\�#��R:�\X�������ȭM��r��=w��|g��!D)���� �м�ā��@�2k���'�kbl�k|r�ur���}���ۦ�:Z'�[
�,M8�sD"�՛����#��?�?��_���X�K��愙g�R���؄�l�J�E�]c۶mQ!!�e8�>�o�B���:�����י�B�-�,~,����o��B�9��EX#�+U����w�7�o^��L��AA�[�̙�>�-��~�z��(���n.n�ޤҽ�O�\������?>�Δ?R��aH�9��)��"����I�����5�jU}������m���1����7_�qV׺$��Ɂ�u�k�Mi�'�Ҫ�j��"_\m��PU��Rilʲ�#=��OmX�x[��k�uoƢ� �Т�:L�b\)o������K�?i�-=~`	�ՙ�`c�qB���N[���4�Ud�q�%Ua;T�I�� �������2EAu:kl:C,��{����Y4F��&p�v1\,є�[���nȅZ9iޫ��H�C�mM��w���wu��ˊ��D4� ��ޟ�B(�{�^�������O}�_��oZ�o�ˈ�EHg]�*ӱҹX�.�ȱ��V�Ԯ=��f��G��C�_��R�T�f@3t��VXD.����-h�7���l?81>2�5�1E�T,L��{z��o-fd2t��*A�h��q�B��j<)e��{�O>�����a��56Sc���TL��ﯦ��I�%fD���M[6��0��V$q\P,�-I�����f �M��z�͆�� (��R{[�Ow߹�ۆ$���o?�Eæ�,�(�Q3h��fqBhq�f{\���8��̟��ｹ��/;ٖvI��E&���F��_c��n$�Yb�Z�M��w'9NܧmN�D.�[� g	�^|q堺��!�D�pkK�ѻ���w9�^��! ��>;�euB�B�M=)�p�6����o����>e9��"���	�
AV!C��8f誯�ˤ�>~K    IDAT�z�1�K���t��L�~����q_1�,�����:�I.0R!g�/��njo+R>�Sru]K}�skʭ�X'g檊��ZVҸ2��Y^�rW�>�����Rr�r��_;W.�}\��35�.w�񗄤g��!%����28��Z��]�l�rV�÷�`A�B��27����8tj�#�g��w�A�=��d˵*555Q�\�|&K���*6�s_�Yeh/>��&�3�������t��A��gD�.~8��َÉrU+��q2\[TݪY,6	?�U�[>,���t`�R�a��Q���t�=wQkk���PƱȱ,�bϽ�������Q�Rdp�F~l��,i�t�i�6-���M��
P���Y|j������wWS��t�V U$�f��k]߭���55�ϗ^q�Gz��6sޫ���٪3�14��%�܋��G�<g�����\]ݶ�0�T1s,�l��2��l���[�[����`x�� �pR�r�=6x&��/��s�~��G����7����	*�s$����K�B��ߞ/v)����n�X��wt����Omɩ{̢k� �
��@���~��eFZ�Z��k�+��r���d�w�槁T�h�eĴ,e�)���5t������J�JI�#�W��qL~@�z���	]���0Zd�uL?��%�H��ń�|!�AAT.��O�p�B(�����B(S�ܩ���b��/�i�y_��&{��`��e��a���O\
B'D&_F8�R�x�d�Q��n�\q=$�.ko����_�l�7��jʁbz" !� �v��{�V�U�?��������:�V\�p�t.�S���&�3��K]
����=[xֿ�U��ǝ�W�'bwW�o�v�r�s+d�aɴ������������03ۉr���43�"�M�J�K��1�R�$���h۶�4�n�z ��c+��e*�,dw��陙ܘմ(
戈����ۦ�.�3�p1����ӻT'2��.@vA'��_�@���^�}�N�&�ČE��fTgEMb�T���2�/!S�$L����BH� ��?%�~��_Z�SxB1�M�K�¹qK�*ӧG�{���٧�&��+�ّ˷���蹿��0O3�e���z�ե�Ll�xbKQ��,1�ą9��� �Y[�t+U
%�VP��9��������G+��?�������dl,�aY-�gY���L>K�Z�ܠL��<�HRyj��,�ܹ��߾MU�����6���������J×ZimV��z�׽'�T��du���bv�5�bs�kl!���Ǽ!T~չ�f�ۙp�c������ł(q���l)e71��P�~-
�Z����vggۣ7�z�ɡ×+�z�u��:�[}��������~�G��ů~�Sͭk�Tk��M��W7N�#J.����x�DB���������+��۱����P���+�:��1���FZZ������|3������|�g���ǟhtĿ�u3݆�ϐaaqYܐjn�ܪK]��T)W��ٶ�6ڲy�YrlݠU���Rd���.�2Ү��!������U�B<}����.�qfNK����e_L�=��=������c�g����U.(��|���V�?7��X�8#��J��V�2�yh]��'������|��G��I��f/��J)����O?�׿1x���i�,##cr܁֔k�P12ud�-s,C�i����7��0�?4cምc�E(� g��r�Q(M�����|�_��C�?�%�nܔ�FԻ��S�}�������=����AT�������o�B?��g��MM�n�Zڸa�l�$�$�h
���8����KR "�����;Ed:0y��h�Σ��A�7/t�\�'.na��z�z�����cxf���ׅ{��Qg�K,>�]�9XZ��(���H*s�e�m���0�2���$á�����z����hν-����U��K� �"Koϗ̊��F����O�����_�T�;��lq�y���شn����&q�Dͤ��[�b�Vܹ^d�{̢�{�I���`ĩ3�$+��u�V��������G�U�i����_q���q����>}�����}UWn�曗{a��ip ��y�E���A4��d�qX��Z[��R�S�d��!G&�!)A]�j��@��.�A�5���-$	.��o������ț�2�����̥����U��{|�ǹ�r����H�}��#����
�d2�=߱�S-��aà�����rt}.�-ۦ1f��P��?�|Y���e����B��.���*��]�V�I��زR�h��}�Ǿ������Ff��##�+����/}�8���7Z�S��9Aɭ�-A�EH������$�b�|���d����'�l����/��Yz�b�^��GDy�h�}�v~�����[�w��%a���1�����L�I�X�^vp���b���
�)����nZ�z�w�Pի��%=�>t����l���y���4�Y����M��c�#�zf�����B��_K*pY(ǰ�;�d�o���K@��&ט�z�5�ĐJ��|���uv<�q��S-E:7<\m��0�0���d!��6�#9�F�ԟb��c_��1 ���^/ٕr�tŧ-_��>���>��V�yS(�&���'�lM�X�P�u{��Z�xdYqL�2��p�^�w�rK�1L���
���1U�C��k�E�'ӈ��]Ӓ���/����o>��f�P�����I)9��u�B��xq����}aׁ�lZeZv�a�92-3�BDl�� pE��4�s�d��Bϥ�eҝ�wѶ�[��]c��S�]c[�\�U��Y�_�-`IlU}ݤO��5~�����c�E���\��,�Rr���NͤM�u�-�S����%�@�\O]V��gb6cW�J�g�Z[K#����|�K�"!kxr�j���V�E�!�����WϴϮX���=��)*q�\lhbj�뇢Rt�O�E;�E�u����x�w�Uo�����O<�Ӈ�J��|���2F��*����u��12,C�0��
��]���[�³�\P��]]Z�&1,
�Pes���O�_����#O�߰��O��G߰��yʟ�ڛ8[��D��A�����<��o;q��ơ��5�ew�v��"�"�0m�"~q=�v,��
g�5����G�˻8�Z�˲U�N�ZU֤\.G���� �O��\�6r%!d6��%���m�u+�|�0nZ���,����Oj%�c�PH�Z���|�Ѷ�{��c��U�����6l\�L_���>�36:v�!쵆a����B�![L#��/����;�ܜ~�m�]���<_'l��� �м����L@JY�Ц���<���Th�i��i��A~�13�*��-m�i7W�ܸ�ˌ+4�D[a�`�ə-�G�[�LFF�V����۷o�ɧ>������|�@4|=7�X�>�;<��篼��7��??2�I�<���R��r�aX�aQY�܁;
C�~�Z��{(�8��U�7oe�P&��
�,R��I�:K�*��L��"�c�f�k0#�̶P�ʩ�x�����u�BI�c��C��$���'�
)6�z���󸀧������"�iF>���m[6�S�֧�)j>}��{���kj�r��z��".�����FNf���|�~m��O��j�y����\'����űO��<�R��<Z��3{��{O>82Z�I�[p�a>4L\�D���ISG*�4����I���A��!)�j�J��V�mpBKh��x�M�{ώ���o}�ǽ��9��j-A�Z~�2kr�:�*-;y��}���{�wdd�cb��\��MccYC�s]�Z�8��X����}������L&�Z���\��5�Í���KZ(��θˮ.F�Y�c�bH�K>pȽ�LN�Uj�w�׬���-+^9yzr����>!��"�mr1̙zG��Y�tb�0�E������qtlY��'_�e�O�ܱ��{;���n�Dݓcs��'&+�Ϝ틈�e��L��X�x>�i�l=�����6�H|�̘f�k��\� �Ύ%G NM�{�壻�x�{�9z������L���v�H#&YvFe�%�,:�K����uN_g{���*^�*e���D�y�Rն噶���臞}�w=ߜ'n�8y�"�~��jV�
Q1��E
*N��idx�81>���N�R�LL�e,;cGA r�\F�XY�z;}/�E���׶�����Rڵ6S�G[u��^�	t1!�)�˔婱�a�c==�?ڲm�c�,�:t�����;�U�C�m�)=Ю��/��v5��{� [NC��ڪJ91`!Ր��nߊ���ܾ�K��Ȑ399������++����&a���f&�g��҈Ct����(�i�8\@ B'Œ$[RZ|��?���=�̝��=u���̶Ede��,�rT�!%{�\d,���8n3I�)\����F0f���{�x�Wy�g+W-{�%�L�ܹ�����kؓDf3�Y&2kU2�95s�Z�w�;��<����o%2[��0�����얚���ԥ<_9C��B(�B�\6E�N��ާ���x���z�|��؇�����H��dgHr�V,�8�$�0�~��b�:l5e�l�$����/�<����s��oor~,���p�󒃞�'�9��#��r�� �oB�M�[T�:T!�,�ѺW�����^�t��3k+�h���e�lSsH'��$!a�ŝ9�3�-;'k�'�B�氢ZUw��5{�kY���s��x�=�5��&��4�9H)�t����86�P��m�d��=_����C,��T��K��xS�٧�E�Ph�p�ށ��=O����Q[�ފ���c����x��?�T���䥴�Kjk�T��:�ܢ:)�dUĜ���l(�d���[fpdՊίo۸�k�C�x�/̘�M  !t c�t��J�
Q��i���p��o��߻��5�O���܎Z���}��MYS���]*�4��k�0���e���6m8z���6�x'��������BR�������O�{�����v�v��)��?-�tS�iW!�v��+�
��θc�t�gM�ݴ���뻞�I	E���U���Z�g�k��`|��IN!b!ā�*x;N�V%)�xi�W��]ٺ5�X_�pn}�d�K��R���qZu.Dyi�<0t��0��/2��ny���<�kǆ�j��L11�p$�W�j�DRL �札��D�%�85xnف��zNvM�&�TAj���$�t;��&�W�^�f�����g�[�\���]����b1�K)���=6�n;~����O��	kC�Na89ð�H�cB8�ǲm�w���r��M�+嗂��Lv}DAխL	��z{�_Z׿�'��+���B���G���W���H�����#a�R&7U[U�2������ӔIi�T3V%����d�W*�8�Τ�$K��#3%���Rӹ�e�5sI�L�Q���V��֒�t��K�^�t�_N_�^N���qMu�0
u�,?l���;�!��+e�V�M��֮��ʆ�˾Gzo�ޗ�{�v�;����&[J�I��������|2}�U`Ps��]Ѝ;��}��8�qEű��zj���䩳;�&�[J�Z?	�Ӳ�ð� ��0����C1yq��j!��e��-3tk7��l�:��^<������=�/暬MD��,�\��șO����M+w��eX�z`Q@����q���B3�&�5��>#2f����nĂ�ֵĵ�k4���u�.���P�rP\)"ǱTk-�,-L"]�s��g}��OBCez]J�*���+����!�|��߫ʦ�S�ґ�Ζ�����߲��!�yi�C����k�bY+�	7L G�OA�X,>ײx�|Q������hu�ٳC�G�J�ڊ���,�����9�ݐL�#��C��!J��X!�=��Z|����`[k��B�u4Ct��*�b�0Ϗ{|�g������Q�Kpi���h%��K6��s�Uֻ��Ʋ�H�v�ͭ\=�3Z5�t�bh�EH������o��?�u]���!۲�k�E���qE+������FS�>f���lN/���9=�*����B��Z��l&W+<i��~�h_wǏ�l^�hk�*����n��A  �Ұ���@,���)���V������]A4W�Z��̄RZ2��i��eY��X��iwt��)�'�-�Sy[���]�]�.Jߧ/�r�w'���B�����W0f5���bW/0抡� �Y���7�%�׻��j"uo��kMDq��ט�˒F\��PU���y���U�*mQ28�?v���������i���Xi17[D^�%q�)+�[[���9]>���Z�<��On�m౎��A���k�a�q��{��Xf	 �@bK[�
5�fC�	�lH�PH�MM�S2%y�ʶMS�)G�~�����Rʾ�'F>�oߑߎ��M����L����. �]q�D�{���Y1:s��f>�T0Ү����Ta4lR�=��I��T��Dש
C���M��H��U��d�e9��`KϏc��KK��؟i���L]p�,�7;�E��� �bW�F,��j5t��:�[�ޱk��ڵbw��B��n� 0��|��q< �EO �%��G��"��$&�d��"W����o�^�|P
�%�p�y�|���]�/�̭�ά��e,CuV��]Kӟ�;�������ug]��&�T���`��e��&B(
��椆Ic���/�v/;p���3�����pE���M�2TUt�?��]��;�1�Z�$A�Ik�8�(㑢PJ�d�{de_�ӛ6��~K퍋 B]�I�w�� �P
6S �� �-�h����_;��_w}�`�Y[�������,2�9��i���,C��uYS�9pI�M�%�� �1!T7f,���S� s�3%�r�A˜��J���=�]�ٵ��;c�!�odt��6	�j�RXA�q=l�K�mScL���@�>Z
騡(
�K�-AQ��<�4�sy��bV<�g��-�}q�,� \̋� �Т�2L�)e��I��_~��+��N���\�̌�Wq3���c.��F�o���t)���8�4�#Կ��n��%#�F�i����#)�ǅ;M�EY�-�ޙ�����ڱ�sy��U|��s����O�+;�鳜l�"�&K��Ps��̊c�\��o������Ҳ�����0Otuu��jE�OW�,�����7b�[:g4V�FBi��	@@ݛ���p���o����=����2� ";�k�p�ms�i��kqF[�ꂙ/H��7���>#���=�
�tuv�q#5�E��߀k�bB(��h���s�fǶ�Z)Q.��Tu�-�������W}.#���^wi̽}��ٻΜ�Y��m0,g�$3GdZ��!D�bÙ`�efَ>Ӕ�/�ג��s1!M.�����������^Z�j�K�[�m"Bp�U�@`��Z�[����� ���kD+Ϝ�z���c�*��q��v.#�Uu��nD\�O��Q��Öb�1K]L�ſ&YR ���*X��47��#j:�[;��?l��z�J��5nd�к��_غ���B��u��X�oj��yxl|����-Q(VzA�E�h��#aڂ#	�q���΁�<�(2D
��Z�2e��|!�=����Ɗ��WZ[���Ӱ-��o)�Bh)�2��� [<\�5�O�:p������w�m-AA�)ݜ-ε�t�y"�3�E��i�Ӭ��D�İbWZRK��&b(��B��r��y�Y�����k,Io��ߣ\֦(�(k�e��oߺ���W�<&���AR�#�-M��ɩʚ���U��+*���0��L�j�Q#iq�<��`CW�	�JD����������G;::����&�NƭP�)�F� �� ��0� 0/��Y�h��ᇏ:����.L�Ur(o,�T���h����.f�I���?�
IU;GUs��M�"�]J�r��$�餹�]���bm J2��E�{��Gٌ�m,ȭ�&�ڋ?޽�kk6"��\l�Xe�DE��ݭQg�B����{G'�{*S�v2�l�r�w䲙jkKq����T!�;���Y��>�%�`ס��  QIDAT�R|�J B(�;�y� \@�S�Y�;U~p��?T��N6�n���y܇+"��:7��];f�.'�b�t�P=�HUu6����y�+��&�LƑ�i�Lり�װou	��S2iW[�T�D�Dq�!�(M~����5+��}k�l�޺��Lu�b�DT�Z�O�Z�L�t�El��"�rf���KD!��aS��EG Bh�m&K���2W�h����{�����D�Z��v�l�q�F�Gq%fm��6!�ߝj�x xRJ�@�&����B!���-f�����wGT����Y1B*T���ulP���k���-[7|�E�w��w�Xͨ���s�D��J Bh���K�@�%�;|>�������;7t�aX�,+��y��$lۉ��A]�"4WT��J�T�2<�����5�^��k߾���h�$���_/�QI���С�mq� U�(I���	�-_����-�om�_������y# !4o(q  ��I���qcة�6�81z׻��31>u���zm�i��H��Ogaœ�/�Ⱦ/Z���
�Z�D�e�a���{��o�kkV�~���|S��u��N��D$�uDd����bfv��N�5���BZ��rQP��-j�_}}���/oٴ�1"���f�q�V% !t��,�K� ��jD�S��̓'��:��ZHX�Df�$#�m�4��8�:n�:�s@2C�ex���j�b8��c��;�Z��ooGW�ͼ����5��?{�O�*ღewٶczA��Ny@d��n��~��(�iY�jd�d���ov��Hl�)��O��X_O��k�~����
!�Kd��LXPB����-�,�Μ�4<<�qhx|%���� 2�BX�H
+
#�;d8��Y`���8u\F~�P�9?X,���y#W0���4�������c��ӵ��:p�׆��ߓk*6�m�^@´�v�<]kP��Q�ݺB�)�����4�\,Ƥn�!#���j�����zj���ou���@O��qVa��B Bh��4�	K�@�2^%� �z&'����T���X����2��[�D�4��0��=��A�lƙ(4��u���\�q���<f���3.�� m\Ji{:z�������[3�B�0,����L&K�H̞-A,���}$����e1�ܫV���Z�\sl1����캁5���̰B���@`@�D@ ]�(6�p�83��D�n��n�k.�jMU�ulۖ�2��cW��D>K����3FDՋ	���r:ŧ�Ǐ=��;��,׶:�|�ie�H
EB	!]�Q7OM~���4������]Uv���PPX��;+W�<����Ŷ̫����u�a6�� ��"�@L@����"G�`��$E��!"����^��Z[8F������#��8y�#�[��X���HX��M��,�t�GmR�mv�qlPą#��!�a��W�����{�3]��[�e
����n��� ��U��A @����n;:l>~d��sC;�&*��"�YF,��ar�!��hRi;�ű�2��{57
��|�9���}o{{���]��]B��>XB�GXbbw\�%ꞜΝ�z��-^$��n���b���i
���(
? ��r�4��b�9����Ɗ�M�a"B� m�@ � ���p�QA �(���)�]��/�׎�N��X^�V��0�F�`�����m��Bsa����xWW�b���<7R��-Q�X6,��"�� ���d��ڑ<�K/0�Ep�D����<i5͂M!�uV��,�h!�[�_�c�j���3�N�e�{t�4����EN���۾��h�9�9K�\>�.��g�i��0�
R��@�hI3��a��q3��A@W�9����A/���Ё���"��ം�
Ԕ+`�_�,o�5���M�A ����j�Q�:g�9��u������j;��I1@�����)�	 PK   �cW	��t bv /   images/a4ba225b-3a91-4e5e-8458-60f0fa258431.pngt{UT]�-�e��!���Bp'�������=�`&8$@��;|��_�Zwf����U����S��,��J�
�!'+�w
�����"������ˈ��͒��P��I�iz��"eh�g���A����ґ9\ب�pNؔ5V����������s"�}ǭ�m4��$���WQ���H��%q�\^)F��].g��dH�*�Uf��UmV�,{l>������)ب��ˠ��@�ㅨ!���x����4`�*�D�
�0��6^ ��P�z�"*���1�v�@���C��sd/�.��#���`��	Q�H;$v��ˑ�r�����/���=0d����g��˩��#A��.�X����Vk #������o��444�eee���#Јk��ؐDH�����sAYKi�W�P����jx���{6p*���Q��r(�.�"7��̮�H~wW��Ut�E%�+l�}�5K��1n˥�"f��o+�0��Ǝ.�f�mB�(**�nB�5�Cs�]��[��PC��5=5�z�-w6jjj��5�y�=DXS�VNV�^NY�ν{�>��j������J���5�L�<�1ZݔH��Z��}�b��f~;HTS�.�����%��0����V���8����D�ϩW"��=px��ӖRh����vt����{E׏�Ν�x�J+n!��d����\V���?<x|�:��]����$�\RBْ�J��;�j�S�?�d�\D��pRRjB�UD�*�`T�YQ5uVz�/��A�߿�����Qd�I���n���FV��ׅ?	q�p��l�+I{�n.1i׹���h��	���11)0���~U�ˢ�F��E�!]@�i�i�≥�W�LKP1-�\�
�?QM�A��R���q���p�-S�S�WU�Ҹ�-PR"��D������STV��b/۷7?��0�N��d��`��-�Y���L�H��ҭ�=��A�d��SS�i�,BA��=J���	�c�`����򒨏Pa�r�V�+�+è�K�\#ի���	yv�׉� ����BĬ!���.���z�����j<����{���-"BBmi�<wk��P��c/`�Ĥ��H�ұ^��}q�q����F#��_���� c���q�xֿ��zO:\�\��wZQ������T�4?x�u4��;�=�#��/���������9c�����ǿ�7���v�Y��3����W+P�-���@"�4$$Dا����	��)=t]�0������$�X����/���LǢ��=I�����椾�����ܔ\2��ɹ8�����q����|oN{7�O����� �ms��R�W�ްOG�Ϟ�ݙ�w��B�o�������{.�j~�ׯ_,�����8]��{f,��5$_�W����I����o���t5�.6�!0y�k���l�M�챜����=^>�����߿B/�L������'��A�eY��~�.{�������m���t��j@A=�lB�=�7�G�ݞ�S���n7�K����D�Ҿ�>)��τU�A�V#�x!.!��ǹ"~�zm��y�>��s ���A�ρ�o��k�N�l�0��f'&VoC(��	=M�lmO�W#?��ǳ����`�n���7�-��0��� ��@���	j�G�+�����~i��)X�x��@��K�@C���=}�J�>+�2ⱔ��j��rާ��s��n�3��f�n�6J�?}G[^^>����LY�1)��CB��x������W�Gj�(�ITG��p<\��J8�W���(S�R8�+����m#?7%�}(񮂨�$}�Z�Z.'+�������.��*0*���ሖ�;)�GD�z._�ԅ�C�;


s���⧧��p�M�A!��c��Ӂi���W��� 7~R������I��08��������Hݛ �0 u�D�.���,�����9���kr��J��t��g�~!1��Y�� ��u�H&�z�	������F�����ƹ?����I���˻҆eY���b�g����(���]\b�Р�خ���T�-�18����QSS��s{�7u�|���m��HDBA�C�A�@Y8�Z�Z���_�{(t�����ݎGi=ꧩ,�BB���g�<��L���l����m~ ד���.�����A%��s�O��^*�M�?�S�9�U��r�m��h��iQ�y1��i�p �Sp쭲6U�񵫻�����@�^�	I�;�\�~>�� ���~�,���,+1<H�����RiU�I�Dg9ݤh����d>٥U��6!*J��_G��9���'��^|\Ԗ.8$,�U�au}����B������?y���m�L|$���� 2�� ���:_N+�\=s�z��(ߚ|QQ�j.J��O"�r����C����K7�t/9g�pA��ӭn���oV���5��N?Lѽ�t?[ϣ�ap&����6�I��^��^�u��WUeU�t%��ߠ�,��i��؂�y�j�J`�R�"WxA�� �T>]���Њ��N�J�z�R��Ċ�`&"�Vw�m=_$u��x�m��|���ʎ� �*�Y����6>!!�+'�����׹�^�:�d�v�k��ʏbi7�7���B4��[��?-ō�1�&d��j��D�V�f5L�6�	�Be}�+.��U��4rUD�V`///tR~�tj9_��i�9*P�;���E�0q�UP�fBP\Լ9��-� ��*)1��;|�N�������������;01�+���f?�B����{-�*`�k�Z��o�~�絯��1Ќ�]P��jjW�7�o�����CӦ�7�����$�)���ȧ�8����j������~��17�y�x���ڧ[�o�c7E���WBIZȤ8��^��F^��=B}�˃KUU���n;���(�Ș�򱲵���Ѫ�!װ�xP�s�;����h\4�,��ie[G�*��]�Y���{�@R!w�2��Z0Νf-4F����	C����
���xI+�E#o4��@Y����`U� ��`~���끊��vԵSl#��7K*����(j��|���dZ�nxl���a{�����߾��RlPõ�/�
�!k\b��F��M���Q
/��j�I��B�R�ѱ8� ���Mc��mw�oz���ƚ�w��f�vi�%�k#�)�jΗ�Y��f���������2RIap����77��2��A�e"LLǥ9992J��1KO'��8�����B���:�v��������\�� 
of.m�W���gWr���O��~D�b�����O*����4���4-*K�ˍE�.�a�pd�!!�u斖usss�݁7'�E�ЊE�&�)��0��������Pv��4�ǳMC�55�&~������r�)���pQ3�`�a�&�b��a6�����'U"�.T@��J��K�}�� �A�������*_������%;**JF�-��?Ư�꧖�	�0YŇ�����)���[��M�렮x��cce  x�d�������EyU��*����������-�/JjB-[S� ���xD��n�xЄ� ���B���_(��O��PZ\|�'�/������	��k�� TW"h��f��ލ本��b;�.a��QK�}��iPz���5(������x����6�lJr��:����"Y�|K���q�o�P�kP�<��/����.�G;�����^ۏ��|K������0�!",�݂f���O��,�fH��HN�!I��#���_*=͖�f���1�ɲ!0�l�+�s�S4�9�V�L �J�0@M^Ǒ�D�Ǿ�����H|���7vk���N�|��Am�  �$��)`�2���c�8��*F׍@�|t�nk8�m�>d�>Q؛���'ȁ/f`HN�����$�a��M2�ٹ\������`Ow~<Kz��ED�5�Q!Гa�o��)͢�K�#G3�a2|}һ(T�EXb�;���!�4�@�Jv�9�t�,ua4��� 7�#���3�i��/Z˥�p��V�=�A��R�\�gD�'$�à�D�� vŨ���>�K��(4P���Y�H{�S�&��S'd�Kq~.�X�<993c����Ο�Bh�V����2y74��ƅ�������("�F���U����+�P�����[�͕�(�*�H���M5����0��*��e�L����9���X�H�.1� oi��o$}��AE@�R��4�X�� ��FHb) ą1+��AD��5�`�k[�i�ec�{Λ!I��:� [���,-i���"�˿�>��ҢZ9��P+3 ��􋞅����;��2����t�����MZg����.��`��ǫ?b	�3�c��gz��1�+#����s�$u��X&��;K�z�e)�Űk����?��jQV�⧘œ���}��Af6��	�Յ\�� #�d�������&�|�����/.~��l~w���-�l�(�N�{���8Z-��پ��]����I���DG���7�7�}�����A���Yx���G�'=2	&ژ�q�GǨ�g�����%ɳ���=�H��Q�u�B�1Y�߹/�sѱ���<��ufVP ��<� ��_$㰾>o?��0.����2�'&��/Cɾ ���W��o��V�.|V�k�6̖�sB�#>n����V-D�G���R�;.ewE��>y������2�a����e��rٚf� �p	E�+҃堔�)G���A&E�+ �'Km�����Ir�	�u(��[LOQek.�d������.U�d-��P�9� �fwAb��{��	0�Ǡ0;�+ ��[q��N�_���A�Ӓ�J1H�73P'��5�a��=��z���s�B����P�U5�G��AY3�0�,�+$�#BZo䠯��3#j?4��|gqu�H[�Κ�@�=��W弤�M�����N)j�)qWW�/
��mn(A:To��`sz�mv���.)���zm��ii��J��Y�-����"e(�(�hуV��r�CJB5�����׳�]ҩ~qG�\�� OgMߝ;vq�㛙*� ���t(�fU��"c���l�iѻ!�*.��>��Y�s�0rc-�Ň�-�� �W
'&����h�8��Pw%��Ц��͙%���׊�9a��gVU�jj}6�H,l ]�����~��/$�$�|m�ɝX�H�2�FU��hè�H[��m�W���0�������_<ckDԘ���5�8����d���{5C����1�����]\m��~����G��`aL�"O��{O��M��v���:i�ͮ�J|I�y~��-�������3䞽˽��MQ��锉�-�-�Tu�b���L�,=��#$��k����Wj���55��;d�Kl�q�:\{�B�n��|�y����=#S�'񳈀�i�y��^a���������M��'���ѩ*==/�m?m���c�9PUj�ß��}��TX�
`����E*(��$&&Uam��d|���y��Q�0$��		���d��d���<�~�&��(2@[u���߫ˬ0���՜#^�OyeZ�YW�����`}�|��U�ߕ/�9D,ZQ����8M8K%@��^�m����)+���a �2t|M�*BL��/iRoia��$���x�~j�k
M?ԡ�6oM��U-0��Ty\o6�-���M̉��$�Yt�����;��84|�N��k*^�H�l�mr�qD/�J��tr�x�tE"��7̆��A�~�qsC�XQ�~9C�)�N��V6!�׎�U^�U﮷�R�<�)��
�!�����p>�b�Q�p�v`L��T�������D�z��-Q$�0�����x
ӧ9ϝe�~�l9N�~��k�|ƻ����t�8�c/!��������/���2�<��1JhKP�����P�y�_GeG�B�����k������r���g�\;���+܅䜻{���®BX�9��<?��^ў8���� =55���ׇ�������z��ń-���H���3N�҇U�b{�Uo[�w�C[0+��	E��`Pw{���7�.3�9�NpC�V̈������C-��{�w��	{��^D�-o�1�	�❵/���O���A���wu���/�Vˁc�i��l\|tt2�Ǎ�]� Q� �;��Hu۞�8��]MMM�sS3E�(F�-���4�� "O����f2�_�=�D�[��x�`�I��T�a펔]�Q��/�=�����Z�p�Z5���55�ۮL�!���u�aU>j���4����wvd�V���抝�U� R�5߃j�_� �{�U�:�����E�g�M;�s�F1r���[;��,�य़b��<}��}���W���1��O���;�i��NF�r�����8ȗ�L}�)��iio�x�]�C�L�����ԁH5��,3B6����l^a��P�:*5^��Hئ�����z�םL"aody&�ļM24r�r���mgc?f�C�8��؟�&�:0-,�M������_#D����a)�!��� �$���=.+ڂo�G�5ESjǦӯ0X;�߹w�Mt�Y�܁}�m*��M�	Dۈ��0(zS��6_�o1ɢ-�{��]m7n>`R@�<= Sսw��[�r�M;�ӿF
||>��
��JK���?��u��]A�nm~�5� �{�V�j���W���5�7O]n6�D����|��C��?܁r��������Nl6;`:�M�M齞��ĶZ�%�i2l7�l/�^��Q�'T��a���[����|>]38ش{��d���Z�l]�ۨ���2d�"?��ɔ^��7?�7|V?&l ��b�:VGr�n���;�w��gC����,S�[�L�C�d�2,t_��,*bb�V�RKH^�N�H�;��4�����i�'�"�&��oI'|s=���l���W�/�( g�k�]��@�o��9��5;Þ��%0�6[�\���Y=��W��^S��<__���x�1�z>';���ᱦ�z�҄�⥊f��،�X9t�������s���]o�|XN)��=ԅ���vf���O�����:r�*ʑs�Ͻ��$���L��P�n�ylww�Ϸ;���	D�)O��7��^�J^Ab�3�����%��D��y�|����e:��>Q�-h�-�l�q���C�l�pm��jyp�N~f7����t��w
~w]�p1�u�C5�D����){	qSF��Ow�Y�ND=���'��;�\b��3>û3���H�sc[�{W�0�v������8�j?��i�+�C0��Ceid������a;>:�ru�ګ���c�VG��J����9Q��po���o�)I9ɑS���3���z\ɔ�ma}���@]BKj�??"��옕P�c�����x��MY���oLe-�#������NW��r��D�$.�9�A~��
�܉�`Qhm��\�+�F>6��f��w���ʻ��n�hB�A�����W��P~N�_ٱ`u{U�-�ނxq,}�H��#�Z�!�����1�1�ȍ/Y �DB�*c��ް�Xpn��z%��{���!���' ��_h��l}Ѳg�B��'��U)�vJ4p��]�GW �Kg^����J�;�S�j�����;���,Ղҷ���ӏ��N����M4(�R�BIUCR���a*+y���>Fl�|)'����d��J�W��נg�_�π�E�����Gն�Bp���<+��Z�E>����� �x����B� �5Ge���Z5v�Q%��6�Aa�x}��'mr���s;�LH���������ͩP�;�Y���3�B����{5,B�k��DNrv�e^dK{Ks�^�>��%�	���cQ,�;**�����Y @2?��H��,�,9j-#�Ў9�-�|���p�2�a�kƪ�3k�*ɅI�Y�q�t����{l�n|R�/�B�. �	a�!��\����湻�S��{��0�T�w�����q����Q�������tU������}�E��7�m��B1�
���� �]��W�q��<�Q]��-��U��M�:�%����jf
�l�bț$���i���}1��§T )��)��a�㾌�O|���i��U�_0L���#L2�H@��$�H�X�,.��.7��"|��B�R���%k0{5�n\k�p�+C�Rji�ag�2E5�N�ģp���*_ئq%����@����$��`�����UJ��V�5*�C�E���x��K F)��J�?�!��{�p���G�+a��&Ҍ2X4���������gJ�^Ӷ,�_ʂ[y[\dL}<�F�-��o� ��Z���a�H�������7�6�*�@=�,~7� )�N�[������a�857�_]���y!Ic�y��â��?��He����ht ���o�*ЩC��#� m�7/�O#l	��P��,v�'��<�b�n�v�zKR�̂��*���ppr]of2�ʭ'����2VV���3�qvz.��G@�P.�N�C+��1�eB6�ϴ�l��8S\|:Q�Iha⍂���b�)����m�|�H/�41�?HA������������kmd
��4j��#TB��,߽Y�D}�`K8�w*kiL�2�jR� ++����PՕ�#�B��3p�������h��	�����Û�	��Ҋ<%q�ПB�^ȃ�bJ��o����*���GZ4���K�e�B��u�.Ɨv���Z?�h������]�BL��#�E��7H�B�����/������3�@�������t5�q�y���D)��'�1&Ü\��v�&T �wA=%)+y� �/�/=3���.��U�VH�lh���L�Z2]5;�N�ڻ���EJJ
�W���}|��P7P|>99)��s!+4���"���F ��%\��#� C�/�[����>�0��V��o3s��7��y9F�3�X�$fIPP*���p��N3tˠ"�vDO��j���p5u���)����>9Y��}2J��>VW>P:x�]�ܻ���;X"��p�>�h��1DWQn���˃��[8'��<������3�Z�k=g�v�u!��D������Ϣ�=�T�,���6��2�l���$t�?��Y�
/���;�-���=� �p�g_�F�{z&pj��Q	o��uJk���d<�,���w����ߩ	���	��=�!�s�k>s/��@�����>�c�Ç��E
��h���rsO��ܒ1#Q�/�BCW^���b,�jjk���C��ѠU������ȣ���� T���Tzs��[<(�Z�d $�x��(e��eddD�o����mm�;Y��gb	1at4�$��X��>���������i���5%�r����I��=6,��t�Sar@�m��l}��Sa.�R ��~L�da��;V����)��@�"m����./�O1�W��u���)x����ɝ����Fb"=xZ����ǁ�UB�;��V��Г߲��
<�k�V�ų����ea2���Dt�,���cgyb߬x�z��[��[�Y��;XJZA<Z���#S+V���w�_�ܧțM��У�e� R?�(�f��͡"� z ��n/�?�[ħD�G�(��KZ0��Ng�gb�~Ա��r)����(�᩸��"����r�Gdd�ک�gF0nfj�T�������8���G,�#��&���̫9���υ�ZO��z���x3&�X�{�DH���
;CtT�}p�8sS8��Z[
��}�1�	���8h%hG�a�@�}bEN�8[i�sZ-�}<�/�)~*|���;_���V�9K�Զ��Ԝ�Y��sWM�Q�o�������%�d"2&!D��x�G��ko���;�u'"S��s,-��sVRw���d����q$�=8,���wU���o�-fj��f����Rh��/��j�_w���{=p��B�喎'����(�I�d��t�W���?��no�t���^���w���)��6�Jz�������w�G��gf���kϿ�S2�����H7��hx�*pF���:�Y5$b�h�6
V��jR)αzh��f����(���LJ��O��I��qT�fc���.a �9�C����&۩uL�ܢ�����*|ܞU:�"�gb�����h�y��=���*�~���
�w��a�u�w���8��F��cX�,N��s	95��+�g��v5�O�h�H�x�l!���Ei�A�o�)�s"��h�=���w�g�P���ו�zB{���w;33���N�0Q�Ԍ%��ģ���׻��1I������/�}k8��h��D��O�kȫ#��>����|:��D��)ѭn%��>�?��1���g�yf�Wp[���Jh�I�f�������A>�m1�d�bu4ؼ�kb��n���7Y#/9��*��c�	;骃>��1]����p�'I�	�H,�0���,�-�gy�\�V$ǧUؓ�~�e7�H�q�ח���}coKZk�?N�����H�l�w9�R���@Q�I�w#t�B�v���v�i����`o|S3N(j����P�~F$�L]u|��s�8L��#�Q�����"��A&�5Hl���s��6A'� ��Q0��v����
�+�եe�m�874@tA�V]����9��1S�0!}��ނ\��T�Fb1��L�]���[�̻6���ڠ�m-�:OD�m 6;{i ۝�� ���)�a�|OM� �!�k���t �)�t����U�Z�<�_�4�qg���js��t��0�=�&,=��@	#����,]їHwEݍ�ͳ����:��%%%�{*�nv�~x����>�U-[/�)�����C�{���zǟ�wJ.KS�*��_6x�N�Y��[�Dܞ�)��Kz�g�:\�����G���K���Vf�;(�m��}�Q53�kt^'v�D10_k2����5���遯��L�	�+DF�&�1�>h���؋R�eQR��Ofu��w��q��e�`eee[�-�7I����:ji���̍	�J9�4�8�I�@��,�`ӝ\+`�JҊ�D�v� aXa�Ԏ9f{��qf���|餛/�c�c=��6���ri��w{u�xq��z4���t0t������z�u_"#:�8!~�s�h����r9E��eQ�!j��Vx�.�E2s����"����B�T�H�	eE:[W5�SFh8'�4��s|_�䔲L�Pg�]�_Z�2;�˕Up��Z�#š����`2���
����W�#{>�c�[ѱ� _�|��״��2�$jw�[�8_����K-#�c��5����`e�ϥE!�l�>������B�M�s�+Ӏ��w�3�l1w��)��m&&����+�{D�4T��*�?�/��-k�o�SS~�e���x#����y�C��;Ѓ5W�IP�� �{:��t]��P]��/��������_���D�_�&O.�rL}0X��E�R�ް����h�T�����(���T$��mt���o�,Tj,u=��c	_a+牄�C�ZQ�hWb����ɍ5~�p�ì��8��|�u���f,>?����M�tO��/z8�}������]�Qx�v����5���1�3%ft�zU�~.k�����	�H���tK|���I���y�I�X�0�mu�gV|���ێ�u1_�:����zs�[7E4&��r+k��	�\pA�&�N(����imm��ҖC#���6vc��\b���T�|i7?��^�3��d���{�(�����u�Y���0>��%?��f�C��ݠB@©P?��E��^��k���,�p�������Ս�����K��<��2a��1����h/Z��6�׿���sߏ><�s��I?��'��'��\P�%�oS�몛��V�l��b5�w�QTD����k�O.Dh�%V�#RqS��#P���7f�$G�~fձ����KNЄ�3GE���v�@l��AR�4�;Q�s"9�]x�p�*�P�{΋z�̕��s�"�L��e����J��P��skӜ�^�ߨ�Z��O>���I���oV�z�
��W�F|�1�Y���⥴�8p�62>�3>�g+����
͗`�v��]x�&v�[��:J��|����p/G���&e��W�_��RP�@�h��6v����-�FA�pdZo͓V��P������N����
(i%����0ǑpD`��5��;�1��ji~#,�Y�#�uEG�"C��
b:�5��cs�Y@�ߠt�x�J�@�݊y�k��+�;���e�B�w�z��i����է��
��|�ڏ���Y�
z~~�1]�ҎfV�A���
��5222���}��Ӆ�$�I�'�ˍim��<�:�]�+jkz��L���9雽�w�ޓ��A�q��b$�K�z�ǰ�j��D�����!���T�Rߔj�d�'�����rKV)Rd�{�cjAo�,�1�!�:p뜢����y�^�}��b&/�xB@��v<8�"��td�s�y/*��{���w�gɏ�L9�_���T?�GW�R��%7�=*���/p�\Ѝh_������Y;X��?�R~+Z���g��t�.3��{�ҷ��[[Wg�FQRi4��E�tS#4�әju�g��}\�k?j�j�ǹ���}��-���p"d�l�<�L����)�$�SLӎg���'N;�6ur�\����|�D���h�7C��>�<=�?e�q2�dGf1h[����R"5�����Q�h��L����(�;�t��=h\#�E����r�X����I��,+�n<���o��G�i���l��\gC[�Ρz�F�{$���l���.��4��8�53H���Rd�X�Qä́Ih�e������+��!#W���k���;����O��$��<��y`!�}��Ġݞ��2{���K/��q���Q���_Ui���JC�'G��8�K�P�����ˏ۷��pYj�|�̢> �M�K2��/��ؽ���s�on�_�K����?TT5��9M ��O�qT��dzo�w���V	�p�QԖ��1>���K>{�������|�
7�gRVr�����������w�1������%��
I��s1m�+K���0o)��E8�V�lE�a��P��8v�K;���	wg$�ZEq��-:��Z����μ�Rۻ��e���i2QI>�f4W\C���E��>T�D�����w��	��ƃ|�+�Dң�
��H��}���Ŕ���� uo P��2U��?Q�:���+4#�t��D�T��n��?�����R�����?u���pޛDK[��_�A�C�oJ��ss���g�����
=�7��� X�;������ð�sӻiϏ���u�<�1�QUz�hh~ux6�ө��`���Dxt�ħ�p
sk8HL�@Cœ��X��1��4��C0�\�<�Bnã* �3'J��M��-��ۢ/{��(��!?�k���x�`E�W��������u_�>�������tt��ƕ������.�?Hp]�"�;3�<���S�wV�v�2]x�yY�53��a��=�:�c�bt��ǚ�'�	�������>�JtG�-=��?�Ń�H�i:f�3~�d���m�R�:����}��jW+b�f�&��%���`Ag�Dr?4��u8ڦ�szk�i{ػ����^�q�N>\�,�z)��|j�`2ǔZ�D=Z���D/��,F��e�*�;u�eW��,���q��5�4�H�^2iW���7�D����lo�R�2r8|�ܶ+�6׸�@Y ����=���M��0,88�>܄�^`�Y����-��4���1�����&�L��x����2>��vV_�1�յ��c�Q1�$�qrU�n***Ɩ�k��3�u��xy	���W��ox��7��c�Kj�Y3E�/$:}}�z݀�:PPP�B�N��hA�NB�;�V�pӻ�O�*qi`���Q��̟1Q�3�a@xc�B�A��0R)��s�l�jdݟ*�-=�z$)nnI�(W�fe ��RS�}��o�[��>@0-�,��.�&���1��3���s��r#^?'�Z4$x�8����8 ��ך�|((����-$i_/�m��C��yE��f��O뛌�0�?q����#��F�}�d|��r#��}S;��9�\5b�(����A� ��bKWb��E�4������Z��ޡ���t���By�vB���v������">W�]	)�1aX�Yl �%�]Z!(������ ���y�V���\}� |v���+�j�5��%�������3H�]���Qt�eX���Lq��Wh������J�k�����K�隝;<����^�J��57�.���m9PAR�!@n��L%p�����������&4�[�������]F� �W�Bys��T���Ȑ��KBD� s�F��1v]�	�f�2��Ĉ"�ir�a/8_�*������>3vb���?rY��6��`yG��4L��c���)r	�"�Dn�ԂܼRΦ�gH�	��<F^��O�{6O~Ⱥ����=�'�	$��=j�oyg"���BpH[�\��,Ғb��7�{)�LM��n�	V����B~�B6�W��4���)������e�zD�_����K���(���(��<[*b��90�]�,ֹ(���J��TT�w�.j��n�6�T\^�~��@�d��w�L�B�կYۗ#���ܻ�����ܫ��WQ ��Ë"��*�����" �2o��\u�3����0��zG�ez�.ɝ7�V]}q*��YH�	q���p����
�n
g�g���[�A�u.w�4F�b	��:ьٕ��d�7�;YA��:ԭkkk��-|�Ց{�p���<���Q�q��.���#B�����JI���<�]�対��&���b�rnl�D��H%��|/	#㔚��Q�r�"�lN�bi1guRE��YUlaAA������L2��=:T�����c���C��w>P �J�6��,����~#J�MRZ�":l:��I�,i�oן/&��H[,�0���BB���~�.�r���,ċ[�]gS�]�d>??0"W��B�:-�{��x]TT�E�sC>R���t�Β]!O�n#R�f#����-��y�\��e���7>�����8
�`4�*5�V��Ϫ�ҹ_�_>g�v�� ؕ\V����g��NWʕ��S|��=^I줚����j�:\a�u907]����SSלX�?a��%�긣��,v:Y�x�� �g��O:����
�F�h|���H���oX<O�f��))�T�`� ��z�:��Tq���t}k�qa�"��cJG[�1P�0;���������GW+��صj]�aHf���l��õ3^+{��q��r���m��"��0�,N����ʳUW#�&	 ����%�?�$)5�gΜc�*���5��ۇ(Dj�"@���m�Q�S��ɵ���)?�A��	��LV\�.���\��p����.��r���P^uA��4^F"$������q�4P^�'�U?%��6��Y�q����7~��8��>?�)������fd!1!����bAV+oG*��K�Т���� h�i����D��{&�ؾ�HP�j|�<� 7P���4�\e���ں���:v����Ȉ�~
�)���\Yn�?Q�#"uG���_�0�*�^���fhǹ����á�OJ�|nj� ��H���Nn|�!���Z^��5�6~�h�����&�������̯y�͖Ji&D�J�V�ﻖU*��)h����J��@�ɧ����1w�
V�5�Yh�������/uQVVs{ŭf���N&>�3	!�4�b��m�����t΄����x�>߾o(++�*]��C�T����R�!��(Nf40`T�|w>s��	WY�ah���Vq`]��P=�2���=!�t�4�`lu
i����s˴�&��}>�V�����3i���Fnx
_!�Z=9�@:6?TD��I�g�6s�V�����=m����1#�G��rED�~�����|;E&Ąh����p`R|��7b���a������v�T-pyLƀ���sX�>�72����� �Q&�[����mK�禧��r���$�F��2f���v� ������"�( Uk92Jy���)�ۏwuR�R�G����"ʛ =�ts'��g�W{�?�~�N�O�)Ƃ�Y&�-~o�J�����@ҲCG�Ҋ�*�2y֊�Y�ŋ�:_)�ߤ�Ē��Br�V�=���E��#>�8�|PT͍w̸8n�*�-]x��G�q�`�P;��q#�N���jk�{v�����A��ÈqC#�T������F��ܽ�c5:^��4�eh>�#������5z���N����ׇ*��y�t�r jK����k�B����`W��M�n��?SѺ�}�O{��T<�q����M�^W�u��>�m�v��Ic�'�m�������649���~������k�1֞k��|������
�ѫ����m����@��_j+�/fg-�x�����m�Cñ�Z9rz����0�|>�A< 7x��џ��p��0�)�R��pf�ѕ�:X���i�9��I�f� ς(z�̤ gb�5FFF�������C �Z�o	S9������s�8<x�p<�"�Cx/����յ^��c5�ˉ�۸��}��X�B�-���=�ף�S�$36��<� H.dbWV��3�4m-�\抢"c͒KP�_Q�d߰�gH��i'��p�!���joX���В>f.ޘ����b�讴�?q���0��Y���C2�8p{w�Ñ�}�)3�̹t����0�۸�^ͼo�ǋ�u�=L������"Y��!��@s��~�_Q�>'|BX���e�	�P=h���=? E:�&��B.�rEj:=")�93X�xF��º���:/�`*��02�o
Z֋�C��=zd^�^쁥�������@����_���#�L؝� i� ŀG��̂��V'Je�ABիߢ���2F��.��+EfS�h;+�|�W��aX�<kTE�?����w�v;(Lմ �hH�-�������Ie�W.MY\6�����ʅV�"����@��_o4�9�����cV��ӿ���`w��ޑH�Y�?v�W>, Zz�^�[��n�8 �Ei�[.��x���@Q�7a���Ի>����#C���0=�	�������E\���I:�S��(�g�fem-��h�p�����[�b��*JC}�ZE� [���"��3|<W����!O\!��0���®8�w��DJQOf�����L��W��Y>�WhS"��p�t�JDJs� �z���J����o׊8�L�'ֶ�׍�.�U���N��4�����s|���e�	@�E����O ]�����z)�!��	��FOo��w�Kn���f�l�]����"����K�j�I�.�2�ōs�n0��<8��lu6<��y:*�V���M�X.�n��a7G�-�,E���Ti��v��ǫ-�-�^݆Z$�ozf:eYN�t*P�Q!�#N�l�'�Y
��G�s}����&��t��R�"c�H��p[ω˗�~�l??�Ie�v��ԫ4z> �:Lմv�z��b&�=��q`�<�ov�TL/b1��?˻;]F�v�����.���R���݌%bR���듊�J#��sg��<���p��;���|4s�\�˱?Y/}����7�l7�l^3�|�@�"�-!��ݾ�7>P���iJ~j�\R���@I�nn��f�ci~J3
[�_� ,��S��LAA�UZ{B���1���\�H��j�p(ZI����CA@ak���w"XT���sX�*��>�Z8�yW�= ��l�[mp�����h��C�D	8Q�m��4���}0�j��d�Qמ�ZW�w3�|�,K{��oq�"���-�6MMs傄�8d/�V>�s�ba�A�Й�����QX�Z�",�O���j�,Q-jG|���W�[��[���@)=�t;�S׎�ŝ2�)���Y4]��ƙ��������'��5�����vp V�%�R�:���5������N���؉�f!�Q�=.�?.�@7LL�}�;����\|P*���OzP���v�i���e(<�s<�í���[]�h���I���	��@��qQ���}�Nlm������R_�o��ԝ��&M�4��]I�5^�����6:6��ˣ��G�eydR�7_Ծ�ܢ�d^�f��p��T��դ�n���� �����v$car��l�#�-��ܕ3l����ؽ�����dml�Eޏչ��٨�8-�F����ij��Б�SZ��xȁ���\/~����+��@��҅,�h}�c�����  �8�KM`��I��˧�s���%�Z�͇��>�����JtR5�K���tz^��C���/YQ�x���g��Զ
p��5< ��+��h�[OxE��ĭ�I�l�$�2��4��������Jj�v���;b*\���qB�r�X.s�A��O��� -]�H~xڣ�wf&�<���h��Ϣ�94%�GGG��ͣ�2��pH��Lqo�4J8�V�$�b&�����u���6G<s��M�ʆ��S�
������6����v�J��(�</�@�)�0�R�{d��iZKƿ�7Ƕo�<�������.��@X)�a_��,�um���� ��5ĵ��JZ߸�׳~�<��s�����Y<6�/-��@|�������3�e�$5���`�f�E�,>�r���Ux|d��&hmw�3TZ�XE��=�Z����/���(�񳥣�S���F�C?b��'�r�r�m�i ���e�p�0��aIV0V�K?���4[�.0�nbJ�Z܂�qONl�w=s�߄�yB=���ƨ'�,��� Knom&���l��� X���Ĳ>�ԴT�m4,J�G�������0Df�p9�f��!� h$��9�'P�kރհk���g��������@5�#?�8X��k���/]s.�V���U�ԋ�D���LU��M�6�0l��4��%���Q\Z�s'5(�Z�l���'8e��㕆s��
#�;��x�?�=��'�f	p���
ѡa�����ȯ��V
�����d&����n;����J��lB��d}dCA��:���D(�)8�xm!eC�Я4����_]"��t\��W�0�N�'��J#�@X\��y�k����߾an��z�>���(}Q~�-)�������(�T����r�7����H[ŭ��)�+�+����>Oc�~f���ؗ��T�E�QFKAI�_�0n}��r�;��+$��xB���lN%y?��L��� ����@�YA������x����k�Ztβ�Y"�3ԌZB����C\��'B��j��8���gr���o_`ɿk��#(!��_�?.�?��f��{t0�-,V;<C�za�.?1�y<Q�ʱ��T!�B��6�'$E|(u�*�V�%R�:�	�/��YXY�b�
�@�%��g\�i榽v8>� �&�*�MӚ'.�F(�=��`��P,�N�*k6n�ǚy�
+��K���{�{��?�<s�r�P�P��Z��(v�U[[ku}�k1V4��b���H+*N�F<Í ���5<ӻ$�B�
��L.��
V�06�+��@+���R/��b�a)�c�X�a����Wi�=�v�+T��11B�C�n�V>j��u�Eʬ����47c�/8��Q�������]ɷb�KSa�&�ø����QMx�yKEqG�g�Ț7��].:1O01x�=��s�H�W~f�f�
��ri��N���A�܇#ኤ�є��P[_���
��(T?Sm�:�_A��w�&q��d˦ޛW6��a�o#�Vs�%PFvH��b��{�syL���W�"�C�Kp��Y�O����%��O��N� �����#C�X��kN�v��j�0���������5�s)�2�a�C��ƙr�:C����_N_�.hHs�δ&�J	���d5���M���5�&�ﾵGhPl��~� �2aA�#�CF���Y�t.f|��S-=g4t`Q�H�M�oľ�$L]�/�-���3J!@��z�c���}8w��>�6�N�ZvQ9?��'��O����0�ؐ��@����ҋ�{*��e�P����O�y��f���$g����A��H�x'N�O�B)Ou��������f�[:t�p!]{��9� Us=�D�4��������"�����|c�wl-o�!�r�Ն\$��K�����)ɑ>�+���"�ȇ�x�ڿ>�wQ�P�8��BsY�w0�����|tTBs?i���&?�܂��&���j��N���V1��:ll�>�c.��ڷ(�#."��;����5�Qxf|��N��r�4��
��Z��,��K��lmm=�T�y�	E�@��\u���2��l\
uV6P
aXϦ5HG9.Oof��_�^y���'\Y]/ޝ�z�		"�+�SN<�k���S=ص���g���W��ZN��rrpH�u�w6��S%K��܄|���
���O�tl�$�J�eK�|�8�9
���|�ȓ5g��X����� �8"hIXd1�&D'y������Bx��ϛ/ʅ��¿|haH4�-��	�9�7��J
F�t3�k]��AXe����K6A�_�"�j�DL��Sq�HA;�;r��K�<Q�\폚M��ǫ=j5��DLқ+���M}�0�A�6U``��5v��-�����C��P`@t����i�61��4��V�U�e�x�T6^�A��T��c�������hK�����!�vK7� �x�]T]����f����M�HP�H��"�L����o����C�����D}�ڊ[`�	�ґ���*�������&4J�(�Q�w�5Vϒ�}h�x�`���8��\���y.�?Y������-_�_�>�|���X���JJz�g� ���	U��:�f�Ȋ}re�59� ¦j� ����Ȼ�;�(;�+��VB�!��8��օ�2�6�.]C��k��`��k29..�?�K4�o�H`0��՚�\KfFF�����rb��q����$7š_��g��P�5��O'P�=�䴍,�|��9ȅ]YQY	_8=�<HK���M$�c;�R.��U�ԟ0J�������SU]�laӡ���1R��Î��2�}��F2�ļ�.�}��`��?��'s�)�T'�p��R�Ԕf�����Q��.�`��Q�`2.�������-���pTT���1ȏ��&���IjD��'4�O�4Uĥ�7�~Y�ӂ���ff3F��i���K>!�F17�{��kr�Uy�D�.��f�;B[���[�5�u2�^OSp���0}�1�|IK
<�C_�҉{+�|n��p\�8���$[�J��5����h=�j�rH�O�c'xj^	���1�;�^y�$1���@�4^'/��`�G�X�O��C����� A�'C����	�#�:���-�z���B�<D]���X/-�w��+�Q���)kS鵝�%��$̥�C�����F/�����
�6^9�^����a4tf�:Hd�Yg��0ˌ�al���:G�R�1�X&��ɏ��إ����?��7��VV��٬�f�]�W���aݹ"T:�Sc �8��{��L0������V�+��UB�-�����qds��`(�<e������du��;��_�PI�2�yL�'�͉~�-銯�5���ͰA�_}p,�7e~>:{�g�����i��u�ȑ��u��BJ��~9�R�$H�7��K&�@������c���1{n����7�Y*B�wSZ��_�Ԓ��L����:����e2�������i)( o�3G�ڑW�&c�o�5Xҋ��@�Xju�Z�k�>�b+�0�֨�D3)U���>w�3j���c,<VP��k���[Ђ\^ ��gR��3�a�b��\��"Ѹ"��޵��kD�ħO������l#�����z�_??F�g1�p�\��@��/��=�ń���#&�fW������=����K�JN���Fg�	�^q��D�na�4:�˸��a�Nw����E��o�'����͇{��,%5^,0��%�%(�<*{������>_�O1I5X��w9c��
A��{�\fSA'x��,E tM$�_D����O�ȋ��bL�*�8asY�Wg�RE`���dq� v���L�d8%-����=@|'Ȩ��ΎR���5��x���Mk2+z�?v�W�db5�J��X-�M4�ɠ�[����{Ƃn�?�u��]�l���|�ͧΠ�()ub�`�{���c`���k�����Q*�M��L]� �|O�.I�3�<��6�V����%��8�(ֻ�����t�V4���񒉛��>Nq���4�4UT������b��M�gf�������w��1Be�����HF���2˦͕�Ef�z�$��U| 
m#�[�\�zI��/->�ޯH�*t�}f���t4{�;�f~��D7dx1�����8P������P���ɔ��q�_Ή6��)+�d3��eݳ��ǿĊ>�r�m�T�ɬ�$��j7ۅ�z���j2�;h����@C��Nc��5w�pa��f}[�J�Fpp��������*{o|�k���h<F�u{-�76Z��HB��<�=�����!�� Y��ly�%��|�i] �e;"�o\��am��4�q>�uǆ�m}>��\6YT�.P����3�u��K�u-��j���f۸ϓ��97�m�1Κ�
>K��}<���5�y�8E��u"GG+o~0��%Ņl��e������g{�oGʋz�'
��\O�<w��+��݉��1���3�*������yb.����$�t�k�_���>��d�8���X�! ��Ylx?E�~�O�����9��A2U�F�.K�r�H|�� ^�h5��ǋ$�F��*�8������P��������:R���f16����So��Q��xŝ7����w��wuǘJ5�HGy$;��=hNt@�|ξMmst��j��J~-�%�6������3�S��	�5ӹtY��h`kb~4�a�O!�<�<7�M�k�Ö/k�� v
�7��^2����z���PI�"aR5)3V�r��#ɅNT=��< '���o���:�BK�?���l��U���޷�m?���6����|`aUZ�O��P������b@�<����u���#kx�O6��?�rZL�=����#��U(gǙ�&���F%&J'�̐��)!� I�ꅗO���4Y�6#ML8�;�7ȋܠ���f#O�D�j�.+�p��������~�)�:�jv�P��^״�B�����ycR��?ܫ8��W����O�
�?�Ih�	��"~������X\/�^a�3�\
�l����]p�M�Hlh��_�����¤4�EW���;�6��<�Cz�ta��	Sr<���w�������J$H���w'+m��C2R� �(��7fh.�^�ķo�������D"^��������X��^��lh�e�O\e2P���OM�/�z�m�!+i��+��/�C��˹�P�x�6���:��_;վe����*	ÒW�ЊQ����@�o=ң���gE����3�ы��r�����XiȧH��P�>�g$����G�����2��%��i�ӿE�"�7��Wu+���@jF֔�h���3���f�?�5��-��\��l	cH�D�>p��g�g�֜a��Hv���;���?����xl�D%%�_��P�-�t�<!��6DBb]�_=ϣ�^�@��P>�U���P��HK���7�-�h$y
e�""��F���a�"A��AC���Gj�+�9[�W@���Ѯ��?��6:24d�P���O\[�'ňB�����O����,b�at�t�J��Z-gU����Hs�rI�����q���x^\fYK��e��K�r��ƒ��h��iw8�KS�b���x���8'S�S�ʦ��7 /(�J?�L��4k��>K��{����-�{�JXwmm��oV~i@@�r��~�|D%q!-���6E��U���T���m�oz�c^��t��n}Y�п���E�Z֛%�9C����Z[�D�>�`�n�`��v/�Y"������⒅�|_O�L��|6�QTRqe- ����J�z�=�K7�%����[�:�*d�0��6�¾���3Y���W��g��R0Ւ27;�O����G��:+J�[t ����AF������]� �D��(  ��!�u�G�*���΀W�[#�*�B)y�M^� >���cK-����k\��əj���9����Nə�{f��v�ŧ��zG/9_ !1���^9��mY���7���"'H{�e���F?�>�~S�t�f-8ɘcD��$q��hom�����}�(>_nx�G�F�UU�f���m����(R�����k���[*fjJ��[���U��l;:1a�Ga@L��5�k�n�i8X�R�����NȥL�t迾�ǒ��"E��O��G�l�7;=eumL�L]^u`��-��r�r�MY��gKض�]@8��lk �i���~�ZG��a4:n G���?U�M���q���o���0�h�9���A0==��J���K6���� w��sT��P���7bտ���U�I@[\�5rS��:錀�C=���,`��v�C�@�Ĭ,�3XF/9SgG(�2@��{S�d����X�n����nBj������t?�C�]�$L�N�͜$�ϊ:��}%��B�t@��?�k�v�)����7��X������~c~5=�����OF��PkF�1\o P�4}.u=��]�FU�[�0\���n*=��x�"�����T*δ(�=U\*pq_&8��Z��f��I9��omhԟX�}�\m��
��`5���b�����pR�%�=,H=O����M�Z���UCk.��3~�Ω����Պ�;l��j��/�:pQ�.���y�n���j�k�%p��&�ݺ��9SBVH�Db�b���iu���h",�Jvn/E_�H� ���u��+0�N���K��h�" G��g�RF��w��'���.�m�+�%'��-%t�5	�`퇸9o?ڕ��Q��8O����r2�P�=�0q�c�D�T��b����dA���G8�l>I�1=�n-���E75\�(=�MA�o����q\%`@��ё�rL�����xΏ�:����W�/�v�?QH_�y^��	�$c���z���S�����	�r��?t}W|�^�"_r�q�*X��h6�gQBR�g&x�c&��]I�z�B�ylו�R �qp�|�a���Y�	K�}�O3��~�@�ZݒOu����授`awe�<�a�l��7��ˏu
�ʬ�\�U�v<r�G�u&_ɮ�h�N���~ݔ4��+����*�T�E���G�8�?�q�1�Q�v�,�|�۱bŹ9�nj.0
qS��
P���>�.�bo�2�o|��VQ^�J%�igӬ[��u4�h�&#Ä�'?�Z���L��Aڣ�%+PvbO�����^.|{%e8�m���t!Wz�R�c�Y���[�;v9 �K��.$]D�ȁ�ՠ߆��`M�d�Yø)��2j�Έ����Y��]�~&�49ۦ:�h%������lg^V���%1��˗�Mo@\��).FKᐄB�l��R���mZ6Gh1U�ι�����J Ar���CHSPԚ�p�L�W{x�m䝐I��"�è�ϸ�(*�C++�d�p�}�X_��A�J<�eɵ�`&(�$�_g�����h��u⚊��� ��Ue#t��,���ްH�a�s�O^˹E!�����ɉ=��E�(�S�z��q��zL	Ȥ1����O<�� �NȾ�ИR��!c$����㎭TM"6"5#_6�G��gY�(�VJ*k��. �	&/94����#Q�Eyy����]T�]��;�9���(��m)^������P�lBi��_���C��4�|�Η�=���*@k^�C�8]z�*���	�p�+�\�dpQE�~Y\�A�4���bI�jR��ŝՁ��V�K�'=j翦y��M�Q2{���B�=�q`�!��F��Μ3�!8��?LC��7y]<�����r��q��fe��~5
>*x�Y���q�]�ܥeٵ�c��Hu���[�R��*�"��)b�o҈/��2K@��t(I���h���ŧ��
�r��"ǻmH7�@�H�qM�w��`H�5m8��
נ"���@�3J�/S�e���`Q�$A����G�����bx4P�w�Д7��[�������Q��O54{�+������j��ܦ4���zm�ʟ"dy�o1d�P0�A;�d.trVmcO.K)@+/�x�	��Ӂ�	6�+P�p�쯝�ŽK�����x|[���c۱� �.�-:0S1���S�<F��b$�s��H�s������,�^Z��8X����)���OD\.I��p�#����V[�5�6����˧#s?/?2k��X��QZ��L�	�:YQ#�m���#����B�����T���OTW�Ї��X;X6
*U��gs[>FQW1�����*����K�%ݏޗA�`�͉8m	��db�k�qE���B�NU�]pu���t�4Ɛ�g��gF��J8�Jb�
�� �~̃�ټ��3�3��)M�VV���i�@�|���S�~|M���7��"����=�P�#P����5�N+��0��ѵX�8�13s�W��-��w8�y#r�^�l�S�$)@����/P��.�F�@"��1�G�,�7�ʩE��B��RG��I�ʋNV��kt{^fq�X���(Sz?�<�������kY�������w�%R��f��K���ʶL�44�����]���O�I**�76�`�s-�&��JH�)�T� �r�tJ�♽�<�Ľ�~0�,����}jnNN�����K,���?�����Ê��
���ωDE*�VN���Ɯ��t��[1���F����i
.X�M�����!y���W-�t,5&'��_j[\�����S�=ަ��ߍ>0�����S/�2��h+��H�����<Q1�H!�Ȓ������~;W�b,*P���d�
w�Y!��l� ��M<�Mp�Pv1σ܊a`?)H�q���|��C�\=D�ɜ-E��'��{�;�I��0�tJ��ԗX����+!Hb���6'֯��f�u�鋏��a�/�%6-RB7.�����*8�3�#M��Ɣ�=A�~f�T��݌������df�|;5b�l�k��^����T~��$݅���񇐚�J+7�(]�{Ui�_wāH���%���v���0�X�A��T��h2�޲z%���0 �%����g"���Q�u��8��?���2~~��DҐ^��Z���dLT� �N���!3��C�*7?�~O��Ưlg��G=���:�Uo�fZar�u��E��	��V�ƣX�ZCBD��0��+̻���]M����1,H�M�����1�h����q����\�T���abDUu,����]�"r������MD82��(٫��T~[��� ��K�J�Tx�����	�$&�d�y
W��yq�c�q���9:�/s��)Ę^)4'�oǢEh����5��KJ0_��)(���@���RR^�ۂnrm�&m�:�\�9��T�&w��l~��B��)����r/N�/�5Rk�1�zs�f0=!L+��i%��N���P/E/���]<���p5��Y��4==�W}���j�(++��HV������X�tC�������q.���rmA0y"X��?���-ه~ƀ�Y��3�ř��)�
AO�e��ɩ��V7R9����Y(6r<��D�V�~,�Hz���1hV.ݑ�ܞ�hKŕIU��J�Bk~�Z<q ���3��7�x��{T�d�_��0E�%l�l*��b��H����232Lߞ�j��+��_�n���1HII)�pσ�
XͣeGqbx��F�1/��%��?��pL#�,R����>�t`d��d3�����ڌ�WW�Eބ��z��@���Lq����ρ��Ӻh��
�~8.[}ו?[i?{^���Gf�i��}�ñ��l�.��i���4�h�����27�n,
]&ETI.����R>��$(�0
����q�B�x�]�z_rt���T�x�E�RY4Y�.�j=�P{���3��AB��=
��@x�ynH�Ū"�e��f!^Ř&��#P�$������[��eݻ_����CCC�c��y�t,6 	� �K�=>�%�N��[U��L2t��:S_���l����
�5�˺�{���6� W�>���3���.�&r	����x+��~�����T2 �(�K��!�@eb>�i3)�0��3���wl?�����?F����?���:�j�"oU�>`lXZވ���.�y�mD^��ӣ��R���7����l��<�P���ڍ?	ڕ�+��p6���̪!\���L��� 9�#o:�A���>�ҵ��h��7;�	��G�H�xe%$�蟸��zÕrrn>��L�Z/��tB���?��'43�;�Q�u��\ݨy�ZS~�C�w},~����x�c��l� [�~��-(%n5@�%7��2��6�O�������3�v�$��yR>ψ/�z�c�����X�Wf�i.`x[�2��.���-_�� @����]����_�w^|�iL�
xW]NJz~����z��;�.5D�j�f��z�*M�_{)��;}�P|��d�nʔ��N;�Ԥf����ݬN,�lc��%��DsS�J�� Zyd�o�Z�n��gܖb�3�}�u�Ѱc��� M�1͑l}�V*�I��+�ǌnd�4�A)��(J�Rah��%�4��Q��'	!�������烎`��!z͸��-�^���#�P/IyyQ�$=h�9�M����d/��o$K���ƪ��,`sx�K�:N�%#�&~;��ڻ���V���p�OM��9�l��l�i��W906q'shJ:���ۈ�;�R��'�L���S{�#��$�6Qs�w�=3Ln�z���caǒ����P@�r$,��Sʔ�3�f3�.�)Q��W���^�y���*����w���9��<eh()/J���	��u�8����_݆�D\�n�{�j�QG�>�IYQ�V�;-Ӣ��6TC�����^7FU�/�n$��S�q�z�;�6�h��H\1���C���&�bp�J���q�P�v#2h���ݫ_���T��FR��+�$�m6����k	j����:ͣ��'Wj�_ r�:0#�"D�xͶ�I�:�+���NLL\����
ڀ_�.�x="極��#�G�6e/�b�h+�(�H��<�HߔG%*�zj#"!5��|�����q|�����zӃ���wڰ�H�\�`����Z��Ȯ1����%f|�XRW�@���-�� t��5l��8�9�����#0�Ԉn�}�{��� P�3��>��*:�(�C�3'��;���G��Fjd��U��,2A٠�~U��5�|���.V�AI&�KI�7�,���~B�ߚvyC��Փ���|��8���R��ZN���+\o����ؑ#�ɟ���W�F�D�Ku�Jop����S��M��H>�1e*!�bP�ۛ �1����!��G>B�0��dRk�" �L��fWdk����V\ry�U  ��-w𢦱:�_6Gab��$��o�|�b�����׿��ɋ� !�|o{X��?{�#N�TaB����ȈW�
�G+�X�J�GԨ#����zwjؑ�!ѷ�� �Q"��Ӯ��v��k��6�m	�$y���^m�)��3�AT�Qlt?��zZ>#
�܌�W�-�|aa�o9uF��q���c�>9�{�WXԣ+U�i��n��6ۭO��(�Y�bs�$ڲ[uC�\r���;��FQFM�L9b�ǈ�4�"�](W�F��\ݫm�@��y'XL�ɛ���7L�!��{�;i�&V�B��|�xV���}�E���>���R�B�a�O�n�%���(�b�u�A"8�v>~��Q��P�)`��ե�?�cMMuw���E��י�p������M���՞���qSK�/z񊒯�%��H�6GZ�B��AD;�/fl�Vi�؃��r�I���2w�J�Z]���{:���'�^�H�b?K�7���
2 ?e?��~-G��DDM3�����ݗ�rL�bX�6�M���H��p4;��S���gu\:x��Uqy-���~�GH�猖CE�o�4k ��[���U���W��y�C�g��6�E��o��=���|�m�vs��ڴ$93������2擷.��#��?Ah�H��ڂ��;}|���L�Ce	ལ��._Qh�O��K'/�&V���
���Х�J�?�u˵�
^z�s�"R��!�Mo
�("t���9��B�L�Z�V�y�w9%x�գ�{���cA���OG�p���T@Ɖ�'R�-Q�?�H��6J�y�,����{��F�:��U��n�}��Q�]Cod(�
;d���؂T����J�n��������(;�Aj��Ҙ��"��[�_Rj,�f*�I��w�����w[j��WW���y1�)��2�y�Ħ����oR��Ѝ�R)���?�H�L�fp���kt}��rK���:���@���K������k_��ޮ��gڙh&��I=�����l���L��i oݪ_�#�jlbb���7�%{�\PA�����Z�@7�Ү�[���k�/IN�hJꞪ�n{�l�o��ئ+��V�x|�1:in�ȃ"� <�-c�n%��/��.�����-��
�F
�6�T*�����Yr!'��j�k�i+�����A���=(� ���A&��4�5JJJv��1���z}$I�aJ�)��%%���%��P��w2k���F�M�[R.D��_HQ1C��v��C�#��QˆFayg����@�]|�zjUn��n�������{j�	$2����nD�ZQNQ�}�ֈ�Ȉb�d�w���Ը9�M�$�C��3�Z+S��;_��(�9E��n�Գ����=%SC�,/6�P���Ec��3���Ŋ���d��i^��N}���N3�g�QHڈ�_<�����"�lj&_M����ۜ,ꃢ�/D��9�|P��$uu����Q��<�8�8��_���l~����;9�L(/��O��O�*�__����bd��U�ŝU��������ס�n���Tw�U�4<����d�I?�**1$hU��oF�Ռ�yP�eu���2��f�R>=2g�O�{��)�f�� �m��Ay4�eË#�w�253kr� q?����X�����ݽ?[*+���A�;������%QB��.,�Ѓ�ND5p��;	o�j~�����&M]� �A[�U�5i6�q�K����t��N�&�j��馗>:��c�	�&����;��j�[TŌ -N��$\�7N���ď�z�y�X
�ye�kJ�������}ZE'�{�!P�����_�����P����G_l��4�-ZS��JS|�gs�Q��+��vf��e���-<%��L��������7�_�����Sko"b��1�F����4�F�SʖX9^Z��ǯ�vyrΑ��@v������G��?�#���ڤ�Hr(��#6�47��f�b䧗�6��b@/��/I#�y6h�,1w#2gz��DBVS`�o�sts���7RDB^�V��h蒑	��볠*$���Ug�JqR�ʅ����*�W�˓����^��Kd�ԍ�jT��^��~�������J��њ��o��'��R��.�s�l@1���	�TyLI�#-q�X��1��q�f�{�x�ɿa�$ಏ���8���5��[4��Eh�^�P1٥�v�����Ԅ��}Qr|��8���f�@��c�0Z;��-��=yh���2��ԚuN��<N��؅�￭���_5�O�"G,�� A0"��(���NA�!;;�ӓ���ס����&�U"�������E$l�xMM��J�`�z[<��!��`b�������D�]a��n�;9��Um`�����@)��x��,��&������<O���oS�lN���X��RX��V*C! @�޻!Y��'��T$x��tbaO��>&�˼`玫V~T̵mZZ�gHԥ@���ywd�O?�ź1�؉��<�%`�cX��L��Kz��I�$����N�T�oC�5�u:	��M��%ܟD��IZ,�W:�)�3�F��81�hV��Tz}�-�ԭ�r7�����6]ȼ�4,x�
/w&c?d�Q}q0)��"���<B����%/�Dd�����D��mR�,� xw\���#L�Vv�}����Dˏ;������3H!�t�:�rN_��Mޛ]&W^ۭ\M�d�9��m���Zݸ�"��wp����IQ��ϋ���[/�o�/�Pr7$���,w��S��||����w�t��J�������ȯ)��L�x<��NV��9bb�8��+m�ip�YШt����UC[fi���ޘ9N=n����6E����8EIRL�f;`%���S����x�����)�<�T�*�׭�1j:�v�
p��}�R}���/�"u{(�Ì�0�㗌@�M�sC�.�2�c;fi��'�gE K7K"���%|�E�E�6�1�����x0��_\T�;*���R�IUs�71���c���j��۶�ƶ�ƶyb�nl['I�4I�mc'6o�q�?������,̹���8O���t���9%x�0R�C����8{?���@(�{�}L��bu�=	Zk#+�t��*�,�_dp@pD"W�D���Jء_�X4TU�t�J	?ME��[�L�g$!��������F4�wf
��Fe'��:h�;?C��Z�B�>�'��frk7s�L�V�OVrqn���?��_�����P�Izz���Dw[y�.�{/�SW��������xe&�2�l��v�zI��L\�� \�Jn�V��~�M�踢�Z ��=���4)W�֐�xP���;�����]qo�)��?��[��4�� g�(�r��,���u3>��a���ARAS)�7x`=)�ed,)*ޣX<�KF.&r��8�����4r��(��bGl��ܡ��y��=T�'���2�*,����WR�}�.���6�3�U��t��K:�h��e�q���N�j-X���ֺv��9�%_h�hm=\�ĕF�O�	H�͚m������=�����[_J׋|W-U8b��@����\�����x��{X[7U���%�agb*���c�\_f���9�J�R�r��K���?
���+*�߷;��1L1��@�����v�N��:��5�S`����+ظd���@һK�R�1*S3?%dhi�w��%�?��P�x?�:"�֮[ao[E�yE�#�;�/n�l^�e���o������D=<8��q����V>�	u�ޭ������7����(�faM�yHHJ��>�j���RE���.m��B1��	?�2���������?U������
�x�K�E'F��=\`��bc�/�Yw3�u�`�S<�!�Ǻ	8!�{Gӊ��'�W����)���3�t�o12ϭ��ذ/0h���°m?�D6u��9~y�{��b�d�vF�%�ڡ���}-���jΟD;�'4-�����!S�_�;X9K���tK2��sn�.Ȁ�*9J�=�5�<����=9��~),�'�L��;U16&�5�͏���9�a�jK���<ǲ�F��]��\�-�"̗��	�]&F��n��qK-?u�]x�H"E���?�Y�ζ8�`=z?����S/�-�>6�[�>O�;zI{|r8�B�B@K=����z- Ec��;r��J�v�b��_8�]D.NA�[1�D�Qn�S
T�����1��'Ua�X��̼��y���"��,G�"�4�g����N���	�!o��D݂V}��:9�$FnS����nW���E�,Q=�\� L8<������;_|��n�H���zT�x�(�����畍���Dᄷ�gv$^4'�s���d�p��Y5H�]�:4P�wq\�`:�tڍ�w_��+� 5����e�e��L�c|j���v��m[]�ӥ���L��xƺDkA͡H��E|�G��}��k�,��Qe�%H�� ��6�X$R	�[�q��[$SQo�L
Z8����#�(I�{ǜ���CKQ�㻝��x7�JI705��4F�\;��aTLR��f�v %�V��tJ���ے�H1%-X[��/V��8��榘H��%����0F뿠c�����Y�e'�c�⋗�^l�:����а_)$;��Id�)���*�DZ�8s��(�;(��K��ݸ$�7h]�LЇ�7�ɞ�/�cL�U�b�w����p߳^��c*�.˴-t��^ʈ�X3GYe�W� ��9�@\�-z�"^�ʪu����00�	��Q<6W��,����;4X�OP<Y����9i�Ԍ\�=�Id��6�):A��o��?r�#wI��cM&�2f9j38x
�����g<��.7��] �$i�@2L ���ֆ��3y�u�}�m%0�ɵ� -8!��d��o�dW�v��8D�T��n��<d���Q_ ���ꊙbp��G:��>�"�s�7ßV��S�y&��7��w��V��i2� ��B�>R `7�j0�kf�|�\{�Y8�ӗ��� �������/����"P�6����D�pI����g*�з*l�7��R��J!���K>�� �q������D6M?�y?���B�V��Of%�Rz���x��q�@N�U1׫�/i����~��o��&.fʑ+aHI/��������>P��E~�`;����fG��Pg��<�#���Y�� @�Cם1��M��-��[Uu��J���_��y�(g��Ք�k%�,�Q���z��E6�Ձl�� �P|����T�f�乴+�i�5��+W��㥡���'y�:�]��J'2!m�%]�2
1�

�~`���1�7�t�<ɡ�jv!�y�ܒ�e&���:;87מPȯ�D�d�$�t7|у�	���������H��|���b�{�!����Xd=_���I�s�%�Zb��)S��`6x��Q�[��I��{Ag�rew��-@IC*�3W����|w.<�t�V��z��'��:�սN�� �Y�a�t�
8��%�� -�Ū<	�fF�/�X%�Lp�e������N�<��#����z�a��+�|@����w �H,�)��^�k(��C��2���h�D��ag&Q���C��R{J
���*d��dӠ�������ˬ!o��U���d�x�?�G8�u��<\������uM�I�C��3�|d-�/ʄ��?��T4=f�<7^GS$����=G�~*�\e��'�뇞��/�DV��Wjm���Ჵ���7�
���A�!��&-����lj�E������T��R�����'�*_Z�m*�E���U�W[<���G&$av�W��[\ᒃ�t[M��ui4�j�y�8�B��h�ɺ�鏖��N	�����N�D��ǈS� �L�M�m�-k�:+��d�������Iq#H��R�h
�2�T��UAw��:w�����75y�hs�d���m�PF�-E���o���i2Y�&W1`ס���/����N��Pߙ(�eO��+ġQĔ����.�F��@��?�7�཮�/��M����U��b����v��\����}����i)eQQ$��P;l.p��B��$�3�7��bJ� S���Ue��w'F\:���k���nT�i�rW��6}�64�
���=8J�6��S��y�K'�Ep4��q�MJ�,5�uU"^�&qc�1�Kj����_*&��s�0���m�kT��R4�Lw\^l���T�qE�LчS��-Q����-`
�x�単��O�Ma�E(�?B`�P�b"��E��=�C~��(��`J���������AA�&z.��������o�Q!/LS�k�B%���Y���g�Ǔ�\�%���zʭv�#�'e"�(�W��.R!��c5>F_gT�4v@.Iab9�k$���`�K���<з'9�W��=:�Lu�T~^������ F<o��nL�B�lon���8I}U��%|���Cm�ނ��e��f>��r}�3%�򫟜f��Ӥ�����x�. �H3?STʀ��j�3ʙy�z�H��Mb�~	�J��8��߰��9�*J�Y�[0��L���:�f�9��n��ڼ
�Y���|�\�P,�5���X~����f��~:CЇȉ���H�!�%����es�$�b�S�5A� �u*��(�ؽ�B2�6�Mp�r����F,`3K�شB�d*��_TT۩��1I,S�@����Ih�۴ﲕ�� ��e����eK{5Wc;�r���$���߻�W������[��S����5�u�Q�=\��ҍ��[�nx�.{�!>8\�a�n��(i|���C <�d�z/
p�{��ӫ����wD��/�-+�xp�Ẋ�$��9>��ۚ=�`�~�ς@��,b&$����h���s=l,�<�NQ��x^j�1����!Qp��F��%
#TSq���?��i�C)���$qzG`�D�����'�f"-[������{�
�.�8ːC��"�Lj���k�+H�B^�M'ڨ}[���c���L�m!;���r�{�ϻJħ{{{�6�tt�ޕꐹ2��=�,n	E����1Ui�o/���l���M:H=\��ȼ��98�����{����8��>\�`���wD"b�� Wa�	m�����^4�dp�y��y�ރ���BH��ָ��̈́J���ӷ
ٰ��C�Y�w>�\Z�9(]^����(����t�Z��=���/��#@K~X�t��?U�&Rur
#��dxm���2�&�\���aɎc~���O�s���a^�Xϓ�]Fؕwg״���5����t_̉�[&zU�<c��b��|`8�##��d�{_Q�{s�[,�F0��������;T���6o���!Pr��_k�����z\���F�6�H��J~���@�;@ɻK,��I�'�J;7�����`���/*H�j�BT�N�:�Gj�rܩ�{��3F���^+V��bL����KQ�i*�5CL�$(B��<=($ur�qG�}}�g?�iYn)N��@2г�c�>�����#��q29D��6,�b����Q?M�Uˌ �#��}������j��|��E��0�ـ�bg��~���C�=�A\H��f��X�p��c�Y���_R��lR��u�{�1�ׂQ��D��w�rt��~�.���&_\��EVF�|�;�� �.����WH%��1E6�Egl��J�dK��(1�+E�#�}R<��(v�t��Ն�5R����ַ.!�?��ڍA�N�>GTPZ�	$��ߘ�`�=W���k�E���
�x_�hNK��\5�����Og�+���Q�:�t���"0�AP�7���1�p/�BC��S�x��SO����<$�B26>�,+%���<ڪ�I"61��fI�(_q��Ei��O=�eB�a�H��'�^_�HT����es�L���7/����ed�%�89�:PrH22��r�3��|�577=�M�Z�
���>�Q5O��`cTT7^���=���Q�Z&G�x��ثڿ�j��t1�P�|����c�d������x�/�`�G�"X���q:pJ`1�q�(�Kr#Zc^�F���=����0郳{_�k��?|vS���߀����p�H����\��-6�Ԣ� m擦�u5����f���{Nn�=�xz|փbbȁ��ft��+�'8=���=�D���>�3���5��^�m���+��k;'r�.Ğ��g.P��b�?�|!���ێ��diO���)�5�`i�O�"^]��q��Ol����l�"Y'�s,��yw�ī�x�O��F(�� �nGUWs|��guf:��[���I�fx]��l~��K!ۥ�^/I`3X����Mbe�(&�c�J���|
�6�.��GGW�-���3Z��R� ������f���0�i6n�ϺP`P��X�����++�L��)�����߷�*
zw3��f�W���6=���b�}W��@�.�� o�4<�]4M�qx휐����^d2�nJ'V�n�ō��~?���ԅ�]��~�������y��JD�������N��.�m�׎��˗�|����h7O���3����?|l�[d���A�������u����aX� ���� >�,~p?
���\��&�~<�HЂ�����g��ĂN��m��_"��h�t)h��p�i8��:)�豭�Z��3C_���(�$(�+P�zz�Gp
p,ڷOC�״�6�uq`�kᛱ��T��6��y����y�X�+�'A���!���)��TjJ�7�5ZE��Ihwm+�2��Rcִs�'Z~��pn�V3�WF�	"�_�� -�[b~Wc4��~ˑ�?�,ie�/K�ϓoE8�<�9�`ywl%�]�k��1�aM\�������O孔4�� ��l)��J��[�	��v"UttC��(5�"�7����V,�$�L�w��}�ɩ,H��&'[x!"��zo�wyT�Z���>y��'O
e�dF�D�4��lΓ&,�y��3ǥN*�����0H�쭖[;UUC8Y��{P�RKE��w�V��E2-2}ي��\�Q��:n���T�=��&x�P�\�d�m�]6l�� ~!ۈ1PZ���2Y�FD5^��)��m<��;�N���p�k!��S�+,�('Zef�	D��>1cf��D>L����Mb���5�-��>���z?8��e�g_��K��VK�g��P��
�bb�r��&-Y�+�˫0!�������;�G�Bϧ~/K����\�!ih;3�b�;F����G+ZZ�I<W��f*��T(��sn��	��g�Ȕ6�1 UA��\l;�G��9�bS��N(L͊U��1*�U���������29��M�f�D��,�g���;	�1�2����{�=2m�/�O�E[����7�T���A���D��c��Z������W�R�%O�W9�\�W��+O�u���ac�<y=��^�|�&����G��Q&��}߻ :����������*P�0�t��_� ��{{�k�o�B�j���]�ou'-?���1��/M�����O5kQ�SR;i���~�T�������D3��6躔m -b]�aP��y���^�\�mOYB�@9����̝�a�V߽d���8���wT/<=]n�(�4�0���pK_t�Mf6���9�ѳ���He���Ƹ\�@�Wb'���n�ʲ\'�zH#��˼�:���c$!55�$�*��뇱Ϡ8����ȊQ*����A�:����`���e�딞����#�A�Q�����}.�4L�|��_�NB��vv��O�&�[��������=��d���=�}}�����=唶|J~��Q­��'������O��v��E	+V��\�qH���8�߷E%\������k<����X���b/B7���1G��b�:Dׄ�6]*�G$JN���Z64�͒œ!��'�AxO�U$3 ��!|��5������V߻�:o�k�\d�=V8R���>�P��ևA��R̥�IUK<�#F��VŜ&����+�cN���֟4U��w]�	L�lQG�֞�,����a���zy����TU�;]��D �61�`��M���	u��*xʎvF-�X����z;��⢶��b��C�ƞjՁl���A��!���Ijj�N�i�����	���P^k,.w�T,��@���l�Xq qb����8�Jҷ�+1�F�2�xqv	 }-�&I���u��Z�2����\�A�j�ކ5ndH����hz�:��~�}��� �7�/�i[�Z+"�ۃk�_-�����1����$��W��M���)A0��k��,�� ���'I��4��x�.FY-A���C�	b�����r`*7�L�b�۱y}�M(4�6]d���[�G�{VT3.����4�ƽ�����n=,���4��x(Lw����=Z��F5Uz�����.��o�g����_
�`(c�F{HAߞ��F>��g�;%{탴"�v�-�|WPZ^�n���@�&zF!����LW)W��_wrbkjUܔΤ�~z���ba-�f B���il�oj
\�:�*���f\>��	�x�������Vr���";buoK�2r�dOy��h����hw�PJ�&l�-��b�)�s��o��m�k8�GGG����B ��ĊJ��?�%y�U����5��f�2�u�ּ�:�iSc�W�P�h>�����cС���b([V�1�n��+���2�N�s�۸�"%��#�{Z<�)�<�p;�]n������/���0����A��a�m��g�9f����=� �F�;E��즴l���[>O)E~U�9y�$"JM�`�\*�P���{t��3H�vؽ!E�.�P�m𹟃��dc�{����ߏ͢}���uWP�#�$<E_]M�b;��+�3��@hC�S��
�w��z����Wi�'4j���SڑD�Ȑ����p�'HG�:]��3�s��\�C���V��jר�f���Z�j�t�ۨ��l���IIQQK&��	�VV��O�{���Qa7�w��M�0ĺ�G�6�RX��Fu��!W�[IC!��(3[d��PխA;H��C�ˆ��(��4)g�*�����.j�eHn�^����2_�ݛ���H��Dό@��2�5L��o`�ELl���uwC�&�5��B�r W��qfU"�h	W��=��D�M�K~��#]e~+#���x}�9��r�;]��=)����=}l��K6�O�bkY��
&����7q
����\�����,dH����h����E��� �>��}�-׻���֗I0� ��ҤV$�U�,q��$cc�ccsV�$
�W�Љo�G�n3�M���=XH�**м��Ҩ7�j����a���= x�
��<?WDSg��f�l�/f�,&[��C���!�$Հ3g�-F�:�*��L{���}h��drR���gv��/O��G���騸^������) 43�sT���HD�o�0�����^U[[{i�wT��|��n��}�����Ʒ\ه½L�i�,��ؓ�6��0ơ.�0���okۺ ��zxʢ�;CL0��uH5Y����ǳUst]HU2ϗ_����]�]܃�S�����+m��GwM$��Gj��^���q�s��ɹ����g1���j���@j��2JV0��
��/q�?���A!D��%��@�b��|��,�����i<v+0��r�����_c��:R��@)�l�%P��4�]���\	:�
c��)�?!� d�U��H0	�x�W����u������ݷ��w��M���I�@�n:�k��Ih*Z��&7����G煇7����`;�v�����_|��c as郦 0��袿7�ɾ:2��N!窲�K�
ϼ.^��q��}X3Z�OKOε�>}o�M�K��������%K�N��*��7�:������������-�>��!185}���*�%$o��#����Τd`�,������(�׍Z���Lٔy�7�02221y�}����L��60P��hRB[�1M�Uh��ys�A�$��kYN������K�×�{����@��B�#��3��##&Gs{Ab�$"��ҋ�����=��S�G�@�=�����%��Ӳ캱ܦ�I��)a��M�r�ߍkZ�'��3�V6�h�y5�h�����+��U��E���.iƉ,�e���Bu¨���h�ǣ���XX�N�r	�>���P�JنŀKd&�)��*�x�V�jO&fL+31*���,x���Ngt���D�{'���2�����/�@@c��-�ׁ�q%���Y��=��8���b�����5dz�Y^J4{����_�E����?��A&t�*̼�M��3̺�P�e/_�) !r� ّ�~#����pf��m��X���m��sO3�i��J�Yf����SCLQIX�bj|��\�{5��ی����>-��0��<n��/~ t�RG͈�x��C��w�@	])�|�}�e�)-G���E��Ώ�P֡fhH�QR�B^�8߬���7xJ��3k��M�r=�uW��N�� 8+���O.;!�rt�N=k?�/���9������3|�y�<xp_d��^DO���~���b�?�9My���O��s}�ӑKH
����f,�f�m#Ðخ}š�7/F4z+��o �s�X���b��mh ��q��0�����&)�R�"��
lt�&�c��W�����tކ�*yUY.��>�Q"�Xۖ0=(���F�2��K�B����W /m�mdn��ɷ�c!�_)�ʌ��f������صv�����D��Z3�{1pY�Q�:�"��������m���:<n2V` d�i�2���7c<(�1�(�ٓ�w���_�1~ʠs`˝�1��*���M�ӿ3��!Z.g���R[
q�hE�&���@��z�����} �`�k�Q�Iw���rH}�'
��o>�je{��j{+�DJM���k3��~HLc����A������-`<��|e��&�2ֈTX����:�����C	Q��`J3PVq� �WUu��d��^G�vf&<��#P#���;y�Z���e%�U�3�z�`�8XƳ4Mp&Z�fN?�
�V���G��h���o���ܾ���h��'7�,=�ǧKnè��$�l���x�<1�1w@���/�ǲ��UX }�ڙh�YE�o�zrnZ�U�-�r���n���������i+���toU=�����[*,(0�ɍ�!]�R��d�B�"]�y�r5+��4��}��=�1g����⛳����!0j��e��D/
#�^x^�ngŵ=��{��`�^H�i��A��b=�5<ǀ$�@�S0�̀��&�H������_MȻ]�!C���6�z]�ʸ��\�o��sҧ ��<5Z����7W�H�dV�9@��nEn�ݶA#�`��@������r�����4k�S�`v��y\�b{;v�zzjlx8�@��Ԝ���$�h���|w�a�+�y�=}I��@��_��ʣ�T'A*sj�� Xz:��If���P�niyIs7&w�ϩ�0�am��ˁX���?�\d���+4���"�G4D筴S�#c%�	X��v����!Zϐ�?�D��'��~{]�����	r'�A���u�F�$�
�i%�ń::��Fi�u9[n�ƫ��ii2���ć�������d��P������}`��r�Q֍n�\Ԗ����Z����.�B��;��+��E�	S!�gvE�Q�]�^B�V�'sݢ�"���Y�-_��T5�O2]s�5��
	"�sG�	 �F�_����K�cbQ��9��R��7���T����
��﹗�F�y�C �[c��<A�nk�29i|��]�����'�v>�����=����vf�b�dp�������d�{:bE��͆�w��T�s���1��\R��-C�iS!C7�롄�m'MPO���d��J��L��FM�K��\87p/*�Vc�4����2v3j�
�a}�����V�Q�l��t6=�������8�8b_.9�	=���Ƨ�o�y�����h�E�%E&l&�);xڈB.��- 0�[1�+[<�u���ܟ�~�*��!�v��:��B�H�Ёx�Y�V�s�JVH�~_�>��/���6A�q��5�������5�,��?���[4��ᰜ�Z�K� �6�7����q��X �2��ˑ� �[5
�uB��b �i4mQ�����3����{F�J��Y_Pn��K���[�A�5��<�c�ڸ,
�)	#��5�A�p���n,ۯ��X����s(�kQ�`w���&�_]hL��a}[���K{Oʰ��B-3/��=Ž�:���B���&jMh�9o���rX�^n�ef��y�����Y�B��i{c^d�PO�I>���W���mY|��N��Y/��̝IҾ��,��=̨�Ȟ����7y<ښ'E���ѐ���(�/Ldy�Q���m�ܜ��ˍW7� ��gi��p���@+44�ܞ��#�(f����;Z�  �����Ri��^�Y��������G<�[�T�f�Y�l�@�t������Z/+���7Kl
fN�Ğ�e��2y������]�?Ы^�4M��Ѯ��Z%H���|h������{lH�]<V�Ak�G��*1��f��Yh����o���W�O�6xP}�v�y	�0W�4֔+p4�TT��ʛS�'�CK=����p�V���X��y_H�)a�+5���`e�
����c����WSȈ +��T���\?��pP�Lְ��}*��I�]�	��[�~FQ~C�أ�Y��4u�PY��g��F�l��Y�e�)0v�{�Ŧx v �i��SeO������B���j�uPa�d����8��z�x�����W��:���H�MǯT�3���o�R�Y^BW��C�،a܇"���\�N��$�h�w�);=<n�<~�^p1 ,d|V~�� ���=�1y�,�#WTtPt����A�0��{5:�Ϊ��Ϗ�l2y���q�����a=�o���V_��f��Ȇ^^�(oG��b_�U"C;��f���*���<�.����� ~�is\�����������~��!�D�Q4����m��~��E�Q���snV�Ix�����x[w���KL!<���m����V��;�(��Snx��/I}� L"7QN����Q�(~Y��S�k �Ƴ*���+��]54(���5Ţ0���Q��viw�}��>3��R� ZL�@���#=��!�H��Dz_e�s�RF���������`	���Zz3��B�W����[���]m-���A�4�cu�\�n�<Z�KۤBC}v��
���J�� �Vad6�QB����DP����x��Z�}&
_���3����k	`�@��%�ЌN���0jaAe�ʄx%����ȵ���C?? �h2B+ؿ�`)�����S_o2}���>]y����T�wEH8�E��/�;g�%Q� ]��]Q���(�ۜ�r5�eۇ0RY����I���Q�v��C��0�F�&��R� *X?��?��U�@z�yq.M�U�l ��f!����6Mc�V��oy�s/�t������a�+��Ya/}I�(q��=�^����!GP4��ʐ��[U��3TMr|i3��jlE�f�U�Cq�8�BD�%�Qb��N�K��t��K��8FX��ք�`��U���/�^�O[0!��Ct���	��a���T�=��Ym��B�c�p��c!#T�y�?�Q��aW�Dt+@����5��>����1���"��(��� ���b��.�.������_�Q��F �a���N_K#`�әo�p�^p�U��=�H?�j||�d���r:�!��]6�3�c�#4�3��%
m>��r n�rz�x���N�5��B6����|'�4�����GE��2����r�ލp�{�d�3�`�B�a:7G��ʝ���u���T�8�[� ko��g�.�*��vq��N����wg�AQw�`�VdO��]㳚�"	xU8���"���� ��H7��9md���@�X�U�������k-�yl���3h�"�]#<���*���L��3��]
�S�{RB�"��:�S-�nX��B��|b.�jMhQ�m���.���V�[_ �!2�`�Rp�kK�!3�Rͧ#
���4���g�(Uc6^G�,[�F��j�.�7���>>|��	���r�ZO�s൶a��͏ y^�)d)�Y%�����T�Gd��[�^�WA�mF�[�T��n.o�v��9qy�e^Ӄ8�i;ʒ�4�[2�k����8zm�h#P��f�w���3��"�n��N��A��/���n�#*�3\�Fi���ŰQj�m�������'�0_���㿃:%	�!�W��Z|�ꌢ%� m��.V��P�D)�o*7[]��Z��a���Â͖��I��B:a����{��!�v���8b�'��W�����
sDt���Ȋ�I���f���~ذ�������I�}��U�A�p�!�E.�ĝ�H�����Jo-П�8i�M^�����$��&M/�����b}�6��r"�kOd�tt���f�sRV~�A��a6Z�#4�2�TR�'נ���66����h��� Ϧ��(0��5a�jgZ�U�0&�jf',u��]�8/�?����t�Y�1�����S������l���󸍌�Lˡ�A������b��ݩ��>��z�4�5���y����WW;�N�at['1];� )LN�û��H��/q��߅F(��M$�i[�]�S�P_>xg�գ������Wl����J�BB��$S��:���;VF�/�/o�=s�!�H��V㒪��⎊�Ɉ�Uop��:���%�鿎���G櫭~ᅉ̼����J�� ^>[�$�/M߶�~��Q�����D
�s�у�en�p6)h�M��q�������	��� ��L:)��χS��/fS@�R�M��M���ox	?�Q�Ც�.`���7���[9"�����.���؇j�2ݦ=7��,f7���4�γ����d�K���b���|��amUL*���_u��0����--8�{O�K�g�jS�!g47"��l'D���C�����1C>�;5Z�:Nؑ2��c��tqiy���m�IDV�.��=��`�:Â�n5B���tf�#^�$��.j�dM��~.��fF)[h `&��38���'7aűQ.�۳Kp�x����y
}��:o�G��Nс/�J��0�1���m���>Cx���{�������dy����G�nt�YG�#�'|���Hd3�#2��� aoXkЇ�q�OiP�O �ېLɧIy'n$7�i'8� ��%Ʀ]G!�p�������zR~Z�A�7�D�"B \yk,b0�=�BtP��
hD�r�-�e��b��o�G���:_�[��c{�B��ߖ��s-�  )��,�]P�"�I-�}��bG1bވ�ʝgF'}ÅNե.<�lF�M�p�Z�fE-���U����!l�kf�`K<0�b����T�.b4����=wr\x�����`�:t���"�ǰ�Q�r#�\d�d��=��H&�85?��@]��hJ�����Cp���Q9�M���c��fØ�CK[5�P�*�~���M&����k�>{Z������jp�y�27�����9���#E�48m�����y�y��@�a�Ѱ[;Ӏidqa��S�A�h�fT�A��9(��Pw��h~�	rĎg�#Շ���V҉^���t,��ZuT�o뚈�h10���d�`�M�`u�-U̯����՜�N��+�7���g�8�QV�g��E��j��:��|�����A["��)#�zJ���(k�o_D
ފ}z��CMM���w6����_�=��\�i� ���Ѧ���[���=4�{B��F�9��A�NN�Q����Ⱦ;%|.���$�#F)4�L�!F��B��7܁6]U@�w!����u��*ZJ�^�_y��c*�ub�h�i<�g��ǉ����y�a)W`��}hV�uZ�DE����)��lGJd<��	�G9�	���[���{�-� � Aį9mKs��אs�����/���c���R�7H������&@��'jPPq�9��qQ+e#f`X����*q,�Z1D�;,6[��-�}c�)^����#����օf�7����G�� G�_��/j5i��f��4����k�D���қb��Z��)�e
�"([?Q��,���9M.�ԧ�ײVFTϮ�ih�7}(z�6Y�M�����d�-�֜�h<�h/@ń&�#���+��Diڞ�.|���14�g.
�AHL3Ћ:���P7-*^��|�@��E����d3?�ۤ��W�	�,bCwܻ؉'ŭ����T�Df���}�>Z|!P���d�&�ZL���5�1g�d<���<J^,���&�q0;t3$8�織���!��a�k�A���-�\׺���@�qǍ[�H�u�0|�*I|�,l���>X�h�Yg0��9��ў%W��!���%Xd;��+���D�j��%��x�U�c�f*65�mtȀVfT�K:5$ebs���>TSW�K�yNrk\*&G�!$FƧ����8�ň����C�wrNb3��X�,|�О��]:�*����uy���+u5F�ݻ-Rl�_p����j�L>� �����	J<6-�+�#���|�t�Z�J؈���TX��=2�.�i�~���TJku�|G4��V�6ݶ�¼M�6M�@J�*�f�R��HH2�����Z�SS�F��h)t��#�u#ـ�	��a�dUu���YE$�1#	�f�b@Z�ܕ�1��#NX�\#��ڿD�D�7X�K٫5�v�
*ʭ��pF�ur��Dz��]�`}d�'��&���)`�u5=�c�O�క�tn��p�Ww �u&3�=OSҢ]��=Z�RS�K�1����Y����[�vKܹ�D��s�Y8h��0c�]�h(�e��qM��p��}��Ϣ�%&9���" �3z�ʘ7�9ڃ��P���z#(Yi����]4����KE�����J�I��]��|�V�$�WwŰ�u�}��Gd���e��ߋP�;x�?j�p�o�j�V�eee��9܀��,B�����~��0���������  @bUZL�6a��VZ��g21�l�)��;h�>�X�c����-G�3��������_���٨�/v�"���Ʌ<�`~��E���ܶ+�b蒉�_����*��6�	�P܊�w/�ݝ ŝ���ݥP�)�Vܝ�Ŋ-V���y:OI�����Zs.���-�NF�eSf�h����͕(zN{,�J؜[�z�n�,ԕ��c�3�ӷ~)V�ĭ6���Ź��n$Q��4qgM�����J2iD�	�1���xb(�%���u��(�R�S¤8���Lf���/{��$�A=��ٓT�x�<��_%G�����C��Y�kدA��h*p�*	�u���h0��:ve#�s�FF�R�'�1[��/�
�؆�3d�Y���b�+�ߚ�����r�X/�3��;��&:����0	Z6��a�����b���"b�ʔ���V�n9@�V��A�;��@PE�� �e˟	���"�lU�����B���]� -U��tp���V~kc����O��A��K�ȫh�D��RՔ��o�����Pt�"�9�_MXի���|�ʲm�I(��"+t?���@�&�,R�Y� ��

th㦕����^��:4�!e�p4�R�Ԇ�){p_m��0hN����d��i������k��अee�f�v^ɑ�Np�x�՗����F�Qq�u�Иl]jj�k�%�e�}"u.Ǖ2|J�S2�6�rud D�aU�R����|���B�3�iM�r^��TX�S�����>\+���F�(Q'���۴;�j;�tJM�1��Ns�ܡO�O��{^_���w�en�]��
nq�qG6+��`8˒�Ҁ��E�sN,v,+,�������(�d*1�����Ү�WL@z$'R�a�p�!f�F
��E�!:(ҵ�a�����f�ވ:����:�I��fb�ݫ�z�h��*	DՒ�>:� ,&;��ޮz֬��*/9�ou���k���6|���FGFF0�g���
�r�����Il*<L����2"�4��zP�cX��Ҫ����~�W�)Ͳ��8��|��>wm�O���*���4�<`�j�/�L�x�>�;jd��$���d���r#���+|�at�U>[+�j��E��6>f��}���jiv�C�نfYu9o�&�݇���w~z��-��L���h�u#4Dt�?;:����>G
p:��	xM<���3ۇ� J:D+�:9��1cp!�7�jj�vS����w|&Jx�Y_���j~M��$�_��:��D��>�k�~8��כQ�F�ـ�]�utQř��z���B�pB�m�~K�_�w/-
�lX�w���=�)0��Ra|�x=�!�`E�T%.8-^bʦ��Cl�C;��g�N�i�|�B�81��(^��ZNT%����
����1�Պ�K�Tzc�w/a�A�	�~��+qNk��Y��tRk�i�;.o*=��U���������� �����BZ���cO�������N��I���!'��;��6X
���l��f�5���]d�9�Xk��na�tI���R0�~z��ݔ�N$���/*�P$�̄�q~���v�[Z�|����~��(C)��3�M����\�#N������G�H�߶�2 �E���Ϩ�F����3:��������! ��2�C��Չn�Q�k��ު��(0w9oÆ�\�������l�@�%��I�D͇]W�N��22�с�d���`��CK�v�B�2!=��#Q����h��$O^w��"��߹CI!�j��.��hb�]`|��뤙Ո�ir&������xB����4�!K��w�sl��)����"R���}3U�(�V���\2Y�\��I<�¼Զ	%��È�B��w��r����Bi����������ø���z�^k=��y}**X�b8��z4qc�OI��u��~]d�(ƒF��uYHh=Lu��G�D�՗���єd��
=�rC W��VS����(�G�U�u�b���`hl� �b����{���.ɍ��w��S��5����O�H�VR_;���{��e���9"SH'�/�M��¯ҽ�bN?]�h�	c�K��WU�:|���j���k��*��de�[\v���u-}-$�ri��Ε��T��q̶����E����j�h{�f|TR!j��7x�c������X�f��7���4�V-��-��)�A'��oN�8���1q-�6FQ�9k�ٜ'ߩ��??���\0�a�-&�v���`���#��n�ju����m���z�#9�n*�r�MW��������� ���
�u �ڍ���y!� B��_�c�-MAW�MKݩ���[+�^aA�(�"8Vo��w@.�,*��g-0D�	A?jʋ�8y���}6�Jb*�S�-53t�C���);��j�q4uji[5�p;����-�g��t������騩H��꛴�ݧ���:��dH��,�u����$zD`U���<I���j\����PI�|���>��&<��XR�P�'Zu�9�q�B"qQ�Dv��K��b��FI��\fО_����#��i�#���vd�(�翮�߁��5��6$	{Cgs�����	y��L��t�7����$5��UM蝡� Q+��:�)��Nu.+��,�8�~&G�s2o��	C��Ȃ��o+�.ι�21z� ^VI�G���@R\�k?z$�v���z��ٞ?�X���U�Ð�m���ݽ��H�68l!�v�_4k�&/v ���߲��7���]��hJG�Ġ!�=EE�%��P�Fj�|a��	�!�?`%K�7�s�Z���(}�t��N��b��(�H�.���~U���a�˅�� ��l��m���w�-q��$�/7H��&�C��=GD'���X��E�(A�����Ђ��Y�?e 4xb�9�ő�gD!�G��η;�jv��F��ފf�bd��+����RdU�tM=�s� ��M.8p�N�����O��b �0���B66��(D�����c�?6�Ŗ&J�T��������f�[��X(W���L�t��I���ñ3���}h�:�+��Y�%y��^���2����0N�h_^��φ���S<"�d{�pS���7�[t9�c��=�ToCp����u[�u�5yVj��^Y�L6���萼9�N�`���""���7T"	�X����6��C���x`�[�In��zn�RD����Md��/��l����h�T��y�{8'�����b3�[�,�	eB������R�z�z߬��A�P��4�X���=�LP:5����u�����!�+��� ;ؙ�3�3Q���b'i��E��̸�
�~�;�HCc��=W�~},q��xٞ6,���ȼ����������
����>Oz�	��}F�J��Mc��ŪU^�tQu�\Z�y '����D$	{w��48ip��a ��a����{�gNs���R�^/<�Q|5qw�Q�O�
I
TB!l��D�ү�=�����܈|,��G����j��Z��;� �~O'���J�_ ����+�d�wQ7�R���*��2o��@ؐ
If�벨5@k%�hĿ��$h\��/�Bӊ�2�u�XȾ7Cf�Pg^6Ɂ�T��\,�
3�n�x��oZ�Q�b2�w�Ctzֱ�y�����N������}.�NG���GSĪFuH(�aTv2�,����>S$dz�?v!wF�����L�)a�?	g^$_�2���;���s�GK����f�s����$9���ׂ�v�|�TX����L�l}7�F�����q��_���>:r^��:��d�����Bm>�w?�$�G��ߝ6Y�!j���j�!���H�&���~�����R��R�"4H��`G@�rkfӛ�e���`ڋ8���,�D�;�rk��R�5��"����@ozA�Z�9���ցQ:����;��ʃ�X�آ{�n9�?V��~��m<�%3f{E��"�K�S�#알�h8f� [X0��P�Ս�yB�huʀ� �DM���L2��7�����ƺ��h��t4h��`/�B�61��e��>:���j��j�v��4q��0�ڷ�������Q�����#�I�:=;��}���k�����C�l�[��;h[�,�d؝�%N朇
�.4�3�(�U9>��?+��q`�O6O��lP�1D 7��X�5]��4�2n�t�������ߴ��嗘 An4v۱�q]������b�����U[Sӻ	�Ғ^g;�\�>���F$�L�!^貣�y�rKS�E<*��"/0�a��n��nzz��-G��E� K��)�*�l(/����2���nc+�T.U�/7��b�0��Z�U��	��M=�*�Q��E_�*)!G�:�
*E�?��E=�Z��[�1kT��}�μx����&V)M���z5TFQ�7��QԜL��۩;YrYa���θ-*�:�����rAD�\��0����!�m����cjZ\�[��r7��M��*�A�T����Mks��o(����z�HI88����|�'�NC_a^>�8l�2��9y��hSp0�Mg����b}Q��D�x;.z;ňng�N䳩���L�O�	cv΍�a�յјM�mv����Wo� *~���1g����n�������<^�����ke6Y/�l����FI)�ӆ�@����K�J��`�J<�,����u,F���a��� @��7��۾;��}�� ��<�8��z���;�ZǓڥ2�<%2S���t!��#�B��e�9
<.�/R�jG��!_=�c����9�o�S�&?�i.U>��%����j���'�f@�3����m��W�����F�&���9���g���\mB�5�7��?��L�Y
�?�B�7+�~2}A���"���I��
o6�]̃�f�/o6���j������~����4h <�%LM%�������	���44?� �����8�ɘ�GїC��Ms���x>�gyc👐�>��y��LI
>�����b��	�e�~�W�J�S\�}�+�fQl�Z2w��D�/ޡn�Z�\;?%Sj�!��*m��hlV��򽬑�A��Ϙ�϶���r��NΗ�e��A��;	�Z�N9��4鴚6��<���5�w����p4��ìF�L&2�x��qr�T��J��y:P���,�$(�^@,F^4�~Q�)�I|��J���{1aY�5�Py��p�y�j�k���S��)5u@���T�{�`Ț���+��������c
H����m�:����ܛdKs�׷ɟ�������ف��ƸZ'������Br��ЃZQQQ:������4a�����UK�iS%r[ɝ ��!�����)ӆ���퀭s��Y�U�ҩ]0�䳻}9D��(_:�ُq�{2e_�M"�N�B�/�#n$2�4VL��;�z��?p$�1}�{Z/��>�px��ڿ�z��������e�����Ύ�.�������[/�F>��p
�u]h*΄=X�\ �F��B����Tc�[��>�����Y�(�߇P�@G�� �  ׼�`)zce�UQH�l� =��$꟢vB^^L� ���=#8��RC�3�	P�W�|����|�!5)��P3�7W��Ь*����:Q���O��\�׍��#}2 ���R�k�>p����	��m�db׮�)����Ӡo.v[݆Sb�>M[��R�,��`�Ɛ.�B�(���S�q6p���0:$1'��X���������Py��v��!@��JY��@8�x�#Y�m�bF�WtT`�gl�������5��?Qb�^
���H��A���c5*���5�q\�HO�`�U;�PDo���f��?�����SƟȟ.�����LW4�k�}Y�z��Μ.	�Ӎe���*]�z|�/��L�7���ӎ)�f|�������O��]1lק��4���Lpl��|]ZٞՉ[H��h9^�u�(n/�R���\U��J�A�O2����D���*�{��z8E3� ���3uBS�^��bN&���;>��"�Q<=�!u����S��a�LtzQ� �iV壿�`OE�����%��=���?�W�lV פ�/��`Z�yzPf�Z����	�_ k)�ZrUϕ0�4��]1stE�(��큰<����0Q# 1��F��(�h�ia���D�����z�"ϨxlF�tI~��(ϟǀ�e��
D��W���ݬ�uf����-(��J�+璵�TI��Pl~�����S�&�N��4E�u3��� �q���h"+p�0F���kwӾ�^#��t nsO�����[(�k�s7�s/QFj��n�c�8���������Wf"a.��+2����������V����Q�����_.�� y|��=�ZK���LN;a��e�G�a����1v:'�4"��"=I7q�Ii�
|L�05��{n2m�Y�U0Y0����^�����F����j��$(���$�&�;X����v�|6��:�[�t�_V�p�?~�]�����5X<h5Ƣ,��aIE���!�LW�`�,�;p�i# ��嶥����Oi<ILmѴ�]��0D8����U����v�5��sUħ%�[��z��%�!@��F�~S������.�4�S�J�hi�G�u#Ƌ�+���} �_s�04���y�9Nl�Ia��e�s�[�C��O9rr����z�ez�xs�9��C���n��_7X0��h��v�">�����o���T`�s��n���%E��т�\��rWoa�vP�J��
�J�M+�i��y�����R������ջ�<��pu�,����`=��ٰT���Æ��c?����{éz+Z]Y/�ߤ����O��cF��av�w�����4����V��/���K����8"�L��֙�M��W5?#��V1y�>Dp�-��r"������䍎���y.�s�i�*�-.�`���@$)A����/_�	���)$�H�_٩���[�wF���vQ*�,��V���m�%M"�X�]bq��}�ξ�K�L`-?ÉX0W��������_9���������9yu����B6}w�'ro���Mty�<�x�Xw�N�s���r<���==b=�\jY�e��8�-��R�x@04��"�@+���rE��.�MZF�a��*)bD��٧z׹3^o�N�S[o֔
�����+��8�}!~�������ˉ�I�����I#`_=O�[��ֈ0O�M|�{��d��"h-E>eI���Vg�k߁�$��+_D��T蒳����d�,t����|@�[�jز�aE�R���b*�-�_7T8��28��/�âȞ�'5	ɹLbY��:��*���ۗ�N��8�8R6PSw��z�*��ui��ح8��._��Q��V�H�\'�����񆲶�wo��'�����������`���;�ӡ0l{� g\�M�	�5T��I�Vc�����,�2`k�a:�u�^�V�ö��>�w]�V[!�����9Ym2N�t����ި��!�?����Pʾ�؍���E*3���y�Β~)V#JNͼ��y���pcl�~�/- {����$ئ�o���ו�a$�A��G��	���F߮5��9�1�m���+D!%������S��6<a�����z��!�y�A-�zl�(���}��K���_�V��>�J�=��m�!�2
.A:�T� �zH,�6��q9P�X>ȱ�u�}5����?q�Ne�D��Կ�@�-��V�d˖Ccu:���z���r��b3G.�p\�3�@U��bl$Y;mm
V
�?fy����9�#g�:��J�v%���w�m�כ - �bSQym���qt��ͺ��wȽ�v�e���)��w�i�N\��!� �`eQ�˨P��aC�L��o���>,d�Ǳu8?ڹ,U��>�}�r`9D����Y�1�<��|���p�w&d�h��*�Mӱ�����h�����]�������[o�t9�W#k���\��n/6Z(w��d��n*s�����m����6�Jf�,m��!���?�u�mY�f����?��3��͝� �?	��|��.��8�3��!Lvo�7�#�Mz���Y:�e �D�����G1S�x����%�y�
�-{����	+��>��^�2#�xXG������-h�^ ��{�����e��d�2��[��>5�ժ�f�Z5w�hfs������������(��(�5Q_���D��Lǝ��3n7�]��bC"'�oG�\%�����B������]���t�

���A'��F���4�Vv��챡SJwnA�Ǥ�f��4��O�1�]$+n��e�ĝ��O�Al���K��*ӭ*�d�=�x9�3Η_'�lo�m�M�<��k��u�j�D�Y�V��;'VkÆOR9N���y����]5�G��2�Z�(�y7Ӝw.�:jP�ݯJW_W���D��?���4UV2�*/�_��o�'����r�T�38�/040�*��F=��l�ti��-sh��Sn�~�Ȏz�0�^i	�� az�_�����;@� �+�v�hdJ������0NK��/-fjd$�(�)V~�)_����v�Z�U��\L��ԯgy[�7��2ff��ʆ�eiE�\W_�=�010��Aq�8҈�SSU�5%�]�o�5X�C_�8�z5Yϗ��C�Ѱ�N��,�����99��G���H{{!����ꆤ�H�(.%�����?L�87�XX�:��|�>zz�l�@o�=���ɫ>��S��HP���H������]<��MMi\����YJI3mHeb*	PU5q���[�.C�e�Ɵ�z�oߢ�:�~;�����aC�I���aU��>�Emg��οJ$��.�w�u���w�D(��FNL��/tŞ��m�\\Z̈�J������3�����f|����+b<]��xO��9�'�kG�mVb�ԮFj|8&&�qr8�-
���~���U����#,�-~6��#-~a�q�>~E��"�^/C�R?�����M9
2�Y0[�u��H�uX`�@�����w���rS���d�r~�g$�f��@��*��b���٫�����&Q�	
vAA
�Ǳ���G1����٦��9�ȗ
#�.)��ƢL����`�y������^��A�4^g&�p] =OS�.�$T=��x��(H�HVk5�K�+9v��m�ϻk��.[�r��R��Z�K��G�B����C9?��OJ����+����Z�4ۯi��罯�$B6`.�%���Tp���E�A��Nr$%�s��vƷ����}=Z�Q��破td�V-8�B�,�v!y�;�z���8�h�_>�E�%e�kK,
�@��y��nX�����/�Sy�y��$ ��+����������#�����Og=2#���Vod����KC����
� ���"��ҭ �<_�|Z��5�R-���%���������rq���4���Y��G��/�=s��H".�a� !�=?�pT,��կ��'	Qd�.�x��U�Ɉ �D.�v�d���~rBve^2��\����n�Sw��8��y���Ͼ+�u\�2� �j�c۵a�{:O�}��x�� ���mkk���p;U���]C��Fot@e�e�nsu�������7p�x_�g�ي$+���0:TӨǁ�����!]x8����;^�� ��h�hp�&lz�c�M�`P`'�Z)%���<���(�'À����_B�ie:���#l�C�w��	�] o�UX3�M���4�������'l��k�o��9�^���؂)�N�k>�����������
yVg�|#!�����c ���'��Q9�_�� �xceM���m8p����yte�f�9�B��r�U]gM�V�P�p|�d��ϵ�,w9��G�!��t�x:{#�z����tW ����halLa���ךe��"~׃�7i{cK��żN�X2���F�?��3�?�	J_o�`���:���p��������;��)%纨��Ӽ�0˻I���x߮R�q&0�+�-���u�#!M,`����wݞ���$ߞ��O��=ؖ�M�F���QG�T44�ߜG��>���
�Ono�����&�_�/��S8ۓ�d��{�/�;��`��f،�0d��tC���û��a��΢1y|��Dg����!���z�}Ƨ������J�ڡ7�bkw�X�i ������<�U�`�uF���k���N}p�&�iխ���/׶6Y�u�����N�.5��\Jf��z�6Z���-sD�?XN��<�;�2�
@��0�;v��)�,d����\��}��Z6ƿ��`f�c<L�w?�x(۱���Dc�g��S׼bJ,��8X�l0Rwuuu�p��\�@'��/�קl�,D@2Mڤu�� uT@9�]���\��i���$��U%��q��`�3�,4`����s�V�ӆo$eY���I͓q2��2��Z���eDQ�+��.��L����g�t� ���0	��ɽ�%�x�.r~�{��+��EPV��1z>��߀S�-ߟu����0`/�7�J�kT��?<%ʐaY����(��y���ƞQZ�|{��m�dr�P��Fcu�A@���4w�q.��:��3�9�L7~�2������4ɽl�T��w��z���)&��ׁ;-tC�/|�15)C�G}�Q���L��(�)է���2�{���������E^�_ϒ
U����r��'8i2w3D���ػ�rjܣs&|�<�襰���Ce�T��_A��n)�븰��EQ��i��z��_������,g���C)4��
pGmݳ�6�i�.s<o�dO�W�8ޡ~X����� � 0Rɽ�6�\#o����j�ߣ�5��l��ɱ�����Y�¢�m���k�Rl��*_�] �g��nCK�#&�����=t0�}�I���.:�h��6���)AG���~�N��4���n���Y+t6��$���)��gw'��Ì�����.�7km��9�}�1�zߖ촟�m�|��.����p�'37�� �$�S��#j˺K45��V�feh��'�+���u�i��
�P]�y>{_i���{�n��.:���ľnu��q�NG�}�bַ����$Ib3��yI:�u��$�����
=��Rr�*<n7��@����갵̑Ϊ���qf��a�G7���S�7���~7��2w�1C�1��i��`���Lay#��9�&љM����
��F}��Z�LfgH��/o1�\���m�X���}��(Iy����z�sR���=�x�;���	���A
��Y�����ӛ���:_j��n}����,�a!�
�"��Y\ss��b�íP ��yQ#Y��ӋG�DLr�1�HՖ���'��Û��,cC�T�,�1�(%%y\1P���t~g������`��w�<;�-ɏ�%��I�%�4=�J<�s��#߭o�L���d��y��IDh���ap��#uց�ĝ���i�ն���0�҉�]���M'X��ɿg�I����]��o��|�<�A����g9�PV��84ۡi�����M�~��+����Q�r=�0���c��Y&y�(�z{����	�D˼�j��f�z����P��:�|�{K��P��@��2j{M�(�]<~����Y���ǔ8��d��9ጃH�%��p����'�������P���P��lo`���7r�T�|ns��[�ĩS=��ŋ��b��gm���e��v��Àh�'2z�Ϛ{�BCG;�����/2a���dB:\��i~��۽A�_�W�F[t�*��{^~��nl@L�)��U�k����$ Kp�!���K�"1jǦ� �c&�q3���P,��f�_�(��)���:�$G�q(k٤����h�ߩ����z��>� f�c�+�O+�J�P���Sov�h�I�p�I��RpEU@�1�Tӟ�%��bWR@�����4��w!��+l H�`�T�����J����~C}�3tjy5�iខo�Ƌ�X`R�U�5�Ҧ�)�CԉLn�<�y����}�l��i2��
�q��ij�qm��%��b��wc��eR�CJ���=��w�Jr�-T+�<�Z�%Z�-�7�8OȄ};N�w�$Db�HX�փ���I�m5�2�@_�(���(��¨��[tf>�#�/�X�<׼>����2�-��j��D'�������n5%���=�\	$� ,$涌L���hץ����H������L���C݁S��R�&m�����QhO�g���Gz]���:���fV�\�[c�E���D���%�F�ByF���KZ�"�����l>�������8�_8�u8]v�lc����Cl=�V�D�ʡ2���E�<��k� (�0�#��6���� ${�g�oq���F`L�M�.�M�����cO���l
������m���O�+�>M�ǨծD������g�G�b�7aI�����cY![�%Wd�X��$���,�Е���Lh���3�p�`|䶭����+R�iRT��	���ݞn�uϣ�F4>t�t21~z�z�<��,�^��E��8_<H\PC���焥!���% 78։8E�~_Y�C��|;�b�n��3��#�[#v�g�n��K���O��/&6�[�;�|�Ĩ�ڹ�E� ���V�\R�@���=�� �=�ԱSY�6�/^G��t���Lf�c"�(v����8��3��0��a�D�hZL�u���pwh��e�>A^ej^�������&�O�5��w`/t�����8����y�M��qі���7�gN;�`��k���3$���+�Km�K��[`j����� �@ 4 H��ʭHVj5R�3���a�d��̏l�ˎ�a*R��傦΍��[��4�_��A A�?Ɨ��, ^Rf`�)VI����E��E����;�:K��TA��Hu��[���.���;,��i)���Χ��e�����mhJwX����㾯�'��.�1��s��h�\�A��n�t��_'����I�e�zmm>��V��3�ZJv6+M�a����B�u���$�����{}c�����P�[v5]ʚ��� J��/�l�-�ӫ7`dJħj��vpX��f����i�<�;�B<Do����@��
`�S��(K�,h	��N��+5+6	��a�R �� ̼����ڎ�Sl��#�*�d���0��?!���0�L%ʱ�s��|��ٍ�ה��� ?k�޲#iI�0��N��d�d-��km6�>+62�����q��T*�CB�B�A;ME~E3��v�>R�Ӗ3h��GuI_�k�;~ �{��T{@�x�vsn�a���,�?>��XH3��Og	��["�<W�kU�l� �ߊ�n�ҠT	�e����W�瑐���J�g:�*�EK�hG��iKج�7���o�C���NP>-�"4d���u����\wW�Ñ3�Ed�J�Ƕ$[: iggO�O�� �7��a�H�S��8G�\3q�P5���6K)i5H	T�6�E!B���D�4��YVo2AK�	yi����O�OSTn+���v(�H����\|�R���Q��ą{j~���!��<N�e�6�TM9u2&�Y�-��Y���|������[��4/k$�|Gp��7��-8���-��7���8��a�2������Ř�8#	7��S��ݍӗ\&}�M	0�ܐqC���Q[A���u��#��%��hkť��Ԙ�P`�@.��ܐP� ���*
g� ���	��Pj���Sch�W���&����UӒ���J��4t��l���t� ��i��Xx�Ґ`M
rC�WW[-�>��j�f֌%A�l�����^VLBl2��B�i��8U������	�[S:B%�jd5�R������U����9A��ZB���s�x
A��j�Ѷ2i����#n�$ >�y"OZ�vLn�k��6lP6;�C!��Jڬ��[҆a?�k�*��5��#u}�}�!�@䘷6���Ax��i*� s
�h������8���]6�����4���ɟ/��O�h"�E�FS�cϔ#.^@u�m�5O���gdYO�E�P{,!ܜ�(HcHg�գz"��b:�p��z�Զ���DbhI,�6ۯ�(�V�f>��d��i�_�7uW5���e~됌�AR���[�!R�G��n�K��[[�!��Q�}X��%�q��t�!�#���.=SA�QhZ�u?��6_a�i�e	�m���$Ĝ�ܭ�0JӺ�g��ԙs��=�ܯt�*�i�6�F:u$\�X��>s�X�IdIJ+��?���vKҖA|��
��>�_iW��}v���%�n3Ys�S�Q5�$RH���qqW��2�]$0|�
�(����U$c����Ɗ��S��p�'�nL|T�_a�_x� u]�'�BFvL���Ev�;[�!9��������p�rv�ؒ���<�o���+���\縥_��_�m�`EL��MsJ�~��t�A�Z��". �fikb�^�#��5ߵ���&�WgH��@�����c��]_�얚�ǹ�B�h���!Ӌ���ժX%�Vvp=�3OK��tF�L���\����3���; h0&��C^�G,Sj�03K;�/S�	3�Zsu���[����?3J\NY�r/9%:����O��Ӯ:���_hkpi*|B���]E�8)���>�4W	����z���k��+鳦�&���o�T�Q1�R�Kʕ�N�Y7^"ͮO������g�e�a�"�жn�G�b+ȟ���PW�,b�*��_DW.Ů*�u��M�*�ބꨜ$e���*؀��`mcO�b�E�dK.�Ɨ��o����S6쯥)ԓ����Yߜ�Z�2���A�/�,�'��ƨxSXr�n�R)HG�o�����[0��i`�"6��4�N�V�N5���R��1�暨X�Sir=Phq�M���du �"9�~����^�}Kh���B7�cP�� � P/p��e!Q���ư�]�^�7*�m�~^I�(Υ}3�ҼF�Z�YÉP%GPSYC�Oy��×n�:��*�V�D�+IrXVC,Q�F�K%�Ȃm��ee��i����7c�o,��]�p�N���y	��,�	���=�j���}�*$��¾m�
��z^��; ͊��O��w�S^��>��;��by|���5�sʋ���z�Ƴ�B����^���#i@XK/����{��>(�Ypxp�4E��t�X+����lG\0��a���0�.eZ��ۇ��'5���(��R`e�_4EI&D���
�.�����꩟��%t[����^�B��N�j˦I)Z|Nxy���Ԝ3���
n7<�JJ?�?�ZS]}�l�^�,�V��3��@��O{�!�eᛔv���}�!�'�ؒ]��O��8��;���i�!՘V1k�gP<��~����}޽���L���r$����φ�m!n���*E��n/���tM<��Vz���*f<��ݧVIK���FT����F�g�Ғ�[pe��d�볣��v�Ju�U3��f������;Z��o���>�J�b�H&�h[���m�W�Oلa����H~�[�ݨp�Z�!PX����>qт@�VTcKIݜ?����K�|�;����fIq�/X{ľIC���@+AZ V��C��� N�;��~��w4��#T�����fQ.��nf�Y$�������l�M?
��cl��s�:z7�c�f?��oGY�&�Ż��b�B��2��e��ͳ����|����5����lF�������i����2 ���8>�*�É��#�k��|�]!�!Jš��u溙�DV�֛/�!M�ݞ~ge���2aN���g�[��׊���|�g��b]7K��BC���ulbnә"[��.��2�0��o{�	��'
� 
3r#,�F�ǲG�5i��a��_�Q��ܱ/��|����h���������v���F��YC��(�x���cѳN�U��:>m<�|�RN������|9�/��v�ݑhY6��>�\���>L7-j�sӨ�>�h:�*pt{����ϤEq�0��wƺ1�x���0Z�<�f�i�-u��E�R=�f��5��ּV�͹�ڢ��fk�ͳ�͚v�_�����0+0��C1"n�#��onc)Y��ɣ��f��i'�>wg�S���v����d���S�m�:>���n���Co�*��3֗����W���rɃ���R��$_3U��&}�W�����FxN����Y���a�i��2����V��@������G������ݻF�E}���@4g((�G��8��i�Í!���}�&�ot����|H��E�j�S\6ܗ�U�m�Z>�r�����G٨��]�&�uS��:˨���o� A$D��.�[Z�[`�DE��:���C��!���;�����y=k�Zg��g�}��ߴ-?y+5NB����<��4�Bj&����j����� ��,H�="%�C�������w�¾���sZ#��U�Ʃ�R��oN�c�S���|�X��d2�ic!v]!y{�{�^׈b�ɘ��ڪ��
Qp���WA)}w�jO�Rc�nE]���1%\�h��+�O�M-"�'F��C-�fF:~(��
��l.*G����*D}�@d��X+�(I�o6;m�+�BQ_����lM�F�-�mW����8����nW�:�hP��D�gB���P��
��D^#y����b:�۳�0E����I��ZȳO�un�.��is���jb��u�<td�O#	N����B'@�Ԃ����`߯}+��j'6�ډ��7<X}�7#�(T�9j������݁ڱ)��	��W1�HT��2�+����-O��.Y]���E���v$�~!�nt��=�sM(Ԓ��S���:*���-�n���H�h�^�VG����̕�$��uf�(d�Q:�G�*!�%�g�>�����a�aVNC]T��&���l#f�l��y5��b�%��f�c]��xBӳ-�-4O����k���[�Z��xG��D�����r Ecf����Y�SO�+�|��=�Rc�-u&N�Q���Vf��ZĽ�Nd{���g�;�u-����r�}�:;�����ۦ�U�o����F�S�)�\Bu��MsMݚزDk��d�:����&a�=W��K�S�s�e&���Xޘ]������N�2�S8��˘���Z1+���pV,$��6m��)�.�VL�ԭ�~Q�lZOk�!@�3�+q�����j�賮�3����EO�mF@�G��<@�
m,��}!���e7��ҍ�-X����X��ប�4�����פ_h�Z�Z��/�Gm�8X9�٘ ��m�D_ܩ�w=�>9u���n����b '�d�ɴ��.�~��)�M�$V�"���cqoo(����+5�(:����z�i�2%�;|���VU�E��4�����jO�4.W�iIi�����w�Dץl�r��d*J6O����>����١���&�9+�%�!(��hN|��Ʈ��\#�*�>t�l�P��������'
Y��������N^F}���/��
*�ꠝV�؀�0X���l�jm��d�[�y�!:�tp��$�8�&o_�0�xބ�Fx�s�u��.�y�:(<�c��79�f��YU�c�Q͉v�r�H���y��=�²��Q���u�K(�e|������z�Z��/]�o��.���t��� �H�[��|_�	� ��ù��OqZWf��O���\͟4;"�\F¬�(�2���(�ME_�x U�#�~SԎ�}$�n�3�c�w&��a�����Ŝ�6d[��j*�~C��Ϟg�Zy\B\Wټ��6_L��7��:��[aAw	J��N�:z!t.��qE74�/0��v�>$D���0��5{B� �Eu��+�
��L����|Q���A)�r��d��刮��	����>7s`X�HH,`���FyT�C,q��5>w���9�c ��^�s�k�Iڄ�&����"dqy�|w@1Gܧ	���#TM����뺤�ߨFr��^d:�}E��� 
�Ƅ'���m��V�\��*�<#y�|@)"i{yHR᧾A��QZ���n6��a�$a���m���[hچ77�L�Ls	�`G�(������Fs{>[�O;b\<"�9�ʠ��U/<�^$�O�Q�fuUYd�'_x�73���C!@�i��*f�$�/\:^����&��)�*��1t��T�x��6��b�$���p����Y���5�ܘFb�I"r���z�]�k�/+9��};��\��Vo�����-���74��jf�5��:�J��_��#0�E��%F�xX�tA���/�--��`��7¸4.�8,����+b��fϙ=6a���7N.��,��@&�:fYS�`����Z�O�݌�᦭��s�MZ���rnu^P���Z�����w�����;�]�.�t�X��[�O������1A�̫�Ԃ�(��Z�ۛ��Nّ��q@�s�
S��#۞A�	Y�4/�X�?<ݣ5�z�u?��/�Cv�No��X�����?h�?�c����;R?k2���)q�V+��I>�Fdt��Ɉ��1x.S�=Ox��*������̈́��5'���G!��r-z��]�eo����8+p����6�����$���q�����~��ۖ��%��}��/-c-���_de'x�~���Y�5k�W�k�!���i��������+^����l[��l��H���Y���;t��N0�a�~u:(��2��ʜAݳ)�چ�|��G���\��T�]v�f�툎x�A5%+\��<U��l?qd�=�����V�o�[L{ץ������-�>��[�G��bd�&W� '��Z(lpY=2\��;OF%���)���T�Ɖ��f9ۯwK�uiVͽ>x�"I�gW�LЌ�G$B��u-�Q�M�b}RHD�`Mi�X}�θ�������hl9�y�i�qk�9�D� �E���4��܀ܜn"�t(�gz�;:!�OF�h�?���{RY72�:��)R6�]�<h�8Wu O`��K���0��o#�a:?&��ˠ��i�m����Bʛ#��k�gq2�z��u�ˊ��O��H���~f��E���1i�G�q9\ǋ�Ow���jhm_K$s�����%=g�Ჷ5p�����x��������أ��>�u?�_t��^����r����krmi���� ]_ȉ�7�����k����w��YK3_8�e���ac�mF�r���r6��0<yZ��/7�/�ULy�7_7�]����Cې��8m���j�7h���Z�hn��'���ٚ�7v�0Ab�����]�/�n�{�h�c��Y-<VCe[��no�X�T�EK�����UQ�t9T�_�7n�����f"��SeeR~�;[^��/f�Q/M�AǍYAj1�~C�QoF��VY�n` ĵc��̨�8�2�,xѹ�sTL�skd����/Ӣ]�{��pfI`��^g�k�����;xP��PBiU��e��[M��A Z���m!�L�ۅ?^��9�N]#-��`���!eD����Ȫ_�8���~I�1�j\-��^�K��)0����u����O��hf�<��£��n:�K�,�>C���-ݠ�NF�Q�H��f�,�n�Y]�g���>~	[k*��}����q8��@ߚ��bſ�j�t:W�~T���ea���b"�U�y�w��}%�J��7^7msx��4��O�����*O�-0���}��^ݍq�s�w1����!�9Lq�r@U�B �����q�D�����܂�9P��_�\O{�<>��Ǜ���7�ʥF:֛W�m�V��S����!�zW��Q8�-h����s<��۹*�Z��d��-�6�%ǋN�H��&5X��Sc��+�}�q��P➌~�=�*Io���pL2�@�u�,��qj�e�xq����s�A��M�=s��2sFD����[��X���#t�����]Oe�r(!b^����s��2{�ԧ �E,�W�-�̽���ӎ����<�D���aH������e���f�����ס��<���g��`��+���e�*7�s뮤:M�b�}��_Kq�¡�^$�x�6��9E�Ýx�E�enUZ�jj5�7�E�X���B@�?B��r��L��a�������Z�槙?�[@��%?��D<U�1�#ñ��,�]��F�� G�������� ��ԩ�2x�e�ށ+�3b��BM-�p���j���ˤo���!!u��NH�X9�6��J�}�C���Bp�[/P��'Qʟs�9�����D��z�`�Ĵ�0���C�v����"��d������B�]0�Q(����6��~�llm�E��i��g�Ř~"��w��`�MKwN�L��O�VK������2O��]�$y.�{�ӣE�&�����)���U�i9�6��=�V�v�3/1:���eM��������h	DA������e�p�ks��7����'D�;F��I����p����5Qd�:9�%�K(bb���9���2���Wt\��mѴ f�:I�)�eh�`&����q9��ռ��YC�eIB*�w��vM�M�L!�����땬@3A��D�}�����&F'�ZH��ח�H��ҿ|�B�7f�����aU��,b����nMq�de���9� lA����O���Z(��D/s�\M�/�*���o0�oY9N<�:r�\��Ar��׀3rW�U1���7�-�-�����^ @G��%�� 8N%|3�=
�r�9����e-��+����l�z�˒���� ��6�Aw��E���n<Sb7���m��GQ��<	C�\ã� �sy��F*��l�)�8�f�Yh�s�D�ՒiK����b�|�q��www| H��U�|⽂�f�h�� 5ukUm6�S���^�@��f:�g:���{TU����g���͙⃋���И��n0C@�K㊎|��	7�N��N�:�
f�Y,�{hq�L���~y�7� [�4�>�h��S\�!�6n�c[Ӧ4^|�lJ�o-u�E;�5�Zp�ǫl'o5���h�r���m�"�_A$f��z&ܲ+���د?d�DK��(Ztm-�FD��Hg��|�o�+���tr<ă<~h5e@��ל��(ݛi�NN���w�w�lo�|KP���j�/]>�}>�?$8�͞���ׇ���,�V4�h �6�J��	�[l��{�M$ۛ^9Q��@_#p�U �n��G�]r���g�>�Q�or����j�\d�����-5`Ry3���<�2h��m��k���Ԫ�jK��i�cû�s��
���c�ۼ��q�Nz��'--c$��1Y��)-�mpϿ��~���OS7��o�K�n�Ѐ翈�Se�4^Z��q{���P3�)	��Y�#���z�6���.�E������ä�'v!?w3�81±���\�Y��Z#�`!U�`fn|�$����-��Nk�V�}M�K�+g�+��U#�Z�0^��2�ZH����.Ӿ^��W�s	�]��H��Ԣ���jU��柯5�M���#s˒��4%gd�Nx��_*��"j�����H�v�������"[QN��<�]d1���A^ɉ��]����~;���	)G��K!_�}����_ݠ��7:��=̀-���h��\ĭ'������4���^�	9� 96��(�@�Y-��_-��ü��f ��vv�S��^��%rw�x�t�6�k�5Y�B�jE����4c����.���Ѥ�M�g�IXv��}JІ&"�Y��D�_C��<Cʎ�e�kWL�}�#	8�|���󏍀�1/�*jz�?	?�G{�,�3#w��o�[h;�����X��t����������[���1RA,�v��ȾN P�dD�~�{CV1V�����\J7m��c7�i�a �i�4d��y�����W��8ע��7]{/��w�
��$`pqϨ$�H#V�aS0�f�)_ط'(#v�׉F� =�]�[9Ti������U]��\���T2�K���_`b���`q�X½�t���'��+<�KK_�@w� ���d�^�Q��Ia��>6���2R�؏���n^egv{c�[��7�X��u��
�}�tH��")�C"�ZZ��%�u̹�2���t�\$����'"$�pj\O�Fq���ǒ�@�Ȥ���?�E?�r��bI��A3O��)��i�R���8��@p#u��5�׉�N �pOj��ϡ�F�ztU�'m�	(�Xvpv��	J��D�m�H�(�{P^�BJ���_�d�N�� �k8��~hٙTKTeKz�q�N�˸N-�S��H�WQ����.��d��K�kUU��4�`��1���Y].����y[Y5�+�l�%m�8�zLsFL���3,��`���ء�$�����a��3p� �Y.U�b3Π��5y��ٴ��ZC"��s���r�k���(:_�k���$"�m��OV�֯�\�9Ɩv��cKj�ZM�?CS�o�v����S3yėDk;M�;����	@��(�BL�=��vJ�4u � P>�C1:�I�'}���?�*����_*0���1#_�od53���~!��]�jޑ�%Ĝh�l�nDL�z�~�Y|D�����Y�\9>�����M��������x/d�w�T�cJ�3+T�S'��G�m��H
y�\0�6�eI�T��+y�d��)��[��ۍ��q�.�FubV �g���P^�`���8�o�#��Zh�x���R���߳C�ia f�`>��!��ק�C1U�ᩛVh ��1�^=H.��e����:ܽ����n$PS��J��Ckf�N���*$w�S)W��1�0Wv�N'Mݰ�v��������/���"*=����r��[�I��#���&<����M�|k��c��C���|�}!��C����_��p���E;�&���w�'u~�P���W��>��ѽ�Ɉ�o&�ng����B�ٌ�+�e��������P��[fM˳�\�(,��i�� ��6��ڍ�0P춃e����&��6�9���}E3��;�˷��N�dB|��[Gu����AV"���E��1��àsZ�nڤ��t昣��;�z4�=2Q����!�;�G&��c�ҵy:��ˢ8UgZ0#8J��}�*���]������n����?�2���'*����וsKZ�ޝN��o����1��s�z�f�m�GH�G$s�21-��a����$wm���X�ߡ*�gJ䕾������T`eEc��?y�����s�4�<z>{tՐ]Kz�h�q��nC<��W$ffFv�T^���엖e�m�g�`�	� j�ͅ�bU˩�Y]��b*:��#V��Y�]�,��;���MQE�jV���j~�M,^K�Z�&-KťJ�x`���~-�9*�v _�E��^��'ȁږW��4{�9�08�����A6�a"��4�Y̓�!|���rP�汱x�O��P�c�w�x���������%:B���b�+��������4��/���A��}F=�����'��!Z(�����ɘw�+?}���-,h�&��A��[�i� ��Pd�T{��t.|�=�G炛�5��UX�E�p��/\������+%�����;�oE���)���
��ߎ���s�6����cz��P�:R�0��t�����7I2��?���)����3��U�s��b�}�%:rR|�SB��lA��^��a0C�ٟ�|��介Y8/m�;�WOL3���T�]ĳ��80�6X�QH}�y/�@[.��6ʾ�D	�k�j�vw�2�~�|t�R(���c��\\�����-`9W�Êi�)���~�A���N�Ye?�{�x&}���0�\?��ۗ�~��}1�+m���������ս%��ID�g��v5�ܩ�PCxe��öf���d�u�.f�C��LT��UD�T9����F��ou΢B{�N3�Fs���keee�b�����=�����'L��b��J4 ���9�-���8���#��[; ��Ci~ϵwf�n���=q<;�đB�+
]J#�o�2��g<��8������F�6jmӻ9=�}��:F�?6pS=~7�@i|�9ߜ'�S����w߻�a��aJ�ama��D%Ư�%�*��Ww�^+kfQAk��RG
F�$U�qW]�x��n�"q��]��M�O�4�t�����]��l���QeH��LAh�C6�@pQ���D\��B�"�*kG�56	��p��К�&{��N��`B�0�?T�F�L҅�[��j�̈́�Б�\J��<�[�*6I����%T���B����-�rP@[~�ys��a�*��ҭ���uI��H@B.���~�W����
XX��т�,�T3�pH�0��A�uG{4��Z��e~+�l:������HR);�Zu����t��@�ء������V��Ws�y��o�.!qI�./vIV�ߐ�h�tL���k���_aF|:������+��hᤓ�sg��JFG�S%��vK���5��?�7Ҽ�KM�S�6���Gޮ���oW2,BԚ�\P�!J�;Eq&�X8��۔ɱ-���8kk�� ɜ����V��cy��c��QE�Qn�[�v_��J�;�f���el`J������+�J'�Q���GC�k]��W%l�	�����ϟ�Fo��uޛ�_�Jg�8�
��������Rv��l����X��11Ύ�����c��y��̠l���'��)�����d?s��F%�����#<�K+���;eǵ�>DG�����W��D�������Y�3x��j��u�.�
H��H�-�����z�m��@+��Jr;u5UaU��;����k]�/���l8�:�@�B�GZ���?��O�_��%����f��V�UȆͲלA8]������m�xu�?ϗ���e��t�����e�e�nD��f�t ;���݋�=;]�����k�FM�sVD-�d�AN@� s2b��S�=[�s@��7cV!=��Z=�"��>�aLh�P�Q�-��]�5�&d`��.(���C-�ݸ.�x�E�F.µ�)cf����9���#�t���i#���zB��cN[�V٢�����*l��/�J)�z�C���^��=�Œ���uDY
���_i�"��w74ìd��_�[SRl�占����~n�"W���iN�#�ј�ʘ�]���St��,���ͽIL@��A�="�Ɠͽ�"ɱ�:Z��D,'���?��>����+B�"܏��m�k���'/fMݚ���v��At��,k� �BG�1Ι���Xq�\I����̫´Z2���@s�3;�bU�������:%�)sm�	��C%�����ˢ�fwϋ�H�������~�
�͌�x3�^�x'y��(N磫���F$FS�jw6�lG��>�#�t�jI�X��%���]��������+���� ��4�u�̗��;��@�딏s��	IjJ^z�O�$�H�Q��~���%�����;L��N��T��{w�7�Ո�N�T���Ͽ��'��z<����,��*�x���rR:y�bW\d��M�"^��ݥ���dBQ@D�$�O�Hӳ����g�8,9)��&9Мعӈ}�")�(0"sII�(+�*���m ���]>��v��^jb
@�x$MZ'�u@I��>�l�SfΥW��%5�����]��bH���+�����!d�)���{O�m�����l^�93�z�m�xg��x<��vY�Ja8D�JL�_s���1������U(BK�iR0{����y1\�dK Ċ�w4P߂x��K<����g/�Hk��o�� ����������`N���n���tLI�r9W:ƺ�x����(�c
{O
{丫�[/���\�Lq[bQ��J��_�{��>��WV;
ߝ)e3�p&��;��Z�B,5u��T�)��T�`0'+�5��!K|�E9ʅD�Gu�Ts>��ԡ�i{2!�c�Lq�E5�k�*��E<��}��0?̮T��E���ZPz2�{bLB1�Ԋ�}������z���ʠ�c�Ȝ��x����Z@���V/�&����'D=LSK�n�����g�������d2&؉&�l)*:��(R�!�m�.lh^h�+��O����.�ˑ�g?.E3�BF?���+�.����ƃ��r��_`�
���S�&�N�ǝ��x}�˵0���E��������
��7q�1Do�
!j�f�/
�0�y�˾>�]j8�R"��Z�gg��~�g�6���<�+m��׺�R.yE��@�3D�٬��[/����iJ��T��n�2qL���S<��>��C��q�h��Ң6�h�N���GDw��LK�>���nT���_���WOP��b��[�>o�}�j�Ԯzq�K�Y���Y�~)��!�N��`���-���be2�Z����`^�3���o�q��}13����3�xy��qo{�|HaO�8�:y�x��}ϻG���J�c>���o2ț�K�e:�L��A��Zb"u}�⯵��5�61�}�+�K\ �.��ݦ]6t\TU�᫾9����3� 7��H�nɶ�F�A�k����>�� u�G�kO�����[����2�Y6��~��4��R^J�OP�Ep�aT��Y< Q��g�i��W��xЎ�������S�%��;AKz�%���4&���gqW�G1���K�K'�AǬ��6�5��t��רO���
�g��Y��U��v�(h
 ��-��񀧆�����_?�6����;n0 ���-��>������Kw�2Jt��_���������;f�a���B<g��,ϒ��ɢ�y�Z�r����/��xW�����y<�i"�D"#�
��@��� [��\0���
[H����� Uy��,�2Q�̛��^')-�V3;GL��t,˼n��;���Jy,�I]�r���z��s���J��fg���G��o�S7!7�8�kƑ���Hk�AN?�� يG�5*\B)�3I`��aD@���g�����nl�NROeR��ʫ��dk.C!K���.NC��R��f<`ع8�<��m�(��	Y�\��I�{m���(�W�v��`����x���M��nߵa��yًx�@�n��@U����t:��G��Z���.6]�I17�&�]!5�ޝ.�;�yi�v6g:fnjlP�W�{�ku�q�q��E(�ث��Hׁ5Q�*7�-��R�xT���Ж�c��9��%�B����- ������C`�e��BS-�/g�P��<jd΃��6�owa,��a���~�,Rw�&�G̲X�gk]�o�3�Ff��v�5��N7r[j�ZRg8��{���Xz_����p=̃��|%�\��[ ��N�8c�>c��L�-XxV?U+AHBJ����^��E�h^���-�iX��s[a^�;�s%l��o��y5�O��;4�?�h�F;�HXcH����*s����{�Rf=R��j+CBV�y�k4��s��xy��P; �5�t<��x�s:�\����N*W/ɭ6<;;ItFV���K�-��쮰��E�Pm�#O��NK�:�o�]8����=�W�I�������'�|-:[�e��Qm� 
Ǥk��Z+@�y	��**�/|�R����$�9����N���l%��	š���n;|����>�DA���X#CZ+FL);�ZU>љ�2tz���/�!у�0I_����4���`s����sI��[9�w[ʌ��|o*�y�!�����|랢��1�K��jO����M	���-M#�^���E�����}nr�P���߰�P���"T�s��'�^�2�6�E�Z}��!�k�ڪ�t�ΩEE��["5T��I�I�7{����lY���t�e�é�
0h@�&y���5L�Bfwtu�(���r�d�L;(VD�� -Ҽ��x����8aA|g���w�w���ҕ�#��g|�3s�xĴ����l���O_D0�~���T�W��{�{�yn�7�VdZ���v���O��}`q���	��@�o�n?��Ȓ\��Ra���N�I�3W�u���p௳|���[K9�#J\��Gs>a. l����e8�+�,��{z�x�;&'����S��L�� 	���]���E3�mv�4}E/D�L�ŭ\q$-�ڷb6(f������8N8�x~Ĩ=g��9��ɣ����e��i�=>���-پM�L���5�f��b�1U�lZ����Q֋ҧ~�îW�������{Y��s)!�钆��%�q�R�E�E�>���t-����-�}ص	�5;�o%V�\�1H^�����y�����x��[UMu��[������%�t(�ku55�n��I �f[y���*����L��u�*)�JJ��Sv�\÷�4��������o� A�Yg#�צq^.���+�3}A,�����F�*e~�S2��Jz�b _�(��?�7%�@֭7$���W-� �Q�*|RE�0t�$��t S�@�Ϋ��޷"�?ر2�z�NV�y?��y�1��No}��08��k��L�\��ä���@yV0]&1]����L��O��7���l58�̕O!N�W|	��Y���)�kx1=O����'G�0��L?��C��[IW��2��[O�8Y�H}⛒HI"�O�E �m�P���fZ��|��gQ#�ܤW���bF���x�F���z�����"n r9l�����@
�ֱ�L�4U�{�B���+�Gc���J��[Ԝ�c�J���W�r��s�A)������ߐB��?�K:+��N�en-�!5�cP#>˿�XI'h�z���'�~$�{�)4P=���: ��\	��2����TP������.��.C�
#U�0����7�@�%^�� ���R.����J��Z�BAnQ��r��Yk�0k�j4/��Mj=�͓�(��
�lo��1��i��$ۺe�Z�������2�d�Ꜯ�
yz��7
�1~��d���6��S������W����iOo�0���W��j�F���'^a(�J�
R�>1� �F��������e�Cη�H���!���V��Z�*��k�Z��B��w!5"*i��.�q)W��9fG*�P��>w��II&Z���
�����7q��S�vH��@�j��������W��ֵ�NX(R=�Jp^�����LtU�P_dt{!��=�tG��,��OXe��E��앆NsJj�Z��}8��S�p�g/��b��.����74����p	z�tG-)�Z�W�y��i�$yl疕=晚�H���.����'�כU��p6�`���n�(]���_��͒b,��=�z�9���!�ׁ��&���3����h�_��G�XL��CQG���ϏM��gd��T���p[�O�r��"��DK� �yn��:�&��jLU�T��uvح`Rܣ���p"�b�7
+��3s�O�ˎY��pP��h��<�_���?wk�|��-�`��\��y��;�G�m|�ᙤU���8������u;[��WU����Y&+ ��S�IeN�x9�A��B���bU��)�u1�:1E�e5l6�u<�.�����8'����5qEһ�ᬩ��(��I�{{X�����S���K�7�Mۭ4�Z&�35˧�''������f��Y���R����<0_�j7�?\��6���x��9��E�h�*�c�O(��-4i�qy�IG����8�gs��)+>fS%�Iʑ�Iॺ�2�Y�?E5�i��P�C(��Ɲ��1����k�)$JJ���ӁP>-��gea
��dH����Md;½�6�q�ʃDv3�>�c.{�ǘx�������7�/-�7N�>=��U����?bYh=}Z6D+A��XV�B�^G�H>��C�u*'J�44����t�Z�������{&F8j���p(����a�����E�q��ۉ6���I�~2�n��\��7؎��1R�5X�m��xAi��d��^0�6�L�,d�{���N���Sǝ������7�.�"�	�^ ,������d��|�[����-���eS�����k/evo!�H�ܛ6��멼�Wo�s�,Mc���D���,� _�獜��KK7��&���DQ3�����b��Y,t>�i+>/�M��z[�Ij#�����$��<��p*������zH����J�
���w.�,�q�2�b�@||��=(����]R6��U�&�y,pz�<q��������*�b�:�� �(�	�����)��""t�k��:~�7$n ��,;FF(�y*��(,7�I,P�9��7qs��(�7�p�Xax%$�e�?��HG�D�ت�m^�rˑV����R�)*�q�_[CcdY���gF�&�ֹb�sg�%�cn*#����5r�qɿ��@w���i�Zm��1���li��w]D$����C�lՌN��2\c�4����w{���4*Az�S�Nޕ�S@���q�e�H�t�u$�x%��e|����z�_|� 4̍Ŭ��O3�y�*����s���)�2� �mx&J��)��{J)�B9S��Y@�ڐ�>Ea�1_/��s�_�^K"R��a.�D�3����M����KlG�������m������G����륢m�/�]-K���<U��͜�W*-e6�do88��n)۰ъP󱜊�����J�,巛甼]9t(Y=�$Ũ�)�9����yG�՜�G�'	h�bm=�<�j-6j�u�?꫁�p���w
f��Y|�U�����}���B=W��Nf|�ö�Dr����բFٛz�2=om�]�Ts�}~A���k@HHH�ss�������wDs?�3����]��T�t�d�8�-�ܚ������H��oͤ��>.�I
d����J̵��|(A3e��}y����煩�O&�
��9Hb�K��3�^�46�o<���\�m,/Ύj�ҭG#�9�']�?�,F�2M�
mD7��Y�jk`�7��#Z���I�Bt5��̞X���,���ֈ���˦Y���9I_M3����&�v��ٌ�ܜe��]n�i���Tm(�������������U�Z�	�����G���G�ᬧd]e�z�&W��c�n��;H��+�o�%Ϯf'G�s�JH�Wp��6��93O����n9���	��r��X�L��v����jXԴ��-��|�C��(Y�.R��>P�:��]p���z^_�w�_>&}3�2[�����Op�K��-���:�,�]D���&j#7nV�U��93�T{;����e�Eێ�o�ۏ�r4���f#�e�]��ⴣ�r�8�����W{�����j�WﻟWGQ�����������V}�w����9��_�x������K�B�L��S�Z��{gg��{{.3�E,�3�%c��Hc������[��떣^E�e�U�DC�^������g?-o�vޟU��Վq�����T�:��� �U�����d��ls����1wWwh��H��t��NV����>h�W[)�yM��!3_��<�Ncլ�<�]�p< �,���{|vR�����[P�}��ś��W{
4����h��7����g��'닦k�, ZŁs}����
�Nx���y4��F�j������_�t^i�)�����p�u����)�_����>�Of��e_�Ŋ�������O��)�^.9�j*I^k�Fbm3�ӭ�!��.:�K��];�l!~�%��h]F��<��z��~f��϶�}b(��x��0��i���\�t��_2��y�I�q��еy3��F&�\�Cy㊇���	�����ی�������rW^�Iw�0�o���T���e椧�c_�V�ng�&U��}g>=��jm��r�$,$�3�^��j���ʯQ����ɂ�D�x<�]��ˇF�?���?��
���F��ݺ�qWY��pz?t��F�C�P�KÂ��e�@7��Y��ѩŖ1�Yݑ#�fe�(�TQN����ݶ����u��u�jJ�/KO�a���A�˃�m	�H�+��~�,�EW�h�"�Gˠ��PN�+'!��D�t�Mo�5��e�M��$�L�[���vw�X�2ڗ�V!���t�q��K��Fͳ�If���dtZAydl�`���^H�׹�l�v}/��}���.C@N�^�x��x�!�����8�eb-��u��zvH}��#��d�^"��d�°3�ִ���?75Η�5Q���GF#�q��T�������M%�V��竭BϹ��0�;�~��x X�`����߶t#�)��I��u�yˀ#E�9҉=*ۦ��ϟ�?]!����H̥�yd��c��,o� �2oP��㗓j<����*�
�Q�w��m�?�Cݪ~��NFf�M�:��q�ʆ'�W&�2Ǉ���(��J����4�-�a��"�)���26�.��fCNY&��7D�d�ZWh�X�d.g���hM��y/�Tv޷L%{rߑ��!ȶ7&���$O��SS������I�����������9��gu��v�iCS��,����s���ِ&�]�}}\W;�D�(�����hR����b��{vs�ypͻ���v�,���NE�t {�������cd,�FA��;6�\J�_��\`]0]��n)�m,�<h��ܛ����ـUͷ�qW0�׆��/n�\=Jq�/���2H���(�4��+�5ޏ||�B3y��͒m�	mh[v�$k�9b�/�?~b��.ֈ�'U�i�0t�;�O�L����'fh�:�Cu�i5�~��Xm0?^ˡ�%I�F�3��1���ˠm�����A�Ifd�="�����!u�1�af%Q{l��(��ז����C\󀣞
�'�i��D���n�e�/Si��{����ta���Ȑl�{/όФ}���{������p�����"f� VUU���T�jԮݢ��j��1j��_��*5��n�ڵ��'��s����x�<�s���~�;ߌ?5<���+���f�Op	n��9����Cg���Aߓ�]L�X����OU�j�]�Qe�����u|�>qO�|���
X6���\��t�KL̢��;�s��;�P�k��T�5�c[�	�qrePR�W��e��~�����"XnR{ւ`��2�,��=6��M�H��-_��A���C��A$�z����%��W\sȳ	dl�/�Q���e�s��i�DD��Y��1
'�Q���|XiG�}li0�
`NŅ�~ތ����(b4��P�Ax�-�m�|@E�i�E�=�(+���c�udF�A�E�jg
w�T�N'2��Y���R��^��L�;Hկg3��'c�l	}��:��� �P� f*�U9��c�e��!�
��|.�j#���L@�߼n�{���=ʑC��@�[{?�j�c���:f��Ə�
�isn%ܜM�q�N�� n]f�bR����!=:�0i�]����;�������EK���y��7���1硏��-��) ZT��8�/��9꿌�g��P��O��fԜ�@X�����cHϩ��`�v�T5y�������z\������_S�nO������ ��[�Y"�f���x���4�㐈� I��R~����?�Mתע�k9'�*�C�0��cj�`
��b#�ixti)��~cs�ϐD�P��-��ʘZ��	����#��w@ O�Fd���؍���,�:���d�RH
-f�{3H%�O��Kx�'�N���h����>�W�G&�� �^�}a�0�14�&�1q!�G�W�b(k(�7���z~`U�9�o<0�l�Uo[~����)�O����h�!�ň�F_Z�=�� c�A���9}⣖�_�8 �qt	�#�&b*�����E����eٙy�����>�=!8hv�,��qt����>��a��Ȉ��O����.�ޘ�>Җ�PJLȒ�u[}!hv��dL�=���cD.K�*i,4/����S=���3�kc����8kK�����Y��.tOi�u"?0՝���g��u��@�:�+/��;}�t?���]wK���x�����+]�>�Lh��
�0&�`X�4ij!~I"灖 v(^T�T����07�B�Q%#�[a�����=��wK���R��t�$��ࢿ'��P�|
a9}�y� �^&�N(ס%N���j���������&z툜�t)1i}"3�W���������za���jqh �>aq�4��fdȈI�9�� ����L>����2zjG��=���	؈'�'���½;c%X|-�E��A��-�/I��#;�%։�fFGR�۬q,��S��.�G�^?Г�����p��[�z�0�Q���u�4�j�+Z�/m�hmp���������W1��[��8}�Y6��e��ۂձƖ�ү���� e�׼�"ȖpX��0T�ӱ-L R���Ij�����G,��<iBDH�Uz�굀8B���uvF��;h��ǅ�$���#n��
�x����lJ;d�p$P���b<6��(�By���������� �>Vm� �,�D �O����j>�8a�i�$�h��0%2�� �1�?�W.�x��Y��PO��I��d+�lr�-��ǥB����Gਿ%�J��xR�w5�꽷ߑ�j��O�?�����Hw�j�s�!�ѷ����	mn?��~GV�bYt6�E�;�T�¹��J�II�k���TDt�g����K8�5'�uU_C%����n����K�0�z�`�}\�uδP��R�N�&��*F�0�R^~�,L<�ҁ*t�s��aRXXY?㾐���O��<�y	�%�0qs
i����e<A5�ڑ����^:�R��r�E�`��"��O����?fݵ x��!�g/PSa@œ���� e>���_������T���f����Fd� ��ʹ�Mw�I�W���W�obX�a!�^��#eQBa1*(I�a�^孤S낓V���� Lh������:�_fFoO��	�ld*�&�:��Cs�siB��%��(n'M��2+�D��{i0Q�(���*j ��F9���.m��ֲe��5��]b���d}��'���m[��֯-q�ϷP��ۀ�{�r�pM���4jKd��bE�B�Lη�U�7���R�c`t����PZo��1��1���<���$2�PUX- �T2T]�Ǎ0Q�	9G{XB��l_jM�:9�J벦�f�ABe1w�C��D�#@�.�ИF1����}�P� ��PN�`L�v�^�@n�CM��~3&n3��q���w7`��D�h,�H=��T��UmC�hyc�<��Z�� PO�� y��ſ�`����ߝP���j1��Q�(ո��>K�|}��PP�!Gי���j�6d��[c��	8D�H�t�x��_h04�F�a'z���y���D��T9c�	��T��V�hIϯ��J����AM�$�"�'����bi��@T���09���q����]��m�:��2e�y�YSK�����z�5�8��HS�$�UT&�&��hY	�宽ST��Sקg&~~�g xA�i�p���@(�3�C
/��"�Zs�X{M�BHJ�~�*�yv���-	%�xGm�k�`��no�E	�^�+B��PX�@�.}��ށ���>Im"{�K��Š�z�H�� �ȪTE U��*��G'�ͷ���X�,r��\N]O�s�>M�����"��I}��2����@�L�3�Sv��-5Ɨ�b������93�$��ݮx$��5�zL�`��f]���U�e=Ԭޓ�)i=��7��D�"fW�-�9���r��I�Ny6��F�ٱ��=��ߝ�9u9�˪���k������׎?�ßG�,����o�s-o��*aٮ?}`�� ����*�{�c(Gua��i �g����^�%�r��GK���!� �J���/JW�U�%�� `�@����@�Z�ρ>�h@�m� gm��j�J`n��ѫ%��R�q1`��%������^�a�$��&������l{�3k�K(=�d
5$�o�,������LyK���u�
��w_a���F����(�������o���t�����zD��=���Jl��$,�0ACֈ�:�D8�D#Q�$�+�"yr��6փFTN���W����i�2�\M��xX�@��>qQ�>ʕ���qQ-���A(_�H��d��T&�o��������ΌX�[3װ?���6�p��$ɵ�~�K���~�9C�#��'���/��d����:e;ru��X::�Q�8���a�9��g��6VJ
�s�%�}��^]����J�=��5��XǦ��?6eBU%G|�cβ֍��6�e}�?%�K(�+=/��]�����������C~����QA��d�s���t*������p���^�gO��Uw���Y�,FP��^�`�b}�,S
�A�����¨�*�i_y6�o�V�ӂ^_��m	��$6�L0��s5��.Zw~B�G�w��(<��2�>$��0E$�w\>^�I}�M@���i�>���Uw��cfg�"���y$W�ܿ�����<�*K�����G�� F_H��<_?�jg�׎�b.���ktM���Aq�u��r���.sp��QL��UYAλ��zek�P٤�?��r���/������g ~���L��������"��`�Q�V�)��#J�`1l���L��S�Ә�~?QD��Hn7w��@P�)2Ƅ��3b�G4��7�u,���Y�5d%�1#ͣ}1�2�����V����^&ӢO�h�g쾑&c��g�]k���'����j=a|={A�'�%�zz�}���?|�)ژ�	�P��[�0۵ �៭*q�S�Bi��k��M�0�/��%� ;�%6�P�Q=k=m��$�cc��2���(ė�ă}���z%yͣ�����m�r���t�B $������\Ț��8�_����/��@��!,�N�?�ΥG����ѫ�T�jV��􉯼9�*_LcG2T&4�\}�5�
�;�Vzdi�,�l��,ԟE>���.q��Nl����W�|�k�;c�=������^�����Ϫ�Bg�VbU���R+?5\����I�����>O+��z
��q��o���7��)XS2;Y	_90���)xݍ�I������!I]k�'(^��d���FX��aw���Ŷ	}����5۴߅�������k�]���?��\���GU��&�3���N&�j�����$�#~��)��o���U?U*�ԕ��}Ń|��,'��8Kyke�q�ٓ�u-�~1=����}����ZNĿt���I/��9ª5p����i��Q�r-�C�`����`��^�Tvw��2�.y����5_CVz�Ś��=��j�'����5g���?H��q[/)-]�r5*ۻj��xN`�_[8�e�f�B �)�V�-��M�+���s�jb?�'3�la~��\{�.�c��d)��û�_s��re���|l������x
K�p���Wy�.tc8�o��n.�犭�X������<�ސ���ggg;��y8��D���Z	�:[�>�l;��Kr [����'$�~� sR+Ҷ1-��)L�д���'��&�h�_k:�w%a�;+HC��l�LFR*����Z��iָ~��i�����ݣ��������2�PA�QD���<��!�Ξ�������y�VZ�^(�X�L9������2����Q7˺�;����#��MϮ>����n����$�	��w��֟������LΗ�l9k����:���K,��\��L�A��z������f���M���#A�Ñ[A�u�c#e��ݗ~�ήa�5��v�N�?���|R����v���<0��4A�����z�ӌ�醶�p[���myoL���+�B|NW��~�Ů���Ǒ�fjq(��^0v؛<n[�{x�Y߷5���}_l�k�kx���J�E���cf�L&�����X9�^~��q�ߋ����x�4p�_�$6i���	߂��
\�z"��8� =�i+��?�d�)e�QN��F�[3��?���O�x����iO^����J���c�Tz"�ݑ�>�[!��KQ[S5Ŏ�qBn��9���.K��g7>�$��XE�կ��g��r�U��?w5(��Ҹ�aj�~��|ن�D��m�`o|fj�ɨ���w!iҤ.��=��?c��6���[���\�=>i�3�^dt��~�����
���l9.����M�4�-��	>/�Ti�0�l0�]vr"x�d���U��'/,�'΃��e�-��k*;��s����AAH�^�CC#��z�g"	%���]m���{-���b������0�*|��4�aͫp1�����|��B��f�Xh`Ž0���н.*�J|2Gȅ]���2�OB�^�=�r2a��͝$STQ�:��4�Y%�Q��M�/�)�2��Յ��K]юch5M��5Z���Ƨ<�0a@��M�{5/^3�S�p��e:|ק�L���}4ב���p*�);Y�=�9ŏH� .R�آN4��r�	�"���lw}�J�������C٩�������Zف���;�gMT���owƋ��eťNFP��'Jl�]S�i�������WQug���WnO_�x�JvyVo"p�a�9V�t��6�OF5\�ew)������1�*�C�����m/��R��è�uRr���l��^UzBAA��Ϟ=c�74N,�@q��1މ�ѱ)�%T�~?�LzU�S��(�%�o��<O%�W����p�M��=��敢��p��ݰ�o{���wj6pEH��+P==����IhVZ���}�C�
f@���R���a�t��ngۓB[8�T';��&����,x������J�ē�2Jh���_�	��M��͹X�x��b����/���Zy�\��!Wn��R�Ľ���7����Ј`u6g�\�[p�T>�D�ݙ��|a^��1����l�r����.��HХU�IG����C�ʪ�k�=5!-��T���� ��������(���Qn�E�N����_���s�6��C#j�t���?��8���==EsÒ�h���F�O���K��M�}LO�f]U��=R��P��D�4s`%^��߿š�0��'��Ɣ�7�(E�eH*������O!��ۋ��,1�(����b�_�#f4���{���S4{�}jS1�!b7f��V�Z2XB*}m�
o++*�W�p��BpV���������e(�Vθ�Yg	����� e�[Oۣ`C�x|۴x�,~~��1��Y]ͫ���qB`�����G|�j94MXU!n;e�]�Q�DGY��G)%樃�ݜ+��ZuEQ��@�lu�\����U�' x($DEcW1�ĭ�]��n9����Wʮ��&:yt�Z�81A�!W���k��<J
�'s+�GJ��� �'"�J\�ݔ�cB�ek��B�������~��Qڤ�|U��С4�߲�_-���0Iª߬�P�Э�Q�qc��n��~�ƦB4�D�˲�)B��0Rt7} '�0pps��`��1�����5�5��.k�Ǥ�M����i"����]��D)I��g��ɦ���a���_***>��\�;�(i�̱�JvF�l}�
���Rb��\�\�`kIXQ�-Z���j�����D�����?F�OW?��{��B�I�ͅo�c�:;�hlw�{�4�E�*A�7��h53�9��C�)}�
6V�>گ�%��.3-��#�_l�J�k��t�@��0��F�B�����:��g`8���y�4���XD�����znyc#l��=�xO_W�6_;�},����f˹��5>^���(AԾ�� ^rz f�acNbYy�/��X�8B��j�c�9��3�{�8
ടu�~؏���l|��"t(��*�a#Kv%e��y/`H2Fa�G�J/S��Z�Rq~�2%g|D�E�������u�^��~��퓲i��)~[�����k->)�C_�|�~;)_x;��ޞ����+vо˓:�G���T1!+ן�%c�� ��r4 P���
]�Z��4��|�s����C�Hy��8��i�F���Rc���]� �E��+a��;ʣL�I{V��M��`Qad:�;)��mU�b"{vs���5�2�5t\���$ݥ&�X�v$����Nh�ڲ`Ns�p���C9u5#MF]�j�ҭ����V0F]M���A�����N�7j�&p���81p:z�٩7bMS��Pѯ�����s��(�w[������,��ۍ%����`U+�;��E��s�@!
�E�7B�����Db.]�)݉ a`\ɃB74��b����~�84���~t�wgj�#ҕ�8#�B ����&���A"����3\c8	sRXroL���j�D˔;��q�]�Z��K ז��;��B��,!��y�)�C���m�
�փg�*v���WcS�V>�d��V��m��b�Y�ܝ��ݾ覲%$���	���wS?�Y9m\uF��y������~K�:�-w�s5;+�������<j�j�]� ����Z�����SM�� 795�#��P&�r�����2'��!���:���A�U{�T.gD�&�J�GR�N�s'I-)�3��g<����:����(kJ'������K�y��g�aT��%�h��ϑ��%�>Xv�-��cX��m��t��3zq,8�df���YK�TJurd�+�/�+ʑ��E�u��K�D�Uȷ�|#h��)0۔��|������G���v���V�Te�|�m��`���ꖋ찑�[O�Q%q��d�w�]�-�	��d�� �<^fm:**�L�ir�Ws\��t����L�$�2��s��[<�4�h:�P^�D.J[=�U]D�>ʺ��O@�!�/���kL����B_���{�G�������zu-�E�w谔(��.�[N0���5z���ea��l��˪�S�7� �S����� �wc�U�A�7##��Օ �����5��~3�d�[�<U�"���~%hs�"�b���p}��25���
6�wu�|��cLl)g\��6�'!�Z���s>�C�<����_��=]������&)��E�ss��6���f?+o��9��d��;&
"p��S�UA�ʠ���P�&�!NG��d��(�q+ ���j���Ét
��oЂ����������:	Y��=q&	�2T\bBE����Sߑ����SP)�
�2�)��� �	�^	��8F��G���1����}L�e]֮�q{��*�>L���@��퍷�S{��AyBL�Ttf?�<-`������P�s���æ �-�U�g�7,Kb��X�\�#���T���w��sSb#P�����v�?r��I���矿x���;�B��lԠ�m�+��m'�E�]��=F�skkYAH�H�R �Syd����Ȩ�R������:?�{�^�7�u�F�����6D#��I*�>A����"~ԨHN+�o����lhF�ʋ�S;D_�����0��dѸgw����1H�Kʝ��/>Y��ib�$A�L?�:o�2~[���X��D�����%c�Ϸ~	�nW}�ֶ����$�a�s�ғ�چI&*�Q���K�۩@���		�S\�P0V�!�
g3�#�
��+��m�Zc�y�3��,���z�']K��5��K�K��r_Wi�z�1(%��R��e����]A��^z�Ue��IբI�$(GR���qVq���$�%�է��M�׾t^醎*���2hE�a��E�x4220���_r�joN~�0R4�[:Q��Y���
�ʻ��EE��� �XH5�|�����夺|ƹ��8<�g�����/՜���f��8���˫��8��7#�f5Qfwt�V�Q^��E�����}vHy��a��Q�O0�15���x����W�|�D-��\N���x!��N���*ݫ�`���7{��N"���ݬ�	�).�!lWOf�d�p��u�-:T�m �h������8�F@��.(a�B�Q��r��?�ޙ�Ӊ�
�<`F�3�m_�Aʼ���^e���͕����.�ޯ�[��Z��m4��~������ �
�VnM/T������Wf��~ǵK�����n�5顲vBH6R<�F�?ى(��x6;U�&Oa�Z@��JZr�-��[��}�d(lH)�lw���slȮ�)�8�H��>4�(wvұ�W^��IϚ�Z SRߣ�,�'���B���*�#�dQ:v�9WSO�ZY�#Od�ߐ1�7 ¼���;����H�d@����e�ՉR�w���I��>��p���@�3�pf4������	��0��H��Y�u=�ݥ�{�t��H-]�>DG$a56�GU?�O���<4o�#��u���]�B���}��6�b��&JKKu�j���)�K؎Rk�}�؝�٥�)�J8>IY�+���Q�R�T�b�%�Z���_�@ǘRn��Y�#Z�Z�DJ�Y�˲b��R�3�W��K�;�����Q�H����w00�Սy�#�k�K����%��P�{���t���/ؾ�.Pײ�Mh����@�rӼd�z��������>\�J]4�J��fڲ���`hTI�I���7ʞ����w�,���麲��K����P$'�9�Y��q�~=��E�)/�äv��ʦ{�}������˗/��(#���]�١��z *��3h1NO�1�I�E�ޢ�͗�z�;a�?�y��λ�O��Y'9��l�����떡cU�R).�F��ݳ��߸\?�)ZW��~�i�u�F�����/߬�|{s������%)�� �s�[卵�g})��56�3j�j�jB�C�����kW�г[g��vH�k�גn䐰6K�#x���YC��W��8vAYk_���&�Z[����t��>�D��Y���2�j�1�O)�����kT2�IG��a$;�:���h��rHW�"���P�
�����y!59����~�5Bip�WWCiU.�Ͳ~k���$����z�s��� �=�M�����f��'�|����Nv�R[���[��eZ��1cg��Ն�����E���˹���I�4��Jt��z�-��ƨ��`(���?n��ڪ�M����oM��/�?��k�S�t~I9xxCR��^Te���a��<������H#I֘�B+x����|37��cZ�wE����å�3'��cV�0��TE��>�Mw�I~ll���ёwޯ�M۸�t͈+��ϗ'�p¼Xc���r���\�I��o���Q�U��1V�׉j�D�ό�5j�Qrq囋�1'�m^��>��8_C(iЏ�s�PUs�|N��lS�]�̿�ý�g56Ւ�5_���4��o��7OqR`����0�s9�j&�����Օ������|Za��L/`=�L�sˁ�,�&R�t����p�� �|S��#�~Pk�u�t�������pf�Ȁ������c���a��l�k��J0g[1��l�(臭������2~��N��xO�ۜ:@��-�T���ymm-_��� ~�QN�Ę����L�4<���/{S��i�>�SX��Q�bf<��I�S�I:�x~��$l7���5$�m�[�H|#}���Q�t[^[�q��M���	a��#y�i�MR���8
z���p�ڪ�.یl�`�0yY#۫��M׀:��Y�d-�-]�P�x���D��ʞs��N��ɫN��aGn��_]��wn���j��tlV��&�_� I�r������M$;��������d�q�p�����j?��ٝ�E�Kh����^�	��53���'�����7��<�﮳N֝�'i����S�Fҕ�a3_���%T��}�~ф����ϡIC%h�|�3L?nl�%s�?4�y���P������������6��$�ۋ/Z��y	�KS�4���k���F4�
o�;W!��ڒ�)e�ŗΒw?M�9l�{�#KJ� �8{ڼ�o,���;e�q��մ����1�L����+mkr��m�"))���pŠ��?^�cae���L�ܩ�n<q����l�S��9���Ԩ.��m%��jtG����H��P���~<��m$s�%NbB��ź��&*T�L��-�������<�윜/��^R����(������2�������yIɟ&)�̫�s'l�|��q2}mm���������.���--�'�o^;��5�k������p�v��n����'w�`�Əu�¡�h�0�������䯹�m���S�Ӭ��|����٩�V@�啳��z:	�죐�/��{��R[忉���=|��J�q�|��pJ�������;���}��-B��[��6�_���ݖ����Hn�[`�QH��0x	��QS�BT=��_PK   �cWh��~� ˴ /   images/ab527b7f-4192-4732-8642-2eb32cc47bdd.png��S�a�����+�����S4�ww	-Z����n�%H��<x����s����;k�%_�;����o�\�j
x���(((xJ��Z((��>�/�~32�AA������P�����p��w�FA��JN�� �~F��=��S��PrE-�xƬ�AA��R�K����;*44�5�3���Dr.��I��^�W��ߑ�O��Z� OO� ��q��eO�2�'5
��[��2�������-~�.(/?��1��$�8>EED��_���>�#�+N���bb$��0P�e5��A$��MO�(Q4�_��oP	6�L}��v�g|(Q�w<�0����u��=��!�^2n�_<�7C��u=M_�j�?A��>��(��	zI�/*�v�.8�^�uh���σ�0��Ze�_�	�y���3Ӱ�l���\0_�ρ��n����.Q,:�#a�[�� ?0�(̼o�B����κ��F_��vD��ojԭ�PI?0�j���^;0�{�WP�k2����]!@V6�+ѣ^���:7�Gi�ϐ��ǘ[��f�Wz��5~��z=J��|+�e�Ȥ��5t�YɠD �ƙF#�<\��[�ܒV���>�r1;ŠbX�zY)��Ӻv�la�nŹ�'��3�l�_P��J7� `�^�[E�|��w%#���P����IM�Q<m�p�ASG�u�iJ/�Cࢌk�p�:秼����Je���s�3q-�x7���Kti�w_�pPi
?�;�3�ǋ�d��l
U���E[{/���ō���[ՍT�c��4��	u����0�xS��������3maDH�kP&�0�X(�����,� ��:���k��8Ή=�|%* Oj�L��U�A7c-�h��{J,�ω�����^b7� L�PH/t�������n�{���L�-�W�SCkFY��R'�A�1_X�Y�c��>!ylq^�[���K�����	�Ƀ��]�]F/�[�6R����<�)opI	c�����>hL#L�MkO����tgX��~�tb�!��ajz��q���&���0�F����&�r�"�R�b�\VŪ�j���<�B�y�"G�3�V?��4�����伂�2��|4�, ���4ec�JZ��\�i^�~*�C��fϩ$;̤�=�;gb�h��
�;J�N_Ä`�Ø��4��\�E��r�Z%��oJeu��XI�,:,|,+ZE5�umظ���z��A2�_�s34����c~$�K~�t�4J<4�c�=u�ʣ�A咍�5��g��cl7'���b��).��)�^�E��mmFyF�a���F��i�1�zָ��(�(���A������~��r 	�yx�|�����}����x�y������f+U��&poq����x���r�����W+�Me��$��M���9e�F:���d+Rb9%9������3��+͛x���H4��m��R�#^>.6.95�k<�H�H#�%ܨoq6���ې��q�9~�hn��ڲn�pa��,��iX��A�7:�>R�/4�e�c�9}_��i�ꇅ��{��&�&"��Ì��=a�h�͎[�+�|������|��a��q�&Q5jL��i�k)���H�(����hu�h����!�AyO�+� �i�">�8t��1<�ٹ�]�3�_^ݵ���V׻M;�mYei���r�R�!�};4��1pT�dv�{l���pg3d5�ꂢ�`@,�����Z� �E����Ӏ}�]��j$�yf=`!j�&�)�P�)H�mY�M�ى��Й,j����x��QhY�R�g��A���]?k�^^�M�%�:����umx����n�����a�B��D����h�Q���@�8>���7����ry+��'5�Wv�-�e��a+�٧$�$�rC� ���E�XZ��J�ØyGwC���?� � ��A�.#8�a���e/���}�0�����Xn��{�X��'��|��.�>�Gu}{�Z���( s$M�Z�Z	�(�S���د(�7Z0_y�`�{f��>��n��r�������|��=��e��(gtQ��[���b;^ʜ��N��Ǯ������\�A�Q��ņ��v��Tc3�_~{�9!������Ŕ.���������?���z����A�ڌag������s*�9fXF���֢n�����h<v��}b��U?��x��ZjhVki�l��������
Чny�8���Z�H�S�gy�X��1�=|6|�Y]n�h-�i��m2e�e�Y�_f\b��,�[pi޼�JfI��*'��C0��~*1�W�����{��TH H��kK�����|\�Wm���Go[�u+�.����/'hGޜ���.�Q�Ȱ��6��+7�0��yy˽Wn�>[}\X]^4x�>qޕ�-��TLvL���E��c,cg)-)ՉRLK�+F����ےr���U�H����p==�<r�	�p4��<�>�9�\�zaz����X�NU7qo�8c=p8�;�B��A�c{̈́��٪�.�^�|�5Fp׻�N��@�⊐o{[A[��X�Յh��[�( 8��D�,Z,���P��{��?���쀂�E���7
�4f�8 ͜d�]�����D��N�?׭��i<>�C�<^Ϧ&�i��\�_�NA-]�:f�ڟ�7ۛ~��`B�& �oJoN���J�!@�!��ˮ�F'�
�d���s�&�s��21���H�$	��	�Ҏg�0�g�c�ў����9/mQ.s�h�i>k������'[?Ma����Ǐ�0{�v��*���p����$Hs/�x�8{,y��I�[مby�v�i�p�����$+��gz��<�d����A�y|�v�����lD�lĪm�����:�I̦���qL�N�Ǜ1=���5��#������ݕ �UN�Uv�U�k0[r�Q��������B�F�����ʴ�G�&�ܠ+W$6V�u��lm��*)\F����{��UR��yy�f����^xjJ
'��X�X�ˌbu�i�u;�j�tS�)=_�	�E�E���j��͏�dW+��4��o�uVCű�\�����[�?�o� TTTGZ�Q�Mͤ�-��嶍�����U�u!797���ȰY��ɸ̦y�X!����r&�����Z�J'�aQ/������v�BWߟ�S�\o�r�u=���'%%��S����� ˫�T�**�%gg� ����՜Um]��ng+[ے��:������o�V!���҂�ۮ�	��[�.��Fو�<�!?�g��T��Ҷ�r֎���������/.O��(//W���)^\Z�B"�������5I~�\�50�E-�[1.(Q����)�!��attT��j^���m��:�.7��K(��L3o`�%���v����p�ԥW_~٭-ߟy��do_^Z�~vv6����=����vy{;S�w�E�"ߏ��[���k[뒓���v���y�<�� +�����ťE�8r���=���@�B�[����!�[o^���'_��Ԅ��h��##�� e���,G�z#��p� #�5�H$R�o�-�G@�[��
v#�	�<�L�Nt@�A;W�㒺�O�����֔^��5�TuP�I�R��S�F�J����6���F�,�?�S_�F��U��=��ۤ$�?�rpp�����m��k+))�Ww�7: ���`gm<Z�Z�̾t�9�����̊�V��p��;gg�j0r���@,$y�	7!5�����k3�v
�
>=�����^u�就^����Ƽ��W~8X��3�B���S�$\�A�u�#?�ՉIIK�����΍�]+(
-UU.J�x�G���p�a�V��8������;8:B9�s�mđ�T=�C����S�ݽxGB	�vg~e�5���i0`B
���H��N�������;��3�Y�f|l*��\�9�5�*�"j�zY:Y @��E�0�o�0A��y��HV66�W�G�Uͫg1c�K��`���N���;5'������.~	�!�G�w��k���L��n$�NRb������q�f���d���ʤ�M�48���?=i=�I�	�U�GQ��2`��z?��i�� 9*dw���7� �"j;��Я=A�'rӱ�q�>yU6777S����XV��\O:[�`�����t�F����{�F%o���L��%$�ׯ���Hj�u��镰y�o%5��̨�rj*gڄ��m�CB�ϙ�n��k��A������7��G-���˼�gNN������o���e��K ��V��p�U�����2p~��#��=S����k�,�YpL�x���.��Y`K�@���,�_��Oj����s�[��G� ��S���7�M60�S ��t	�:��?���2�am`tt/}G$ӡ�R�������Ow{mmF���p��U(�y/6�����%,-%Ij��ݯ�[�+�g��k���1[
:9)�	��d��Ŵ�4ņVXb���s���ܞ~�΃j�߇cA�Q�/��������1�t���*+?���zP4�M2��ueA��U]]N���F:Lt;��vov��@3"� ����t��?������N�P�Mj��3R�izy��&��C�4M�=CcAG����Y��oB����Y�����]����a�њ�zO	�]���Qte��2�D''ޢ��{��3���5�g�g�י�9|l�����TUvD�hG\%��'�:���|1�?�?���[a�	8��tj�KPC΄�m�?�$é|w;�.Eh\셞!O=	<wMq���Uz֎;elA��%k=�[r�x�q�E����^A{��E7�O�����e����	z�ֵՃ~����(�n�~��p-���6�9��²&��s���ggS18�LK��k�޳k<���ErZr}�6%;Ư>��g^�� �T���	�Dܞ�;ϳy���<7C�~�J*�f�6c!S�ty��Y���fv��Qo�{����?\�]:�it�yhj8X/��e�k����h���&+a"�"8��JR��A;;6�2�1Z+�[�.�_c��6ϲ��:�Z�$�F�Ϣv564dlp�Mg�B~g:l��܎�|��w1,6+�+�+���D�6מk�T���t@��#�%j�W��z�Ңpe%�T���e�e�8���٨�l3G���B?���,������s2�T������J�Q=+����A���(���1{�@5���\��33v�ȵ���i�&FK�l,��&�"��1M����4w�K��k·����`��g4�{	2�+��j��VI�pXU%��[�D{�ȑ�8�ENj����,���t���W)�M�V�x�;�����A'ydZkF���mF�|�'<='�
���H	2'���~엕pT�G8  ���\b~��jyx�� b��鑔��W½^R���䀹h�c��}�qR釬�{1�j9�򲅄�q���%�����J�6���/x����a�/K�>K���~��!ə �ŋ��],':�"��tшZ���7���Yܑ�L�U�S*��j�mT�@�\�F����"�kz�c��Io=��VM4n3^�xﯯ3���|��J
J=;d�8ە������s��z��E��ƍ���'�� ��3�B�������k�Op����@s���Iy_�<�y�k���?�
�~/�<EQ��V����ЩdTbN���Nø\t��a,_�B?���C`11�f���Р\��2�G����9�`}&�+�c"����Ұ	���?/R��㿳Ǒ���/���6:�O5!zuHw�v����E��b/���&r���f���ԱD�Fd�%zY¨�4Y�.�	)��@�����0�����'�mq��C(�z�RX�B��n��^�0W�5SHd@e����o���8�H��.2f+�4ئ��w���[#b>��w��P]X IU�b�&�{����x�*'�}c.�Df��kg	��S�U����cMW�	���NT��!Jk��q�a�x����9a�����t�w3���R�"�(��.��/�׼��;g8���h��U�m�}P$n��T:�������7�|���E}��#p���NCq*��V�Y�+�ue���	�:�pf޻���͝�]y��̊`"���nv���)�����O��Q4��<���bp���a��q;����8����e���5票O W�����t�:�t1�z�ۿ�i)��	L��'��-��QW˞���B:�;�,�%�>���lr���Q\~��jn�)}��nR5uH�[`#&�!�X|c_����X��/�H�撂����ȗ�$D>�
2������Q��>��c�p��V�y��� �n�&��
��c��/�c �c��n(����x^��急�:�����k��P7,�֠�u�}K�=�%y�"��Y�����&�P���j��Խ��z��NYJ��3j�Y#-}}��H����%���V�?>v�^�;�q��������~���s�yV۶�0,��*���5��0���"	�a����~!]�zwט�������fأ	`����rĚ�/*���Ў���"���'4|Z��,��P�����tJ��.��fA�6Ӫ�?����@�oZrɼL��lق�}|YrX��R��e��SP�x�W6�",l�[�2��9T�i�v,&�CG�M�k��t��ȂH{J8�p��| ��pV����$��=�e�+��(��nN�q-X��c{����L��.�Ay2�x|������1�r�b���l��-'j��:*L�ݭ�G�� �.(h6���k��s�����]s��_j$�"��@����+`��~?�7�V�=�����c{gh����Ջ�И���j��������7��c�� l_
V�"|+ʂ�&�"�r
r��a�b(	x�=i�p�]���b�q���ZY�E���n<�Sۼ�E���x\:�i���(JL<�FW\Abs��j�A�l_SF�Ņڏ��t�>?�yt����"rQU/�G|4��6I:������q���$�g<�k�9T�vB�c�L��Uu=�n����r��&j��e�O�(���F��v�������nQ��2�` N���v��RG�����؍K|+ܓ�̐
��h��Q`;Njb/�p��S~]��T3�%[Ȳ_���Y��z�	!W�H����j	F��$�\�����_�����u42r%������1��9ph���`\�G�G0<'�D6�qGF����yq �?���o�� �S�����Qc�t:�@�}����F��L�=6���6�sC�[�O��A�C8:uֲn]b�[�l��)�c�<`[/Ae�^�@1�,�H?����?�����̻A���:8�ְyJ%z57��3����#���D�����ݷح�S�M��1䵁�+�9�6��E�ܾ,3j�>kN��d���H��ݘT�:�S�4O���3�X-;0�%L@���j��eKpjw���}��ڈ��[�6�5��@��:�u~������O���;����ų�jɠ��]�6��4��mzn�z�|��9���Jʀ���)"B�0�؀B ���j*
���~���|��EMj��\����*"",�Z�jޤ�xs��r�*eߪ���P���i���s˄��ْ��(O���ӿc��^Xt�?#�*��Ơ���	�;�]�Z������sh�E�)յb�c�0��]+���ZԲɚ,�v����ٙʏFu�����sa��J,�����J�>���U݋��#���7$�+aWA`�� ��Ԧ����7/�0�*�޼��~)����l2]ƺ�}�BVJ��3+��T�0�B��	RdԱ	����o����g��``P����_G��a��s�	�N�a.=���dpV���GT(3��k�'A���Tb�8Ӣe_d�C�|�0(�'d���OuǙ�9���u(ϩ��FHyFQWcc�s.NT�_��c�b3.�M-;#����`F�S�k_���Yܰ�A�P)�l-�Ϟ��;�ω�D}��X�(�^7�$��	�7�mU�]�'�E��x|[����UZ�L$D�_�����[;ˊ�eC��|�x��t�}������c�G6�,��t�֫GIe�v2�p?f=��E'��.{���J��HjQ�6p�����^����\+����%��YBE�������>�c;�g��z4Sd�>�B�������2L��,�Nk�0C���v��@H���S�[�f���7Wu����r������ " *v�8 X��4o�߈�p��z���86l�#��!�k�rD丳d�+��b7�i3�חa�U��lv>+�9��-^��l�L�`&�IBR��g杔IdJ�g5ˌg�hN��5*��!�6p�9/�B�\���J/����b�=��J�ֵ��ߠ�#4_���l��Ռބa �p5�0�W�~��/�W���ƃP�),vg6�Q�º�r�->���s���ARX�d��+�N�f����媢��1rmme:��7��S��{����|�b���}��ߺ��1��o4f�1�a�Т]0���ڿ]��.O��~������XAwK0Nһ�b�U�a�i���p,��g?C���>�i�#���W2�R��*������������B"���#�yC:�-e��������EO�/P�[1��큑aeC�>"=��Lb��L]���HJ��f�Czט�Z����!T�҃��ԇ��+c�T�	����Uv��+�Px��e4�I{u���:������z��r&�:�Z3j���Q�e�H�r�9{��ѫE����5�f�����F�/\.b�A����H�����������I��U��Ӧ,���`C+��rcd�1�H����)vM�ݝ�Q{�)�9���Q��g�f]�ʦ3Q{��6DY�%V�G��Ԑ��	�F�Պ2#�N㩞.Sod����ߏjJƦf��i��YG��?6k�Z���
ӛ�Q)�y���m��oP�<)�;,�`�ܗ�M���s��3��kX_9�N�ڈ�`:oB"1�Ԟ&���0�έ����zd���LWq��+��`#�O�+��S�Yʄ�/5's®�k��?�=�&+���B����)�.�N�6���mJ�с������l''�֯I ��R�4��X��4x�^;�WźETGGx� X� u`�uM�C���~����ʕ�N�An���?�p��I
�P"�^��1SMР��>錂hn�IP�<��
_�dV���s*��e>�v��Rr�槧egB�j�̪���Z r�&�9��u�3�n���|t�.���c���a롌���Ob�xGo;�PǼ�n������7���Z]q���NK3'�|L���f_���c;�q��Q�<�Zr���-��`��x�M����`���h� ��(��"��Mݟ���W��]Gp�y^.�>�-���+jB���m��
�4ט���w��C}�����],�wP�y�~�&_��f���F,������9ʢ�.��Z���Q��yy�\�!"�w]��x�ݪ~I&���7ث0X08�{��{ ��e�	�QfS�M�̺~�/0���H�A�^�����5��з�l{� �5;՘tͩ�?�Kz��
����0WC����\�$����V8�B��O����I���q!����5������,�˫���)�;���/���GQ�߼q�~�����/[6'�Y[/,2�a.1r�o����5�O�M���6���9#4������3����g_T<�é��usff�<������cؽQ�.}�{P4�'��n~ڨ4��"Ee��J'������ג�Z#zQa��%�W���f١#�E��c:w�� e����-/��P�|'U�R�V����-
�ю�i�`��ݧ �@ɗ]��K�!�J5����u"n�.�)��Ku�#D!;~,ɧ�Wm1���N�I\9�X4ϗHD3읯��Ϯ���վb3�گ�%r�.�ɩ{�
36��o����%i/�:��X���j�O���K�*tή����
=���J��bV�r1�:X>�͠k[ncS��o)�*6B[!F������j`��UsEΝ��^�k��%��K���mv9�]�p�`aD��􋯖��Yf��Lʐ�	1ۜ�R�
��n����7�����_;��]���qcۡľ���ld:�Gn�ڏ�L���*��-��L�,$>�z���6i��Q�9���Ik"ʥ���ĜY߅JWĲ)1�;�-�N�s琞+�Y��D�AH|���m���V��]۳�G}f+w����a�ۀea��Q9�����Q!8+��^��nZU��!՘�v�v�c&��iٴh��rYz؄�<Ɔ��z�0K�O�t�;�חQ���F��Q�� �h��*��vg 0���ʊ����^�}^�\����-?T3Y��#P^h둿>KQA�UP�$u^��l�5']X���R�n��Bh &+e�g��/���]V��]��0|oA��C�O=r�۔���LNGjh�>����ӯ���6�	�T������utu�G�('r:�5֜O�ak箞���`��\�H܁0��`��>"��]��\!���T`n�&1���z�a�Q�k��Y���,;��w&�U��a�x6..
����$��S��뗨�LBD(VE�s����vn��XB�\;�3��E�0���Ma�eC*�$�6���
E�@��@7���R�֧���Q��D<���1�^'�@�Ӥ�J��˭��U��a��R!��8��?m�,��5wM�tzYA�3ѠJқٚˍ?C ��CH����	��G-�7��
�	K�s��4y#Rk��(�@a[Q�ش�C೯��C K�8�UL���2����Lm_��`X���CP�����]����+q�BH���ܢ_��U�E�\�������4T��i�����+��`�D�g��`��
�&R ^�I���x��\���Ҟ$�� �fy�A[Y,؛�	!�� ���$��O�OC:7���+�r���P�0*_}�^�$`P�3��@f�q��� e��=`�$U��YP�VA�kzC�|�1;\1UۍE�����~�7~�+L���p+E�+���E��luq�J�d�d���C��bw�CA���$�m��bqe�kl�Қ����Ǎ����n��p:�ג�p��AӞŋ돫"�l*B��g~C�������,�Ŝ�l�`wk2�Y�����puȌ�M��T���5-_.:��lIO�Eu9�T%����v�ϧ�8�^d6"���.�;��-9����ؚ�*�(��7J�K"�sH�����?H~>�3o��{��M% 8����:���}"�2Z=����+۱츀��&o��JQW���y C�dZ�+�yޅ���̞�@���Aj&k��(4l�Z�f��?־I�I|��LB��������ǣۘ� $(dkR!DK_����6ׯ��l����{_�n�@��F��<߳��I�j*�*|��ʏi9�Ӥ[Z=!&�pu�z�~�Bݽ
py:^�:�^�l��p��|����x�<o��9��mnn�7(�뱲Ga|���s�끝����s��q;���4���R2q���[!���*;�,3#��Tune��g��fr������A�_���ѹ��Yh(��$��4��}8���?�~Ǟ��%���J����(a���ٲ�6]��[�D���*��|�_��o�?�(� ��"�'�Uʦы��I��<�����VS�x-�"qE����F��祓��&�x���fq�E^����������!���F��L��<vA���ë�fj���q�DxSxKԧ�����F�c>���sV���CU���O�n�W�#���y��&�_��v�I9�-s�i��d��~�L������a󨹑/�;<x���4f8���g2Z]��PQVi#���+�������HNT>�!����UxC�m��11Geq��2�m��|׾��ʟ�9_�]-��WT?F5m�*/��(Ks�	��NPi��i�̄kF��<k�F����!|�	���ޓ4�m�u�Z��;a��v�?��wwݸ2KQ���vG��w(a�g�c�.�Q���֙$�K��j�o�G`�D^��/V>pu�l@�n������XjҤ����"1#t^��6�)�U�\1�J	 *&��y�J|�	��������&,��p#�*���jM:��Li��5/��|� �`�AkB�>{E�����i��A�|+`7�u>��;�����]�����3���<R�{.���"�����_R^W�?j
9�5�1#�|��
Ba���Q�y��{�B�`���zn�Բ�2��6S����偞�q�G`�k�a{�x+�;)U޽ 7�Ӥ��rnf�h55z�As̔��jF�j�����rJ0$S�-�;���$F��)p�0�}Ça�S=�F*��Q�'K�9�Q��:2����-�h�g@�ba��e�\����.�m��y6������lJ�x���y!/?�1)�|�ik���q��=����BM�|��>f�#��|J>����9'��0�����lD��������5�~����H�~��;	���@�Xp�l�����������P�a�њ�R�j���Ն�3�@�*��jc
j���GO�΄�GГP�$'`ߓ���B�^d���[�`��G�d���oe�pJ���~N��"�/"olѩ�`�]�{�aY�|�\�~"X&�!���|'�)8��Ž�X��.��b?0�����A�Y&�a45ME�϶TH0m�=N��N��H�,:��)��㸱nr���A���|t�āJJ�7�53;�����Rbr=��3>�ei/c�X��Rl��/���fꉫ�����Л�s]Ͼ��3?�M�4�Y�Z!9n���Q�6h>)1��e�v�hY)y.6�:n����y'�C��꫚F9#����`o�RdW��[�b��+�9�D⥔(�J�j�'U������7����b���ɩ��Ѱ�]�`��h[m��r��;V��~��$�h���0%#�
<�ݍ?�X8�����ϋ�_l#I��j}RY����*�@Y���sI��<��j9e�Β��v9�Z9�����jQ$���G���7���
��yC����䚁���L����'M_%{{_{�(qG��-�I J��A�$d�f�O�3I�.�Q��%f����R�oN%Z?|cD���B�)�d���1��a|<�IKJ9j����Y��T�d�˘��*3",�K�jt����v�g�Y����Al3v�""`"������PS2-���"k�Œ��_�w!��ʢ��(9�I�>��,�IV�ϣ-x ��L1�����W�wǐ�#א�dH�#�z�8���?�XU��Ι����jvf��{O�fn[�Ԑ���ú��	��kǚǃ�0��yK�r �������,����o�i}�4���c+�Ed�u�?!���\�J$�V,���2������k���EH��v�+�r����J�D�g�m��z��ar�k�p+s1�g��f7��ƞ-����Z���H M���z��ӽ�O�[�ۆ��eeR�'��j����#W��,��5��Pd|/���5��X�16�c��O�������9�nR磓7���_��%x�C��X҃V�Sц����"[�p�i�:�U��N)����H>rm��r���1¬���r�Õ����ͦ���AKtO�|��c"Z� ���39�� �
Wrbw���X�����I���dk��4_�1�	�/r6��� '?�z�eo�?ˡg������I�&������+�j}ˎ%�K�+��e/^�p�I�kP��Ot�<�' ��_<H��<��&���q�L\���A����@���۽���o�)T����	��$|��x��k�V���%�9[��E�\�_����"l�mhT/ne7�J�Ô	'��/[��Լ>0�t�2#���L��� tu���u"�$Py>5Àv�>��_�{�:A7�D��*���&z��z��L�*��/3��B��0ݫ�S�Ip�O�i�4���oAV"r�G�5�,mO�w��{}p����w�7I5��y�U������C�6�?f�����R�o��j�U@��Uy�p�#�PYP�ᇏg8���Y��bWR4Q�?�.���K�m�C��܏��:�Q٩2O&=��.k�멊'Z�)��U�ɰi������ו8\����c#@WyE��D�!g��p��:t�Ū���,��\�a���E1aT��NJL�����2���w����6OO���VvV;j1`۶��ne*�[�0虈q����hF�+T���]).:fTωx)���Y����2�1�ȴ�i�?�O�z/#��5b���A��҈�^���@q3����K�1�wܷw"��9��q��3\�yJ��;^qsC��n��18�	�~{cH3�Z��H-J>�p�S+�_5%��7��D�s�ļ��)��ݹ��\;�� �"IǗ{�Ȩ�V�Z��-E������-$���Α�B>ϫ�7�z�Fd"?#�z(�y����������#K�t�W~=M���7��N�t��ۧ�{�uV{焌qO穝�]�� Pi�ٓq�ʪ� 	��1Ӟ  ��A�:��J}�}=���>`�mv{-8'�E&
���+�o6�Դ���k���.jL��_�^۬y��=?{C]Gm�.A�DH�0J�z��9}���u�V��E;�N��:��^��NHHi>1��������$e�НB�N���z���`��g"jy͍$��-�ң�8�e)8i�s�*U�ظ�h �1��Z�����w�7��3��\�1�0���k!�J6z���$n«8B�V���`��3~�61�ๅ�*��Po2�1grz����%�c��������X��C�K�А�oS߶`F�0C]�л�y��m��Gߘ�%��&�Y�4dd����Y'���9�������T�����(��u�KX�P�j�����[F���q'I�Fo*�y�qӮI���#�L(~���_����_V���a��?��2#L�Q��z5ep�6�$N�lᐊ�i��j�������Jgl]��2���M���s���2�g?Z�p�Y�Ys�VV�0hÐ89��/�X�0 ��Ř�M�媰C�.�<��Nh}��!}ݩ�)��Ue�!J�1�ߐL!����=B�y�11����-��9�fQul#����3��֏�j�=ù��^�U?O9 ��녯:��w62��ʒQ9R~��Z�I<~;��=��lMT7,��\/po�Tvo�I)��u�wȪ}��s����,��O�=�!�����-����ͧ1��D��yWk�a��B����#<�%�f!Ō��($':��+��z.-Vi��:���广�5�s��o�H�-��0Σ���价�PLOhE�D��|��|,J��8�[�';�@F�.1"ķ���<��q+X��Թ�;���e�Z�:f��c9��ω�%��r����/Y���c#�\l|�/
( 2��rov){_�9z�L���DJq\��4d�)3'vG�.�±d_6��;��/�s�Jc7�+s9��5�r�e@���la���/M,i���P�Y��^x�*PIn�+�{/�}����d�&ps���$��D�-���I� S��z����Uk6�������dB��C}��o�ީM>���	�lQ�� ө�g5@z�IZ�L���N�a	�q�	O��
���c�8�/�|C�L}z�թ�L���S�x����@Dk 4Y���	4��@��朣����O��=JK�Svm��Ǐ�#�9��n�v����LZ���������9�Ee6�#���%�c��� >+�`޵�k��U�g����Bz+���f��Є�/i�	|���F��=;��Nd]U�}�
�lF�(��`�A�A_a�V�{I�S�U]9-�HӶS�mGŜzcwT��c��wG�Ǩ�|L'䖺!�Xߗg3Ay���eV�U`���D��"��VQ��#d��M��Ô�-�:3���ߦyw����A>/�T�n`�#�t�|� ��WC���`������z[Ρ(Ω-o���l:9�X�����T�L�ra~��7����Qp9kvH��.������H&}�p�Z��V�4f��W�����3Hd�&22�R�.��M�q�Ae����6C�Nc�]?��ݯ�^�W`���*c��!�;´�k�+R�?�U�Y/�>a��	$�h>�h@oZt��fA����l�Y���,�K0�����	��'�M9�����������Xww�nv�]����2��J�4��%�������Yq�Y����� =@¿���̑�)b=��kwhɚ���r�ޗ�X�-Ky�j��z�(���{���|���:���|��_j��Es���[�kH���Nx�e-˙��	h��L#���u<i�S.��]T�Y*Q��R�Ғr��߰)<U��Fu�a�3@��� 7�6�(����O������ȼNH����ږ*Rn�xC}�=��b�4�����c�%���Sx��%������r��K,%XBYHq~j��
紛g�����s-Ґ��Z��i�
S�V��+�0��h�=����ڮ����B.�q����NZ����1>��T��k�т�%(�.�����SY�)���|�%O�BLF7�'��S�RyY���D����eY�����3��g#S������Y���W�	�N�R(��`�2n��λ���}��W�O�r��@
�*�[�%�7��;st0>�Lt{:��8҉6G�hp\P�8?�ٙsF�y��{�������>������Ê	�ޡ��ex��ș�o|���e8��=B��f���|΋kG����S�s>+}��GF��B���3a����}�y�^=M��lE%I9z��s�(v�6̂�>���~+I5�[D��9��Z�w�&W͛7#�M���K�`��:.w�����f������((0���p�^=t��-�u�@p����V�����R˖�L�74I��lQ%��q�a�GJq�MM�(�"��&L�� �,�5���%̒�A���*�X�t�&�M7�Լ�ꑣR#G�HUVU����9j�$1k�@i#̬���]��J�ƅ(B��G�'.�9���h�ŀg �@b�Oz��V�癔/�Р�I���$N�/>��e� oE$��}¹u--/�Q��Ŋ�y���O�\}N�A���_9��Ru����� }�}%j��pQ�H=�ZB_���%G]u�Ug���[G}`Fs��(��PR�� �2�Y��<MW�!��sP�f��;E4e똯5��m����:�c��N)�p����殮1�9�� z]���s2��:e!xp 0�u�߬� ,&(��B�M(s������[1s��Wk�|��Z叙��d<���T�u5��-����ܗJ��:I��#��.��:Y��/:���^��%d�Z����xȥ
�cm�0�rXR�R��+�P-��
�+�l�7��J� jkW�x��=�ޛzv��5��8Vˋ^j�edd�(OB@ن͒�:l)�j��1\��ͫ'�·�7JO׃�.�j��6y��F:G2
2�-�l� v�gp�hm�'\��	P��C�8�}&��!�0a����e奖��s�!�&�� ��>���;DB&�ur���ӽٹe�X$�n�O������3^� h��9�90z� pLE\�r{��&# �������������|$븛o��?���!>O��o��S��isܕ�߰)����kZH;�oCo1Ӽ�uf��\���}��Ï8���ö�R�K��QT;(������]���7��@	+��~�7:����Z�{�DE���Z�z�˯�2��}�q�i�.R+�˵�-����@�� �g��$G�,pl��"2�a�(��E�"c�Mk`� �oy=�vY��&32d��k-�2�,L5A�/�Z��3�^zk{sjΜ9����K<\������py����$��;f���ɡ��m�@�L<C"\R4�38L,B�k�ȑ*���A?Z8K��9��cǎ1�z�J�m�B^;C���ue����js�A��40ꕿf��¤� �,W�t��f�V�l�;�H��V_��F
���"��ύ����$V9�>��sJ4�u�`����'�42���:�Xxc�O��Z:f�a�Ʊ1��~Gy[HN�|�������e˖�16�1������?��/�;������;�߇ª0�Q�Is�%�̣�7�}̖���{�	����*d��̼�T����'��Ŗ��+L��}�U�&L�A�Ƕ�so��-O��/�9��� ����g�K�5%3I��3��ǽ�mnl�W���Δ� mo5TN>�3��{>���uL.���OkH ���l�I��An.c��57S.G�/�j_��ύ-���-_�aH�%y+y�塷�5e655�@�P.`�<�2�C�  $��W=��9J�\$��y�R,�,���lmoUY۰Դi�M!�﯅n�VSh��j�s����e���\���� _`b��!@i2 Q�쇒�4i<�F]� Q���!�dD��D��?j����7��$�1�	=zUJ4�P��8�6�CcF\��8!Bh's��Ŧ�I=T)�"��L�����Μr�ĒlT^¡I� G�I��\)�ul��$�@$E-�ڃA�I`Q
Jl0sd���Z""�� ��< ����(��^]w¥�^v�u�_?�T�<J��(E�4�-���D��Rta�Z�@s�A	J��E�l�֕W����/|�P׻�m��v����U�TY�2����^u�g�#=4J	^o:H��"�:˺J��/�r'
���:��r̼��Q�o��p�q�|��l��񈽇�$�^:�t����z`��;#*�VJ����"�;��Ӕ��ZS#[����B�")� ��G8Cee�|QX&NL�?>5~�xS�b`��@+�T�_�͸qʋO������|�*)uC
��O�*��I(!�ҥ�R��a қ�A&�d��J4E�t��w�B\G�����4h��U���fysGI1Z��m����r\�e��@E1b�V<��p�B��bpc�`���oI5'݇� �n�#�(�K $�K��/2���\� R�{�<�G� C� *:�B	7���a��;V��ݑ`��!�1�:�{���9+^�^��C]-��}�W2e�E��de	M���]~������m�8�%���FmԬy��y�^N��g����_�Ee��^8��֍)濐Ӿ��]�Y;�����Hn%�u��q�^��9i��7�,��N��S���H��>�v�<�~�q]��_�h��ٳ7_�K��ɟ}yҤ�w@���9��)��Rg�E�{h}0��ZKI45���H���8)U--P�V�!����%�<�KDch!��)T=��N)��f��v�K������m�4ܚ��(ecy�3��~!�Q� ۰�,�+Dv��d@a`���X�Z��5Zat,^S�<xr�"�1O^lq������ב.S�Zy� �M�6!�II� �`�0�aB��yuuJٱ�ʗn����rq�&�v���E��0ą07�hll����T���u�(|B��B�^B�n�LF�6����L���l
�	��b��Y��uq� D��& �^��x�D�$ ~\� ��'��s��$�zC�S/��0V �={6�EAyYŇx��N������w�t�[��!�O���P���3�l^3ق���$޹��P�j{Y�I�<��G��%�_����G�y�r�k�zFO"Dqn�}��^(�u�D�7�2z��Y@�K�4w*H��@4�s(�X���f���u�7��s�;�x�֪%����
�����K�sud
�-��$2b�H�h�s��9��z�
i�4� �&��6z��ը��S%|��=�vy�A�ծ�M54��V��<1 7����EP.���t	
 �P.QX\��6��u^�p�t��A��eb����RF�Ώ׋a!nsS�&@�k�%�!�9�t�߃�&��m���߃o��$��-�f�q������Ό���e�/O���` yPo�-�� r���䶐� ���I���@u�^�L%쎢��2d}���TȿZ =�,<f�XT. �?��d�ji�g���&ARs��N��Y2x�����?_z���?�����_w(��(���Ws��C�i�2����W2�M���.a|��u��R�ʝv��V5XyWr篕�o��꺺�o�j>������,av�+�<h�z�\@\��끧� ��s�U����w����Ǭ�S?�c^�����Ry���ROw��v��p�Vm�V��QSy�R3E�z-�~kYXzȌ��J�6�3�h�4�Ԛ[H�����8�ϔA0y�bd`
��U�$�ݺR��BE(C~8kQxK��y�c��֩jX<���b�e˖����I�hu{X~��+�d��<����i���><a,[��s�����k���� E��I���202��\�8+ �z�k���Df\s ����Ϊ�=`′G&Z��j�¤�Jm#�/4>��Y��O �a�M�<Dr�!lȵcp��E��ʣ�M�W�|�
��k�����hѢ��暫/<��ow��7���pQ�lȫ�~o�m��|͛%^�5�]��j�YS�ĝ�Y^�����fnkl+�@��w[d���WǏw�֪��
�+�B����u\����S�(�w�%c9���n�a��@���Q�[�y�wܾϺ�����]'b��i}[���V%�t!m�A%v�/�H�Hd֍)w�X�X�k�
]2{��]RR��-��zq�WV��
nP�K.Xux�xŠ����6Dbv��NY�=����U )�ыy�<f&Ac�
�b�y��.C���^t�7���$/M����È(��� $ɷ���vywN.�p���8-��msj��lǤ�\S�h�g��L{�ǬEy� 6=��1�;gБr��(�0a8'_cq]�F��w�8t������Q¬�k���{*?��<�|\�0��\/����ӌ��[�
�YdB��s*H��	2������18�t\yb���9bĸ�ë���V�X��=����o~���T\�F0�-c�G�E�(��\*3��z5O�G���5Ohܤu���$�<-�Z���B�J�\VvU$\����v�G�����(������D���Hh�� ��uE�Q���A�b�;6޹�59���0JN[�ʕ5�?���W����8���~��|�?o[���k�WL�^���pN�ÄR�Z�c@qIJ��.�_(���Fx�����}�݆t������2	�h�j�֬V[5�R�Z��	'�����JCqw*��LCb�s�7B��2�`Ew�T�Yr��
ף;�a�"Z]zX|"g��Ѭ}��d�Y��äR�d��m���g@�ո7�����\� �E0��r�z��`Pj�%�](a^�o���΄�(�I��Zg_Xj�ۢ������眜�8�=�߸ލ���ְI��P�\;�K�R
����1��>��o��CM}�Rt`�����m���H� Ҟ�5�)0���C�cH����>���$ �ȩ��`��+��^HH�M=�>l{�2��>���K��g9)�2E:v����K/��	]��#G��j�s�Y�>l����R��U��ʪ�v%�$��-6�k1nQ�N>��v�� cx$.�]k��l�;'x!��0'�|*UTZ<��G�Y7��{uCp�һ��i1en'��r+�SZ1Os�GQ��6�q��0q��tۀt	i�&u���iXk=5���'uڠh]���ƺ�n����q��.�z�'OX��6��1w޼-�Ĩ	XB��>P��*s�k��HT�˼�Y%X-�61��zF�V�g���K�� aF�9T�����!J+�K��BiC~�w��S+Nׯ1O��r�j%hH�i�RU9B��ܔ��R,4�[g��Tf��I����(��09��51�D���{�a�)~,8��P��.ea�`� ��%�Ch��kJm0
50`t� 3������v�4(k/!sO6 6�N�Ϩ��qa�Є%�$-������(S�%eh�����߀Y����z����vͪ�Emd@J�!���&�^@��j�<ZvBL����꜡&�s������Bt��I�����*���Ѵ��(r]����:u/�znm*�kVUU��3�;kҤ�7m��v��jZ2�-J�}��v�mw߲e�^�s0҈O(���4`�{�ኁ����3Bz��%�%O=��G~�n���?���8���9����d�X k��ͣMH�l	ԋ����!�G!hu�����ǀ�	8"R�8iJ'N���[�ҡ��l�w�Z�GI��\Wg�E:H~��;dY�`6i9�B�>��/�4�b���ʂAT����X�z����-� ��a"��,9b,S���m�OJ[u�F�/%���J�6����	!�֒�^~���R/�)�J
��딷M9����ZnY^v���=Ә�HP.X�B�O��pX��2��m[4�f��tLڠu�(�0!C`v��G�}"?����{��~��?䭙4���HGJ��g҅ �IX�NuL�0�=c�`|%LX�A.޿1���kؽ��MH���Ir(�c{��-�"L�f- 5������r���i�G��|8c(9~�~k%aH�6�����P�A�a���/Ͼ�t���ְ��C�/J����o���j~r�+���RFv%)-�NG�|ؼ9]��(�%iN��Q4j�]wݹ�>zO:� Cd��6�����0O�:S��kH�A�՚S����B�0��>Ԅ�뇗�:u�H�J�,Y|�'>��/������Y~��<��C7,Y�t���PE��э�'qZ�HO&k0\%!�	 }n�폞�V�~���@q-��#di�ȑ�����AsvH1P��.��#p\�h^i,��_z����E�D�*,�mM-BZ�L��^����55�z������ŋS��e���>v�h�4�4	��KRH��W=��j�q����XJ�lB�z�b����Ԕ�jWG�1͓�)�:З�]�@%����b����'G��@1���H/0Q�[���xz(k�A�-y�����c�E٢
��lP��E�w��=4�V���z7rz��jĬQot" 䬾_2dd�=s�`<��P��-Lt1Q��
�P|�<�|���W�v��W��@,��Nzu��"sAT�M�p3�)б6m�'�(�ۺ,
q�(�wS
��Csb����8&g뭗�R�r�R,�E�RM�11h�fTϚ5��7�r�{֧[�U�E�k�sf]2�Hc����|o�ٻ`
�8e(r���Y{줾��%t�sJVA{.��*�T&<큇>v]���	}:���:7��ftd��Ð�II-2g}�qr�>H�Y�9J^���B��_�Sݺ^�q��,Q��U���ɭ�L�@�jX���c@ X�#�ĕ����5�3���=NY���2�[��w��NZ#�,�;=�Cȇ'��B9z��d)ayB�('����1�A��E���~��E�HM{^�{���|pt�]��;�ҕ������� �p8N���׍�E{$#Ԇr�wnw�D��F[��E6 �P�pp~C�'�8���d�D ��0�#��>�s/?-�~�	� X�nlx�6�W��=m�*�x6�ɀ�,��[��!4)ٖ��T�.r�fh�WTL����{�ѝw���J�A����	t�A+n��g:;�7P+�!(4�!�E+d��y@.+#uַ�e�]��z�{qGr�ku˿R��,�#��m�w�,,�`P�N`�I�ҢK�c�E
2D0�ú0:�-�,WѻrE���������͚u�׽��k�u�]��ҳ3{3z�X��z0.)E��4��l�/�����k=������
��B)�7^���6�}�R�
Y�d�����D	0(J�񰱣�.�je"�A�P
V�-����<��0�Q��mD4�aj��x�tA����R�лr,kx"�#�[��eI)�e ���N�tOx��&1L>� � 5�ayiٝk=J�wD�;�1���ԥ#>���~��t��!{ϵ��)y"�W��}\����<�A>t�޷+v'|�ȁ{֞
qC��!�����Ţ�e�p����Y�[0v\){� ����ئ�c�p=��H�`����[����H��L�p�[-X�/Ϟ�%f?)�'��������>��QN�W2�W�-Jߊ�2Z\v��62��dIޒ�K���d�3�I������~��d����H��C��c�=�1{���4�F3��aV���'��|&҈Wi�.��ּ�(/��g|�{ϟ���{��\M���X���p��Q0��U������C:����a{֨�tp\wb|��}+�՚#L���7�.����kϞ�{�uw�u�!Z�'�UP�j�`��"[�:��Z�チ�/;�p^��Z�
�O������VK�J�R�'�%u��ʅ��CF��@3�	���T|�m�Z_@,Ej}*�o�c'GRY�����J)�c�-��3v�e��LVW `P��6m�8ɻ��Tx��f=�)��b�Eeg(@ڑrbCD��)]��	�;���µ0`Q���f�{)�IƁ���J�a!������ ��E��g�_�IET��?p
^6�Q�P�D�1M�j�E�#Eh�}t�v�y�QC(G��N���]�Bh��O^&���nq��nU2��cԍ��$@-�U�,�����>O�x	(;�<H�P=�(䪵�-�������c�}Z���/b��N�}�Rf(_�^X��v�QnP
��ۧ{���0�C��&������W~�+_~��^D��7\	�뮏ϙ��\)���!Nk�� �w�;�x��.qel�̃�n��z��3v�y�w��J�X$yk4�4�������[�uvtFH�>:�VP�a-#"X���hx��P�8��	롗����K��u[o���VHn 1�����	��T���9�98[��]�t�r ;�'�5`]Ͽ��.g��Q�-$��ף�g~!��`�K�<���SZnY�)��y�\8�$���A
�*�%ʛSGN+<xy��oaeWd�����+�X����!���o��Q*x���u�IB�ND�a3
B�`��j�=��Փ�9�1��p�Q��%����2����,x䡄ͭݵ���5���].x����չO�Ct���QNz8?DH�;��5�b�ܞsW�F�X�!���s~G�;��&�)�{~�����,�������uP�u�,��Eܓ�F�8Pg�*M�L	�����о#,4h���Uj!��+�g֫��_�΀�����Y׷�5���͏u���N�k��[�<�G�JdjL��`Y����T����nC]���}��'?^�馛�se�ʭ4OJ-<m-ǜ��s"��-���;�3�Y��%so�$o�/��v��v���U�2U���{nv �浞0+��P����ք�
g �筷�:���O��Νkeb̽��	�T��O��D���.���e_��g��څv_������eVo��|MLx0X_�R3���=��k�S�ںB��#(�A$�\��πBoj�˺����~�u+�N�P_.EYX,�R	�Z�	Bۯ���,�g^o�I��-/�'P�*Do8�1�|ˤȻlQM+��@Qx�x��ۅv�C��}-���7���HC��o��Q�37�T��fSҔѡ�5!_�9��h���I��Խ��Pu����5� ]\>�#	!�n�8���\�� g�*;6Jh��1��y<�����-(Y@z�k�+�@��F�2x��[�0�`���}?���X�,^(v )��2'-⠾@��]���99��zk�v�� �?5���m��@H���MMi� +�q�s5#E��>Y%M��{�u��G/Z��FW�U���O͸����Ѹ�E/l���nE2�%�����?����:�7�� �R���~�ko���gdel�Ai�o�d�e|��
D(6��-s���~���m�Ֆ��)���?�`��[:���c^p������wXc�N��w���沔B�z���!�g����nr_	H�B ��{��Q�:)�=wݥ{�}�����?Dy�q�Y޴���,[W���8e8=)����t6prb ��5��<�}@ *��kI���(�2y鬜N��\�dx����~ŔhYi��{�\!$�;�m��`Ņ:j���q���W]��HtCg�������w�{��P&�a-���)J��I�An��)��z5��Zjm\W e�f�&�7���A�;J�2�oe�M�+��T�.&o(C
�σg����#�w��V�	Դ!���u��w�s�͈������G(�s|��-� ��v�~~;�a0�|���dLq�r9x��u� �b�T���P�n�0�0����8�r"g~��E��Q�!7?`�[ՀJ���#\���v�i�
l�<kC�
p)��H��X�M��T'��tcɷ�Y��I	#!��T[�����УjO����?u��ĺ8��7��r���x��+1л�f
\kk���B��𢋯�Hg��bUJt�<�ví$s��a�鸱�X'�	�]�!��C�v�i�Ԙ1c�mq�@䁩Ȝu����㬑�ŏ{��g?�?׉d9�Tj���-�W>ίw�=�>�ɪiX/4�)��Y �n�2�E� �)���� ��)����
]^��D���AC�E�Q��
u�-y'[��b�
��{�RbS�����G9}�8��ŋ��h9(G�3�\qI�~W	���Y�!5a��d��(D�$y�����\-y"y��?�*�_�(AK���y��� I�,�DGШ/= =�k0w�3^x�Ǜ^������kL���`���K4��$ ��0�X~������B<��^ �r�p������0�H8�{Ӈ�`���[�@�7v�K.x"�؂��6���G����|ٙ��D�'z�+����)�`���c x��T���ܹg'���D&��ߎ��`<b<�}y�ٯ󈚚�Jf�<���KI0:�{J۹���$�C>��+���`��2�)|?��B��t�9A�Kf�ا�u�]_��O;�C	��+���:��l��LR��	���ZK���h0X;�� �`�ƌ-���t���u���p�~ I9��;�3��9?9{���w�c��_���v*M���iW�,����i}m
QY�)C�;<]C��A��"����
]�U���l��QZ�����n�� �S����(n;V��+��"O���F36 9 ���mZ����l�6�w��یi,G:��4a�d���B�ER�Y�kE�Q�V�\qY%}օ_�Ʈ���g=k���{-w�?���H���M���F��'(���2/Aަ硓.G:.��zoO#�����[�ZW5�΅|�5�q��Ƿ�M<Z&�B9�l��y�P�&!p��wY�eg<��4́�
��l z��_�C7\#�¢"�!u���(�`����27��' �?�ު�U�p�`��ş��K�!�H�����I�GD�ܿ)����_��ڿWQ���G���*t�\7�&ׇ,d;AM��O�x�����_��qǝ���W/2R(B�"��#�ږ% .漝B~w�%��B�\z�e���_��>f��&͓l^���*LJ�G��6y����G+ʔ+5S})2�.*ǔ�����-Cx�L�z�]�߽��^{�fZ紇�ƚ�a�J�VuD�0,늯�b���R?����R.�}�ڼ�8D'=
��i;���h�v�m�m�Sݺ.��Gѷ˞{���g�;@�kyqf$�<���6�?��#"�3�Zk�P^��l*�V��� e����W���,�J�Dg���٪�Z�Η�W;�<S;*�����|��:�����3��,G�R��\�Z�64��X�hd�Jف�Dy������c_U[+2�6�䭋��y�=�K�0�ߡF"˗�J�X�Bd'�������t-��~����6&	!w���IiC�&j�UO1x��*X��q���>��8�9�$�Ҥ#�\Qx�s��o` ���(V�s;�,p}�c0��s����9�B��y{�Oy�zǋѷ��9A�{��.�;������RKOS��:,A���v��
Vz�C,e#�u�w뼆K �b�����4!�o�5F������19��(J�ާ�!����}�b^�xi�q�7Cr�M���� �Ƴ���m1bT�_��FGq�=���ܓ��j���"û��� c����X��iU6�֙��/�s�)�&�Y+eZ��d����-yV��r�^���R��2fq�4��5f��~�>������Z��֡V����w�]��\��ؽT�u�(��d)&��k�W�����b]�p����T�Ԑ��Y�͝�}��q� �j�[K��YQ��M�й��>|��/���b�*c<�A ����j���:ZacDYR��9����}G=�ݖ����B½4��o��ƠlVk�B1"m<s#{�<D�B0#J��g��R4P�ukT�&K�_H%��@˶l�2�[���[�H�fB7�l�z`�G��-V#@< ��3��
��H&����D����,�ߍ"��� 0�$�H<�L�FL^fb:�W_����C�WFY"����"���^�������l�|���ǽ{�ޭC���61�~���6!o��ɱp�>��!�� �C@��]��N���pd�_;Q��ݹ�5��^:�%�;��1،��4I~=\2�=}�"D�<���%���9r-k�O�U�X�Rl~����T:G,��'紮V<7Ob)z<�乘�qi|�+
���-^6�J��E�������t�6�l3k�m�4%=��y�Vխ�]_h�c��H�F���WI]��â��x�\y��T�07p�����H�P> Ϫt>r@���S�͕)���T��
�5��!��)@�o'Z�߄�=
5p�Ѽ�c��㜾Os���@֤@��s�82J
��-j�p�Jcq�����a��W羒1�*�t�F��Du^���=cO'�D���t���;�����|��o[M�[m�o��r��>�lي���M&���=U'CI��I)�������'�u�=������g�|ou_����L�zngwv��&M�(OGơM�EIT���P<���b�֙�.]�P\(TJ�,�� �T���]�t�#�<��z�^l�Y�j���#�M�P�Z�,W�U�;���hRg1޾E���fĘ())����Z��֔&Lv�;5V^&���4�"��_+x�dzh� Z���C�^>��>x�a`��0���>J��[��zt?wBG���
ڜ�u�N�#���k)�^�	�}m`6[� �X@|�	B�f|%ނQ�21�z|�������x�b M�*V5��V�mX���6���p����r0�� ����A����Jls�J$��p�E^(��Տ�;�M����/�C��L�&ya�`�f�Tt��.q��s��.К���w�^�R
Ŋt��b��7�������m+��)��2�im�cH�i�3�7��x/
��	����B$%��>�<NǂX8[����	qM8G��H8N�11������Y�.����wR�Z��Ϛ��&�s��|�V��1c��G�CB�p�	�����w]��T�R�I����}:�/^
},(y���a���#=2�-ͦ9��9ty�yz^t~�ۀB��ɑ7��݄J��y|�j�2Ҽv�8D�S��s� J��GN����^W\$p
���������1���,]f![�y�z�slGNb�9�NT�v!O�Z�߀a�g�d�\�Z�H�^�Q����' ˙4�(�a�eM�֗�'��/��<��ka��.̠d����l �}��	����0y�s���`���Y؜hCF���23寝��^
�@?ir��[/�E}/�8 ��tF�##L�EX���u�e��Ct��|t���uv���~� �2�Yމ���#D=��D'��Ҟ�EF��҉�"aFZ����*� �
�G�&S ���3��wYM���E� ��qh"y2V�D�����K�l��O	)ܓ+�]���2�,[��p�0j�������_��BX�V���hM��N#��������?���W��G��G�&ψ��߅%X}����A��("�#�#��RaJ����ǟz�i�4&���5g4?��)�^�R��9��#P[��Q5炁��,"J��T���07�W2�P���IRD�kF�ˁ�'�kk'���� >e-yyt��·�z���l�D:���fٍp:5�ۺ��� �4y�)�"�	Ayr��dO�2���=���!�5[��ɔ/A�KJ��/� ��+��X�O����׵�BX�'�"�И�[`<���s�Nek�|����6���[ZJ�(���Io�%;�LLd��D<��Jˍ��b�.m9֥���@�/�K�d<���1���t�?���j��&f���{�^U�e�"��T4�~#�5�g�`h���B��},X,�*���q/�`F��&4�ae2�<� �I8����z���!W��0v�#7K����N
<L@�١	�O��)��|�s>"!��}�pye��4>�M�"�,u8�|�\�zѵ����"µ�	���	FƁ5�A	�PF�%�'~�l�f<�d2[�_2e�¨ȐF��<��=�Nx2D����X1�k��(N ��,x��[p��H�0�{\�a,<}�z~]��cU���8�ئ,|��c��6=O�0�]��?����o���PZ �2$��t�Bwk8�~][��kh)AAR���%h&oJ�WϺ[o�O��[όv��M���ܻI�}��A�n���wk�-W7�5zޝR&=�qoiYy������t?}R�i�	U�%Yt��΍�O}WY�֧s��uu���늖.]Vk`MM�F^x�f����
���(��&��H
<�Y(Ie�bR	���ˣDx�z�]����5�؀ǲ�OzN�2�ɀ�I�*��m�%�����J��`��OHkqM!�ekU���S{��sa�z���� �C�[����%�F"���a���G�!����/���'?��sj�5VeɯXޜfO�'P�r^ə�^�r�]��K��c�u�`VX�Ec|�č�DD
��k���g�ak8k�E �f���oR\���6kԈ�t��i�S�2���)@���[��,X��0��
��K��Җ(	�Е-�
�J���x��O���<y��"4���ˬ��k�u���t�,ArP��9B�� 9����!Zs�R�.a���p����_}���ZQe��L��>)r:�Q�N�W�<o�Q�R�Q
�Z�B؜5���!���U�v\/7��|"{��ڸZ�M
Κx̌���p` /Mh.ɵ�E_�I�@o/��0�׀E��!�����5�
�,D����И�M�{���U�<�٬��e�A��1/�Re  ���|dB�ڝ���-lA>\[g���.z�w�i:��PBŁ+u$/%�\[�(��㈪
�^�ORM�?hݫg_�����Æ��=���<���!�4�H�f��1��	p��&L�|t�5R,��
�'���" R6]2@e/u�� �ճ�Uj�[ϫא�]]z�}�2
�$�N�W����e����FK�u�5U��Ke4+\,à�� ?�Os�WсnEz���5�Q��[����un6s��� >��c�zf9zT9�Q��Ĳ�F�S�ؘ�pp����g~�k_�,Cx��aZ�*�<���*x-v`(�E�����H�9j����e��<��s�(]1X�����E����F�m����r2�ü�����_���C�Q4�� ��K��[N���������qjW�����{Ь���Y�1!�4:|}�3�t��Ze=�K�yҤ�����f@S��<�G�lU�W:.k��=Zz���&M�� @��[���܌�;!�a-1�㙘��6$?YG����I�����ֺ��1衷��h1��~�uj[��AR���~/Y�Qr<�5"�G)�P�y¸�wAH���9��Ia��˖Z�{�i�ɓ��@�L�[-T��Z���/\"��� ��&��!H���&��Y�BCMN�W�d[[:����6cl@CH���r�����S��]prG�21`^�\K�J9V��d&Lhg�@� H�S}�t()ݣT����c,�;ʕ	��,�!�WM�\y��שkep0p�ǱNJ4�ѥ�*e-�`�˲�:�6��~ ��}��j������X�Pz��%т ��~a`J߂�a�t����a$��/ }s���
>�Z0��&���� @�x���M�to�~3v?"�&D'��½�уrFi�]�$v��0)���^m�0�Mj �!�o"*�aN@�{t�z_X�TX�#E�Su)O�g�aZ��.��!�0�� T�	!��|�_B�aϒ~�:=���UX {ɂ�S�L�?�EA��.�S�M�>e9S=گG�ܣ��_R$��z�m��]c�u�}�k�<_���Bsa��c�x)ڔVk�����X�QM�>ƿ����!�,}��o��Y}��e�:�rd�����̔�MZ�@X�*)�*͗Q*���~�JcXw�dє*W���ǫָ�%�{�~�X?�>[F)ak�j92��7�++G�x����:�%�Օ�t!�#D�18Li��I�:~����
̨#U���NP���7�<3s �
ֺ{���y�%��B��$�	������H�PQ�2=�2]E���HɽT�RJ o L�E'��d^w)TnmQu��4�a���G(r����j�E�]2E�Ϟ=;��.��f̘�R���Uf���a]a=�nlxة̑�?�x�vX'�~�~�w��>O��Ǒs�ކ�1�9t�'�=%ƌ/�40��O�g�[Z˴.��i���0s�I��v��)��?���]ͣҸE��K��<�
�J�s�F�S�Ԗ"�B�Pn�������>�d��2����G��(�a��haQ ��c"��&o�^�x1����'D̓f����S�_�fqg27ALBH^!_�Q�ޜ�-lU1�np�/�;�= �\�{n<, 4�	���!8׺Q�Jy�0J��tj b����j2)�0�0�$X΁�#�	�b��DH;���A;��e,(����gl�(���$�p��#ic��|���k�LFJ.���\�)'�^��:ϲ!�����Fɦ��l��:N��{��C���Fb[k�=9��<B�{;�-�D1s�y������ ���!�q.�x4�f�-�����0b�2�y�f�T�נ@s��]쒫�ʘ�R>I�?0�r��I�C��T����\_�
������H�J�)�����PzƩ�V�aR��Loi���:��ҵh�vPIUeU
HP�Bff�^}��W'�u��(�}�����s�}ӟ)��w@�U���3O�@�,+���RLٺw|�D��5Cxܟ�0�8��U�8��*5P�C&DC}j��!�K2l�0^QS U�<7@�d�3�/���~�ue�I��"��L�IE��vt��hz�x.s�$���:u����~�mW�=���|8G����/oU��K����Ν7wbMͪM���no��S���=E��(�T��z3R4�W��m4JhEE"e�|���'i��)��8QrИ��Һ%�����:���d�9Զ��Z������-���z)��=��V[m���O?S�k.e"+Ƥ;Oec��y��p�up����qmH�ť�ܳ��ښ� ?�[�?9��S
�_�"�0�� 2v�U�=hB�����U*%�#T�"C{f񐐵a��^C����y؁d�sد�W+A#���n��F)R��l}�Ƞ���F�I"�a2��bqEJxه��>�	@�۽]�C8��C���9_gN)�'�{(P����$p�{�f����uq�w�����Q�f��a��(LRo9K�K!0�sN)J��B�
$p5��r� <Ú?x��4t|�Y '#s��F3ˤF�~cZhҕ�)�Ľ5�6)������O`9����{ՠ,���@zx�O�kJ<���{[nL��"M���PzG�jE�� �T9�s�`(,��^%����1֭z~�"�a8��s��--"�sx�%}4@r�}�ί�ļ��!bq�4�yh8��e�x\k�i��1o2�0`�J�3CQ���M�(
n�Z�������nP����Ik$e��5^�(��1���0�Y��fש�>ÐN�M��ϼ�fv�.9׍��㵑9����:�
�>3����s���/`!�g�J�m�I�=4�ƚP�t�ҝ��׫�8�أ������;3�xY����=��39�h-z�'��|����(ͭ�5W���J/���)
��wN��<��9��[��AǓR*��x�+kk�>�w��yJ�C4$(y}^�ut�k����=v�5z��A���Z�9.kIP�� /x F�����K�QӐn�2�G�,W�E�N��a�0��<LB�!��瀜�T���Mƕ�S��d!/�A[5�m5�Ƽ�@s׀wR~L:±f���G�5�jO�9W(�Cx%TR����R]R,*�5!��PH%��W`�~���dUcpt�99�t���V'MDga�ŏQ��h��5���F�����q��B�2��#_�%�Hu�:��!�ijiG�"Z�JT�o4������RD(Y�!��yF��Q��B�0��9���j�lB��I�vߚ���D���[ɺ<��������9{d��c�u�l�.�gL��t8�7�(/E���c�/�˂��d��h@��N��2�
(�&������C�����vf�8�d̀Td���>������eN�O�LUx�����������h�2]��"�d;�~7��B��"�0�����s-�'(t3� u2�?2Faؐ�_d*\C���lƞ�$���8f��(>J�sA��ѓ�!�9/#ՙ��$�};-sW��#R�9��>�`Y��,�|�K�������jD̕(n��$�'���)��p�5C�]��t������Z��o�ض[o� iH^�������/~��+W|��̚Ҧ���Jӕ^xq �g�&�n��6"�����u�E)�����3yJF���'d/�):E�����t_�2e
i��D(�X���CU��	�%�����K�8$r*P�C�����oh��[VUU�Ѻ�)w�k��F&T�(
gc~K���B<�ї��W�ާz����42�@B��B�a4/�K�<��.(Fy��'�\�h]�v������9�-���{7����By^��+<Ϥ� �@
����r<r0Z���gU��,�
 $�H��mͽڀ�u��((�P�g(@<k���]&`��d@#�^�"J��!]�E���(�9u�
�K)5����l��J��\�O��$���P�`G���ձ<o5��a�!8R&^�s�y��=��{���ꓼ~XC^1(qo8�W�����|�`3��Nt�{�i�)T%�5/��r�J�E:� _Mυ�2��D9Za���i�u9V�2�/\y� ��ɵ��
��J«��}?Qp�������c: �p�I��	���ZV�˽�5�}�W��4`0$��w$k?�x������1"Hf6v�X�TJX�-*����QF�v�҄�h@���ɘ�ܙ@!�m�]c�Y�N��[�y�TJn�ȑ#	Z�a���<V�#-���nG��D�9
�9Ⱦ��᭳�b�+���]�p��.��oh������������o�z�5�]��ֲ1����m�*�X��p�7c�CDOT��������mmZ��<
�� ��1̒��>`	�>l[+�i��f*�;��;�P��u�v䡇�n��N���,�Y)�R�f�`ǫ|��P�q	���N/��*jߖj���6���
r�z#'�WT(&2=�\+��3�a��pW��]� D�+J��py��ڍ�Ih�ǥ�X��ۧf�P�	��[��̱�֣p#
��MT�����.^K���Av38�"�ɍ�
/%�	P��9-&�3@l�2G�b80��	���:
��k����B����p�<�>����2��C�=)B��(�s���YlX˄���=��h9>��Y�(%!%aކ�`b�4��QPPb�/���,J����w3�,�^Jz(�sZ�>��ٸU��\�>8v�-��2��\wz���~I��5<x��e�%7�������<g�!�_��w1*��RtNk��X�,b!�%Y���c��N>�j6x�����p�D��6����ʰ�{�����%|����MW�2���<�` �CP����`؁���P��͔J"Ǝ����y�i'2����'D��wL$X��~p��mo����,�2\���pl��D^ؖD�4��t����+4����+<�bԨ����EJ԰���q�G^�A���6�t��'�֫h
��9#<��E;|�;夾�5�\*?�ŋ�~�a�Ϲ妿��������H9�5ZG��ղ6�(<>J|"���-j�ٍ��P/�/�F�1/I�u�;0�	�+���v���!}�͡�!H�%����O���|/������ctn��C�,E �`�~���=��+��� [�N�ׯY�w���W�FWۚ5uZ�D�"@Y�NK3��,g����&���2,����-
��� R�9�w ���Lxא�пtX�Kz I^`�%
O�ZH��� j���{f2ai�[����5j-�l ���@�2��xٚ��eRc���<G�{���4��K	�#�@'F uH_p�\��,�&C�kB����0�����3uV��� Df�{�M�m�5�/r�Ȅu����=���
�A�����yȇ/0��"&��d(�PN������^P�%䨽)[ и�ܐ�kob��Ă1Q؜O�}��B�������#+iԙ2
(�2��������g�]J���˄|�`=��jc,��!����~�t��}���{�9p������%Q�7UM�ɏ��v��ͫN�R!bc�����{i
��,"�\��������`��߫{��\�͓u#Dҟà��K
�}QH����_�y�J�,>|ؓS�N�gʔ��gΜ٢�)��_�s�<��Gno�����h�n�=�j�v���<�c�r���(b��p�������̯"����?|څ��/|˧��E����4�k]Xx1`��`em�Q���/'�O����Ůu�Ԗ[n)L���Rzh�v�5'�<dJ��s�R�����Ǡ$�}X��Ꮊ������8��%�]~�b��6f���ō<��:�pL��x�+WFȐn�b7/ ����7_Y�_��K-g���k�:���:ruB6�P*!�aA�A���k����1��[�|�Rk�q�!a��MXt�<��laƚ���k�2e�E�M�"�/x��pLBY,�x��e�Г��W�S�~��/�kQ=�k�"A�{�M�%t�LNGC���`n��W���P���x������ � �ʂ��>�x�,��$��r��p[`�n*���V� ]� �RO<�Vl4�	>Q�P��5���Kk ,i�
�)9�P�+�(:6lR����깂�N|�JFpL��%�5�#��Xdˢ@F�0z>�{"^����:���?r[
ů; -twsՂ'���x�Z�{%"Ae����7��I��n{ϟl	O�k�ςkK�#O=�{,X������wJݮH�3lٱ��F�}l^�w�3C�c�i�A(�]�ށ������XK����'H{� ��q4(���mP ���<��y�-��a6k�kn�ɀ���DѮŚ�F�����֚��a-[m�e������������{��ҿ\�����E>� �zI(�e�Ü��==h�Cו�{��!��")�#�9��^~ů>��։>��W�{U׶�:�q "xDN97
��.��� �(H���*�g��rШ�1"z:�.�3k��4F�
U����ǤΗ�5m��n�G�a�|�Âo�m��6;��s/���>
�g�y�� �I�]"��D�{z�uQ��|�@F���=���5O=�R�GV+o.嫧�%/0O9�b�h�`
�-g6�eݚ^�az�Bok��헂_H?]1�)�#P$��r���֣�����A�r�Jq��DL��^�kR���PƦ�'/���p +��nY^�q�wx�}�p�2��R�
o�bMr@\v ��!;)�ʥ@��P,`gO��#<Ȕo�����6�ɨ���a�b����d�(_��L,�ʥ��,i ;�X(��wA�buC'Z*�!��gU²F�cT�+��g��s#(��اC ���P���}q'n�
ֻ�%��ayk�#X:��sB���X� 
m0d|�=�Y$�C�������b�y����)*�`$�0rV�5[z�p+�V��3����[��!�߫�M֎1)�#o<`��ݴ�Z!_��V�����yo��~��ނq������f
���zp1W����H��%ݶ"r�%�TvԥB����?���}�j�A0pB�2;z���k�?�teN*!D�(�91n�@̸#�B���,X����r}}"a�j�:Q��^��6�>z�֑�2�g��W�VW�jR��}��1�{�纡����u�zv�m��Ę֠q$�9�� ��:@�qƸf�{���Tq��I�Ɛ�́�����f�����7��ϗ^��O�m�T�)MCe�D��Q$�9��-�pܨ�Zߵ.�V,-u�׉�����y+����+T�LE�YG�'^׮N۶��dc�07
�.*0�䑡����T_'�����l�_z�O�A�s�n`N���iM��4�jyJOҒ6*t=!��YXYֆS���4Xi��9Sye�T���/�wj�[��@xVV�Hծ^%���8-vKE�Q�yB5ٚ��PgE�A�	�
dq�g��㼎;0�1�Pz"�H���NP���Aۓ�q�
��j��5�Tu��:O6�a�X�X�ҕ&�M��Yo�j]jB�O׊�!y>c�����}�F�9u�?OBL� �`)
/{c�z�[ᮺT����J�n�]� n? �Si%?xg]`��q��R��5��u�`�r <q��Opddc��-�a�p�v~�	��uԕ�`y�e!�Z�RU88�� =,׀1��Z�ϩHb�wDDzx����)bd!�4��w�Ls� �;`Ώ5��'GZ;�l��Q�%o�?#"DJ,
a�B(��b�D���H�3��۾�	#�q�k���/�,�Me��5>�$��\�;����898r�г*Zծ�:��@��z&�dD6i�fy~�J����<w	�O�:m����[��;�WU��מ�*K�V[m9{�ܹ�u�c�#"Ox�8���l�^�����x2P�AFKp<�K���x��m�ָ/�w�y���k�t���[n�Y��ǟ��O<~�ց�iT�=B�
�Hy��s�πj/��d��~:ed��P���X����#ϚVσ�.��l`�(D_�`�·��h�M7YZ���5��#��d�\�Á���(�wY��U��!�B5��H�?��ň���򬥔W��~�r�e�jɋ����4���ݬҪ��r}W�"�Z�1�w��E�bY�~M�!�/Z �NV�"�R�Ǐ7�!�B5luBm���n+�UYg6�t� ,��jUi�4:BD<Ԯ������䩱�~2��� �x����H(�Jj������3'-	��V�k��y8������cc��r+�5�mPx�f(a�ĺ%�E	�ѣ6X��B�o<�M��m�
 "���1���^P�p�������jW��yeTY&��~��-<b$�E��`'����30��c*@�9s��xx����eHρ(H��0z�8-��2$=!\�q��B���Cv;�\��Vt�H�Ps\�GG����R0���^�x��8���C��5�FO4V��p�d\q�������.̮\��t�� ����4��4�d9�_�����-(m��}WþH��+t3�P�D-�!�,$��)iY�)
�)�h���z��_�X����2����kѱ��\���V�XSQY�B@�ublW@gEEewհ����Gtq臺f=�ԛ�ػ����o��[nyE����LS$6�U��H���y]{����h���W�ㆌ�o��p Z�GQ�i���h|g���x���Φ�m���=�JkR5嫌U��՚[�Z]�l��|� w|1O�'t�
����XI+G�����g���i���.V����\�&�n�Zk�ʖ���|l{��X2���
Ӿ�YX��;�nu��2 �ε}�5����"���jyՈ�Sի�a���yY�Ĕ��Y��^!���I����S�g����)Q�Ynо*�M�y��
�+G��R�X|�����%d � �]��Ȳ�=�3 R��x-�4���VT�sRj��z[TB=(1�� ������g&�9�_ ��xB���Vؙ�4�&`�:�r��~"(o�&(mB�(]rT��uۃ}���T-_��9��rs��a�z��ƌ%^���aN���<�'Ƅs�+�$%�[	�9Ƃ��v���qOɣ	Ș�� �s�� ˁI.&?6�zU�;���urp���@^0��=xl�2R
���Ҽ\���=�5{[��yc��9B��5|����`DZ��=(�Z}���!=�-����]r�C�SL�?�8Qг<�<�]�q�X�X�x���p�üƖ�|{���8ƻ��}��āV��Φ�:�+vnU���-Tap9����M�Ꜣ��VA��K�v�:OBgc�$#�K4�EŃ�5p��[��Mǳ1`[�����<���� +Mp��|���n��q�s���U�P���x�(i�]�mg�zΫ����	P����-��
�v����{��wo��Q=su���ߤ�^�����'>~|�V�lw�x����b���`3�slc}�B3e�zȆwk�;+����W$�0�=,�{z�w�gn��sϞ�2���ϯ~�������Rw���.��m{h����/���z[�4��R}��Y�=R�c�G{dJ�c�o�������\�K=�W�N�*��̛�#GU��˶:���z�cF�]=r��Ek�ү29��`$!Y�XG����x����<uփC~�n��VU�X��N��m܄�[ ׮�D�r�����R'+����Դ�$�HR�c\�l�`�]ȫ�W�+�w+	ҀX#ϛД��m�/\�05�z�ո�_��XB��ݧ�M�R
S���$�� Q�,�� 1��hޒ�5O��j(A{rEYt�k7�_�+[��k����OFOg���58�<,�M(ʔ�/�}Ю���РG��s~zI�/�R�O˻I�:��w&�C�Ci;�{C�Ɬ��BwL�������ԭ
�劶2��kG<��=��6�z6�RB[�r����sc���Ov�s���B�ܣ�eVf��=���C�< �0�"b�y�����W�iBc�@$0�ß��g��Or	�~��g�}�;~��_�I�a� �J�)!�?���6�h�ǥ�:𠒆:�244|��2d�e�ؐ���lh�π�N+��Н�y���Ο�2:�����
�1�!�Pղ��7���Ř����хJ�@��'#Y�]�R�Y�_3�-0�7��uh�k�߭���݄� �DL���>r�(s���ӣ��
�D˻��{j1��������{���/��J��s���8q£�潺XJ���b�k������;�3k�G���ZxtT�P!��Kt�M�E3_��k�����_��w.��o׉�sL�2��īrt�
�ְ$U�6�R��X՚F?t=9C�k���2g�Ki��N0#���6���� ��5�%,%W�[
����+k����\u�������S��С��]�3�,Ժ6F-�t���GZ��>����<u�i�n��G�ӯR�g�/Y�Q�N� ��g<Y�d=��ʪ�c���Ыd��R,x׎�֪��F����A1�N�Хh
U��c4�oR�8��b/��D�Չ��U,�E�X�1�
���E^[�{�3�jn��D1�>K�r3@tn��*X�S���o�:a��~�(Q uN��I�($f���`�*�*��5�(����e{.�f��y�D���1C=���K�ƽx[x��.Dv	��x�lMD��S%xҒ)!&Yg�nQ���F�{��L�$L��n��ЁS��7M9٪�v)�����G:\Q�% ؝D&�[��
Yxy ����}�ː�s�x<+t<D�/�ʜ�n�͖��=��ɤ����&������'=��6��-oh��C��w�a�%��w�KD�h��2?��&��>�Z��@1i>�g@��i4�a6��mޑʱ��sV�&bQ�s��Т�:��7����3�{�����:�������O�x�x�?��^`�<j˛��E^�7 ["�D+�'6�=��'�y.��a [���torú^(�#�y����-�ܼ�n��u02&J������$!"���i}��	�A�D�јCG&[l�5�+��y�mޒ���N��b�i�{c-ݣ��7V��p	�L�D����e���)d����#�[NƤI���r��H�LV��=̃�pD�Ԭm���.R!�NH^䑫��r��h�aPTV	/EN	�<�r2,�9'
���L�+:AV�:�y��9L�:��iG�k=úY����0�0%f��
�K�<�K����ݫl�}PJ�"��kY<ddC ~���IM|�hv9L㽚-�@�)+&&Q��� <?�'���sP�Z�����x
�fFψ����X��+@�R�:]i��tԹ�? �,���9� �N���X�v8����y�l�-��*��̱�EL2�W�7��.�:�ss�1����7�.���)�V8�~]���Д���ujˡ�q�<��r�Sp�H� �!&�)�MzS���[9x����Hj��al�)�hIxR��5�\�8���.m��+�����Q�z�<y��|�Qk��x(��et�h;��̗y�>����=fL�W^1�LO���`�ȡ;���C/��uC`c��0�(��^x�����_��Ϟ��Wmf���X��B�U��wRj�>�Z��J#����,�*z�o$d��k��G���Ӄ�E�U$Ŕ/A�j����Q�����Ɩ����R�_��a��ZEZ�+��p�֌�5Z��_ZXTQ���]���s�8�yX�� QD��z��(��h�,]�K!Z����k�<��H+O^c~Y�0q����(���9��`��;<kB�]�@��1���%޳ܽc�4C�λ �~�	��J�\�b�n~w6��F��e��ePB�"�����dg����[_vz��3��p~�]�k"���-
��ڇ�0X�ΤM�qdʵ�]��_ȫ����Q�<(�0NL��:	���y�~��]�{~ݿ��Bt��J$e}�5��g�����+	X4P�,l�M����*�+|e����ÖA�1�z����ՠ����cD��ZYQ������;Kܢ���;���?��/*�6Ś�h��,��4�EY���U����9 ��X�e-HYK�������(��������*7\U����<�˺q]�<q��9�\c���I��j5Ԛ3{Nz����贐{X�,��jR����7���Sj­��R�:���׿����.?��O~B7��7y�98Z�����Y���ʺ@���g��f������J��k1&V��]�f߯_]0'_y�q�j�f.֠��A6N�UzT�z`z���-�CQ���\Qqj�X��ݗ��!�<����?��z!I�rQhX��L}�n��%����n���3�G���Q�h�,���`���h4O:DpV h1��"�QC�A>�`��� 79��|ޱ�-(}+���Ȼၳ�}�D� �k$7�}�r�Z�Zْ�ȅ�0��:��cq?���y7אJ�w������d�gm��I����V�'��`Pp�,|\����'�B8n��\ �!�pFz�4����I	��F�5�t�M_��t�F�r�*�М����p?�y�5)����%~%��=�#5�n�������Qk�ω�Z V����lQ��@Kc�PQ�Z����?)I�ޖ�����u�Ys��p�j�z�?����]��[=	��۵��6\L:�P?��d��R賍U��$D��,[�<5q�D0��D�{�q0��̘�:CGN��H(�2!rE�����׫f�`����<ϖ~���B\]_<�/jM�/����2dX�������*M^Ű
�*��-3�������Ӄ�S�D�aCg�Y��!2+3��K4xʤ��2*��_�CP�X��~�@@�򺧋��[y�m�E�_H��C-U�J�2g<s�r5��c�|Q�n�𵃡��C:&(x�LG����o�1��3A9�3�9Z4 �|B8�+�3ԑ7N�6t�(A���~{�JO�ܳ��]�R�cW�#K�Z ��!�	5���	׋�t��Ϝs[V����#"x�I��D�D�N�!0�����`�#k9��8���cxEF�\)�-����D����O�P?��s��x*�*��!�#�F�&u>�o-�/�v�~���z  ���M(��f�u��AI�c��+7���흕����z��'4"G�a�Ux+�U��a;ͩ&E�?����4���+E�A�xt��s��E�Y��w��5�;���?�g�κ�=���h��	M��,&�mƻ���ZOhp'���,�踝6�P�N�:���x遄�����ݽ#����:����K���
Q�tY�*>���|��?��/�œc1Ko�<t+մrb�&�3��3 _B:�;��?G{W�[I�����B�o���>���d䯪��ikoј���3ϝ�z�m�c�%f}I���B;W��\��n�0y��F&`�A���&6� �b�%Q���b���r�\pBG�x�EV��a�<Sz|���'��u ���a�c�	�{#��VN<��0��Ԥ��+�l�T�pz�^��	Z| 9y��\���vO#0!�`x˫;���To�E�'������9?�z�,w��%83 iaRީ�=���t��>w�{�\��OlS�Y"��nmjT��̤q�N��d��Ȓ��PK�����7U��+��[��n�R����n,��$_��V]��#�_��a����G�����y�ʕ�[(�W�zͪT ^���CT�4ʯH%�2�� M�2pp���<҃D
�z&��;��n���ye�։<E��|��'�w�	����]q��o�m��f]��g�ZUۦ�]�'OR��v)���@�f�ir�FN�Pj�sN��NL��/��zi��UY?���'��Zw|�a�H�8��mv���}�����u�)����'�n�$ƏU�p���!�& �� ���v��:���蛟�ɦ��N`�۪S��D[���Ҳ<c�� ��+a-�M/����8�E:#��XV���h���E��ވŕU�{t6ɠ��E�6�.sT&[���&�,�Ә$a�pN�Qf�P_/����@���M::�>��h`C�&��.g��P������^L� ȫ�T��Ĝ�ՎӃ���p�5b����2��l� �.����D�'�}'��2���:)��M���?~��l����ګ����7�����r-��r��ӣ�;���5�����p%��n��}��_���k�;H��O��N�4�4�:
]�T�uց��{�w!����/
�K�!��r��F�3��+���f�����;O���?�����eĈ/�8�Zo
5����rY�=ƻ@i��	Jk�p�zt����Y,}�
�'�&���RwO?�wm��ɱu<�X��1�����n��m�|Ёo��]�Q�zR%ú��~�V�Hdh��ʫl-�!�i�u�����#��Gx8Yp
����˔�K���B���a���j��GчT z�^����j�@ݮq˚����	_[�4
�����ה�`��`��@��YΙze�q��ː���irb�[�K�B�Ä{º%�����f<��JN��:f��@�	G���������;^>���2JA��^E�<@��$t�F�d?���J� 7�R�ϊX�����S��%(.ߓ��#������=��x���8�ȅ����{Z�6|���zy�(uω��XW�ZF��O?]���/8���|�K/;���~7}>�s�3Ǽx��ͻ��C.�~իf���_���]u��;��7�|�B_)�NѸ1V�NU���y����Ƭ1D �U��C��� �:� ����טt,��[�"��bĈw��,#��J��:�W�$�p�=l�'�g���2�?΄����
��x1�uO?� |C#�5�����@{�oxߙ�M�ٽR�ֿJN�/Cy�Q����!��w4�{(�� V���4&`ba����\���@�P�l��y��+?ɇs}�t��L�����sL�=+%
}�/ �������wFr�	�\�Z����S~�{�S��	G�=B}L��g�p�{ͼJ�,ҝ�q�q h	��-D���ʶQ�	 ��DTS/��$.�Mp1��v�� [Q�I��{f��'<CV7y-�W����o���������D6�_����(�wU��G�9��{�w��.p��QkJ�B�KWdN*����|U����?�������/��ҥK�%�TP� ̙�Y��j�rNW��\ɢ��N��w�{Vƥ�]~�>��ו�m��Vkn���m^�������=5~��K/(�M���}7��!���65c���(�}�._i���!�)�����`8�#�}��zYo�/|`�Ĺ1ୢ�P��b��/����������> �tP74�O"����0Q�T��a�U�2�� 
�;/G�m7�yW�{|�N���BJ�Q��O��FY������>�?�Ma+�a�ùnJQ!�?���h�ak��t`�9�0�}x�N�� S�Ж{ҵ�[�x����By��b#���D��Q��8^�<��g>X��)��x����q�"!p�P!�ܳ)��)���ӱj�����|A!�'O�8g��i����;�^�).,���=R���1�p&S)1���R�񓡉������|P���%��=�
�tQ������Ĺ�맞zr�����U���V
=)u�}��W�U[�r�k��vo��o��W���~�4{��O���&�⃫����h���p�00�E��s~�3R����8찺����u��Ck[�sPx�Gy˖f���p| ��9�g�$8!��D1CU	9k�=�A� %�� �忞��2�Pˮ�l��/������g~��k1���GˣFj�(*}_H9O{���S�;��qm k�V��@?���������RL�	�1���=�E�PJ��<mY-$�e�L6��(|FFUe�y��*c)4*�NBS�EBK����9�a!��k��m�[p+�R���u�D$K��E�I%oWJ\~>���K�B��n�4V�(7S� ϝ ���d�\8�J~=�q-^��J���W�לso^�D�
g���=?����[l�ţ�o���c?zT�]��`'R������p�[Q�>��O<:{��[d����\n�T���C�83��ԩk��}�ݧ��?�{���̾�k/����_z����ټ�r�Z��F�J�B'D�*ʭC|�Z&�[�礸���;�x�d6�l�ۖ-[����(�j̠�q8Vȓs>�~(Q���`��h& ��'C]_�Kfp&�2yw� |G���9�b
���q�w�����k����!C�uD��n<��H)���0J�!��lp �S�����fn~NGk���7o�SW�zy����O�X��ô�_���B�6�r��T�tK��d�n�>��2ՌB�P���6����Kx*G(r��
�WSOM>G��^�P��;9��2�0���pL������9�h���g1JX�������K�s��隄J\x���k�/��r}/Y�hVǤg�rL�a�	RRV��ֈ�|����D�
�axհ���S�O7�7G~��n�醫��,B��_Kh��(��G�a����V�nJ9�Z�5
��2b�4c�[�ny�%�|�W����c>�і[o���~����G)�%x�!2��@dТ�T�X�"���`��f�:��ӿcm]ӷ�vۭVe��F��#Oo-�a|���I����m�;k 
�N�<�wr���F�#$l�u����v�DS��5���9��үW)�)�^�&�G���M�T"��&L�S�]�4�K�%A�Cpww��-�38w���[p��K��]����{��Z?�ګw�^ݻjF��&z^l�>>r��[�7q���&-�_�����?\{���B3���:�q*�
���l���R9�l�G�4X;��lf���'�'rET��&bhe�4&7�	t���SC�N�M�\	��T����v`6�����ӆE����x�p_���ŏ�\ #J���8������,z��lF.���׮
x��ϰ��܃u�̒�<k5�E�e^���+x%S���R7D�2���2��X:�I
��6�sm�m��ǻ1�����y���z����6{�1iLz����c=�ه�@N������˗��3���/���A��Rr����}������W:�E
Y#\oT6��[1��T�a�{�7O1���f����\��ڿ~�'��eC�H�1�NX� X`pH��
���Z(��D����q9�
���B�b!K�3��'�%�x~��8�^�(^����������ٷ�}uS�|���D�h��O$����$�N?���Ջ�E�9�Jg�R3�À�RU[�Z���ƍ���g�Iߺ^#� � �&���&�+�$d���y%"k>�(��S�W���^=.S�_��P����F�(TՏ�*�����;hw��&5�	���))Z�sAt; ���i)�0y�Ӹ���� ���r�#>��9�`���q� ���=?���6@�WKE;�7�-�4��ؼ��	7䁽to�G��g��QL�n^<�S&Y�,kv3Z�l�]�o��}7isFVbGJ���c�Î'�",x�-�y����1�l JT��r^^Cj� O����T'�����f�i�.��h�*�!���z{bG����� �v�%ثTl.m����~�����T7���?u����jC^�C��tc�;�St���'<�0Lߙ�۶�O^H�Y�+<4�]LM���̓3��������*2z���&�&x>�0% �����%qM�?��u49ylD���E���t/ޕ�_�*]���0fJ܈'�6�μ ��mT�CF�*����n����K�ܞQ'ײܿ������jn���(��grTOa!	1)�!����p&�2�#FcU��`J;U6�P�'�,��e�a�j��S�vN^㤝|�=�5��P<٪����-��C������q�6HN���U��~�����ț_k�fڸ1r���v�?;�W�/���CK�������QI?��6A�}����R��q˛䵗��z�`kuh�,�s��v�߭n�z}�z�c�2��eF^!��PD�cw���a�iZ���X�ke������pλXOV.2I�x��m�������װ#>"�����S�N%-�\�������av���j�Q�������s	�%
����d�5UI^��-3�Rv�������q@���s���c�/D�xL!��I�-�4��` ���Se��l|���3��\�J0�\4M���������	�yZ�ᑺ3�`7k�x��c=jǲPx����I�� ČA��D���M<l�ڂ���|����#*کt>3�f�H3&��;I�SF�gb7urW"ƴ�O0�S^y=)�wt�1���V�u��ظ�Q�5;膚�=�u��x��e�\_d��8��`'÷EƉAP��k�i.c_�[K�ͥ1K�v6���7�
�����'O��cƯ�
j�eM�$��-v��UkU�;�ɛS��R^�ҍ|��o_ܰêϕ_
�hS}�����mٗ�IE����e�R:�Ú�|IXkKm9���P�����%�air��x�3��H�1<�q���;�5�w��y}�����&���{�\[�9�RV�G�'����D�.W�Z�~��L�+�((0��^�l���w�2�c�]������%�ik�c�����8�4/gX�2�L�N����o6%0���=�rF��c;d�x��uJ�i���9B���Dw,��9Qo�_Ю*S�9�+����B�mS���mer�cy�C��2�ϥc�4��%9*8�ʁ� ��⠞v.�r6^����}�?��"�7�JJz�m�[)�}�0hs_F=ȾN.Vx�IGS>�w��}><�	�ޭBTwkLR�1&�Lro�Wن�q
7��+�w��N�o@����-W�9y�[�7B�7rɴE�`]���Z�iy�큝��̐3�T�J�5�d�ʏģ�Cry��"�|8�/��[{���$E�$��bv�)ϿJmI,���%&�5q�����
�ɑD��jn�����0g�?�@>�( 1v���וr^o���0���3&^3����u��-�q���BsT�\��Y�v��a7�Ӎ�Q �ʕ�^�A�3f����@:�
��g��=�!\�lpF���|���t�,p&���)�Ξ�Cf�"K�ı�/1k�"���p�Ԝ�����>����,������3M�n�Oxދ��#e��pc��Ϩ��O��"����KuI���Ж���ͷ�����ԡy5 � 7�6iR@8�x�%b�s��43;>��=����I�f��������'E�%�D��Jd��va����{&�y�<�x��E��~����|bɎ�0�ʺz	�n�&��I�� �^�7�eX�f�IbO'�w
���i���8.����'3s"�������o�W��ߟA] R%I��j&�E��a׉�1QbGeYE����@��]�����i����R�{�W!��KunQT����S4��2ޝ��ؙ��U0���8W �p�����܀����1�}��¾M7^���Q��A�Q�A\�#57�m�+?���5Mm|e�O?�Xtkk%:.����2�j�rJwi�\3�NߪYp�ׇ���.]$�u����I�}1%��7�+����ɬ[������c�`?/���E���=�R?��w05I�\����b���}��]Ԁ�ti�gv�ߴ�k��/ki+*�ސ?�<�4���9
uU�����"`�L��v�\)�V��/T=��f����+�T\��@���^n�+&�:��/�N � ;����G��!����57k!����כ�O�E�R��dȵ�ПΘ֓E��~{!�1�ŊG4��Jk.��6�3m]l#�&�W�6S�xm�fii��%��t�ϕ4�1Sxb�t��giC�@��И�p��:��l�*���
QEz������X]~���o�R�c��d:�/JF�ES �9��(y2$|W�PTI�R�B�O�o3�C�.����yW��w��#|�C���-���,A��OЎ�a���8��|�w�
�+� ҈h���֪��t���c�=����E����&�Sm�X���%�i���ڎ��p��Q|K~����O�����W�eQ8t˗�Q1�[�kw�*�Gx.���F��ڻF���fg_�/|{���5�b9y��_2�.m��7)��[%��r�m�;������P��*���X��>��=5m}C������]��ǋO���`=��৳�����S�d:Ŏ�jO-���wb*�%�wISs�(	�L*�kw�v z�_��8�C���� wnx�1���� ��F}�w_Q�;V��6��񆰱T"������)�$j�E']d{	��Pd�"�Q4-� �==�9@�g����v��������A}!���j�j�=���b�d��u�g�r�C�Z�6 ���;�y�������ͩ�Q4=7^��e�Ο���L��s���AƽB��̻�b
�1#�l9�$A�5�)�inn4�E�ݭ�KIm��c���_�����&K�	���O�)��U��-���f2���~�œy��ԝQ�C��EBγ$I.��d�f�먯q���8��"/�����#�����߲�����Q�� p��B�gjʆ���+�U������n�����SL�8���o���p{𘂛��Y��W*B�Op���g�i�6�d@�-JK��W�$���{԰_�z4 U�q7R:���/�j�ܧ�\`Gi�R�߭��t5��8�Lf����1�%sKv|08┙��c)+��������w5�!"sZӉ(�;�٤BQ�9��S8�h��ߧǹ���!��W�I[����@ȳ�m��/2��/��
����0�yӻx�1�g`���S��z;�"`z�s��<���E|4+�`$�7�тp��?�n�RUpt���;�	9!E��D�Mqx\�h�	5�0Ǫ���x�fO"j������S�Q!�u����Ps�4s�?�"�����R$�;��L�KU��'DGSܾ����q�Lo��W��n��8���5[W���	_��x�P��*�xf�7��"���~��u�4Fɵ{�|ޡ����]?N:3��#S��@�d�ǅ/z�s׼6�)��+��y����<�u}�êw�8+��ӏ������$���8��&����L<���y���g��"���x|i�Vi�z֬�й��d��Qd��-RR>�7ҷO�at�An��\���?ŉ$
�ߛ��T�|��=����#�IP}��V�Z^�
{(
����F��`�/��)Y�{����"�
�G���Zf.i#�2���F�����"B����inVn���m<b�K>r���ݑ2�!�!i��
�����?�6��H�$��ycz��t�&L�+n�?X��p?�%+1�8倱����:��ː�IG�(�a=��)n��ן���B*��0����B�2�KCYCmF�4>�'��n�j�u���Ų�I�Ĕ�(�\
P�b�W�t]��#�5�={��|�"��O+ �Xɻŏ�u)��Ǿ�|v�0)t$ј��Ū�V�FAG�`:{;z�.�H��{T|�R'��.�p0�RxR�d6�W�u8����<Dҭ�̥{gR�پ�r��]~�K��q���Mc~|Y�E��$��_����_�jZ��v��Qt%��ß^�X�/Ԫ��� ���|�A��pe��?��U�A*S�`�	�)_����sD�W��nl�S_��3Z�R�����<R�'q�[�C�u7:c�HA+�����75��� ��Vo�ظ��p=���<]��n�L���֝ ߏ��vS�w��XX��밓Z�/Gf���� B¼�31�Nƫim���B�X��vM|�aUp~�pJn@���C����V�^��i�WUw���R&z��"_D�aN @����tC�+4�5�h��:�+���/��M�z4�l3_�!�[��J�t�1`���+��MѦ��!eA���&�^3���]���8�]]�R�¯�\������ԳƳ��,�i�D]C~�7���Z-[��1�a��඄�~#P�$�!}pv�BB�<���(����P�	x�� �Bw��	d/u
�D<r\�
߿�X1˱��sK�2"(˭8��k���zv�c=G�eRiG�f�*A�u7מZ�+��η��㓤M�Q霜�2�����G�ݑ��F���9����,k��2��*��,��v��ȑ�����\�wυ9p��M�ؐ��U�玮Ȅ��_��%S�����P99*4�P!�7=�4�9��'��/��� ����J=t�X.4�֎�P�ۑ�xZp���E��s��|�{t9ڂ]�}�Ku��J�SXl�+�z����\Ћ���c�}4�[	O�9P�ţ���z���,ZQ��,Ba;t˳���!�;Iz=� t�������&�i�ʉ�*y��>v�ѵG�w�W�U���ǣ'&��t�R��}BI�t��\�_'�F���'5��'G� 	�;�͵�m|8rĳ"�\�>�9����Ս�W��;��Nѵ^k�N%��ӯ��M��y���M4�G���M>k�.�q�a�uI�ᐝ��B%g[O���B�ɒ+l�li�锎i�UN4py[ݍ�ae��z���(�������������.�A9#G�p�C���4��c�x`.�
���hY�^/��NM���"!��:�D�J��	_��~�0M��6#1t8�J1� ���5���Ư��/�%D��Zǫe4{�0�~j��t�s��6ꂞQ+H�Ry$/(�L�ۦ6=z�s�U}03D� �֋�_ޗ[q��ypC>'�S�G�'�(Zr�oВ.I|��=���߸pU/ϯ��3�~��qޟ)O��O�[=>�Ο�4�	d['C�&�֮��X�(�*����Jq
���
�JλN��kҮ�R#���D����ȳK|:y��L:���n���&[$z9-C���?`YT�qK_�u+�����x��	j�\��î=_��WP���}�Y�ew[���bz>%~�/��S섧 ,/l�]X^�~��G,��Ԓ�y{�?ڐ��un�F�`�|������g�J���^>V��
�{�8���l�\;V��(�c��hԧ���`g)�)����p44hU4vp��ݻ�D�m׎Q+���H˞�}<�3��?�_�Lt>��ʣ��Զ��d��V�!�^�.WC5�@y�̭���g�����$af�ۮ'����A�7�L_�^pf#^&Eɗ�!+��{g���������K��U:�k��s�}�}]ޖXX05�����\��	����٬c�= �kmu]��ː<Q �5׻�@c����Zu%�灵��^� ߛM~��qE�B�����EK����r{{[V��cu{8����}�٩c��pd�9nR7,��<� ��V��/�(�C��x1l��1����o�{�߅7Yk�,^�z��S X�ͧ��ۧ�#�8Jd�y݀�ǲ����"�j�A^���Ur�bU��ekO�W�禇�,pNR#ӂ3�/x�A�|��[��|CA6�'OL���p�B��g��nQAO+w���E�4�|���jRN"/�� ˱4�ĭ�3���^�H2��g"��g+���9����ˀ�� �Ù���e����gl*�fWy��0�N��m`Gؿŉ�G�ߟ�/��q}Y8-&UL/�'A`b�rf�L!5�1
]p�jr_Vט�v����g��;q'~�v�hTǞ�VF�4ְɺv�f�(�3Z������m�����0��9��{��e��'m8?��G�qZma��b�Wx||�  �"�튖ȿ�o����x
��<���{�z�)�<-����d��@&&���X��
f
�$��M�F��PIE�Ƀ'��λ�3�wFF��_B��K��x�!��0�Y��������Ap1:�oݥ���=���Syϱ+n2u��C׵*!���%�1U�p�tz��T�����j��fVX�X���h�׷ĄuX��Ǔ�
Uq:s��f�]�=��2�>�9�^������ E)��^��H�c���o��K�%�:P/�VK
]��$���=S��-N)�h���?{_+ѓYb&�#��!` @��k�;)����C�9�=�(���AΧ��^���f�Ux�<��*���D#�j��S�I,Σq	~732�5Ώ�ܫ7�\yz���%H"7\���m?��`J��Q)�m$�����^S�S:H���E�4O�p�����]�+k�.���u���G��<԰d��8lDA�C��pؑ	��@��|Yz��~�R`)���wR�V;\��6w���/̸5�]�<S�)K�C����ն�_��8s4�ø,���_S��E>5�=\����Q�)2�l��O�����'�������g�c*�)hCf/�v�t~��]�}rK!���YI�P�l��_Z���4(�]y�c�0c����Y$�W�&׀m��_��܏S/|��$]��� �~���:W����j���,S�A=�y�K�X�H|��J��#EO�D�"@"OA3;��)�8E �}t�����2�;\Z���2?�!l~�s�f�=���`��#��ReY2l����l������)0������e:�~�M�<|@�_�M�d��C���y��_�DR����[l�e66fp6�0�~���m�������{�b�!�]?S�����v�A�r�í��B��)���Ǉ�V�C~�2�Y���&��`j��f����Kg�������1��(8J����	頻2y�l
[{���oYpa�x�����`�#id�&��v=6�1qP'L.�������.�� �G��yD>�q]�}��6!�Zz�&�X���w�&�*�2|����������µ��vz}���(�%xB��K�@O�d�a[+έ�O����n�|��1�Y���M��_��15���;��������a*���g��X7t�lPs[ ҄�A�\']�HMFl�nҚP8�v\Ia�ʩz�.N ��J*�W(����
]������0���c��Fφ�!��C7����3e���q�A��S(�j�Qs���~� �}
#�xF�s"����J�o�����(F�fa����}��o]2L	�~= 62�����%����	ɕ�w"�FO�=�|	�$�4!����V�ȏbo�x�������{U�*�ɐ{ ��E�������V�=~v���iG�V��C�m�����jv���ud��+��E�#�Eh��_j�v��aj(���4���JF�]śG����O�;+�v9�4nyk�c�M2�폫�, F�Df�z�+s����/�xtɐ��&$����,�E>���όc�
��Uۥ�؃���s�I�|3C�������Ɉ��}N��P�5��DNMN�ɶly�D�p�N�K�� Ȋ��[�{W��ҡ�{�ӽC��D+S�>KU07D�)��Ve�A~/Gb�lSt��1���ӏ���󢷇��6R���҄W�j��i�����O�_�f<���K�)� d_�3�H����|zyw��x�6Q�<W���$Q���0�9����9�#���DĨ~y?+�e;"J��蔵FI1�G��m���̕������T�q�dV�z���s��ij־��l�^i���H�ЊV����`�^���/qL�e0:d��5E�d�?(c�����"�)�"�i	�aq��T��� rx��Wxc1�)��ܿ��߾��?-JD�z�p�y�̣���Q9�p)�I��Uh��J����(�w�X��^�/���L'�t��?\f��k��ʏ]���Lޓm==K$�].Xt
�`u�������̓U��4�	�����ֻ��<D�j�����!��'.c�`Z�(x7x�m�����m�����4�>��.۹7�s�g��V����m��5�휓�)d��)�����v��l+��1���'��2�n�W�#��~ذ���$^Ņ}�ƙ��4��C�*�$o!|��gt+wz+79��6x�d>ڍ[�'L0��h�~�Ǉ�b��p���Rc�Z7�{h���}�V�L����_�����w�W��ǯJ�2TNP�kՉUW�]^�ڟ�M���ţ�.��YM	�>�'5�zo�pճ�&�Ç���Q�^���)���N�ۓ�����[���+�X8ۑ˟#[k�Z?!��B���\k1��CG�^l���LHݛ�2�/Rr�gX����ڻK�_�k��YD'�OȻi.rs8����	d�7��K�"Y�@\�����ҙ[f9w<ұ�#��ģJҘ��*��h���\;�V��cb�TϩD���H�P��BI[�2J���\����O��q�6Q�A�_�p����Ka>��_��Ȉ��n3?a,�0hڻ��Y����uop��D�)��&Yb��u�-�eg�h�ԶWm��Zl#����dڝ��y׳!V�R�֡���_Dr���YBM�Z�ـ�IQ
S�BF)����4{/Z�>��X�)�R���i�˙W�"@[� $�D�>�?W����"x��̼(b�U��aA�����)�5:���ȁ��}"�����m?wG����Rqһ�<���J80-��S����%j��wH"���~M)�����J�-<4M���f/�hĠ>��f�
�yǿ��w^�C)�ڂƬ�N����s4D&��5��qé���?)	7����L��{���Z#��Q�{�R�I�����]�)eÜƱ����t*��σԧ�=g	:\�OvK.k/�Œ����q	R�SkR�q���u��q���d��C����ԃv�jG$h|A�t�X?N�"~�`�q�V
&<�2���B���*�$�'�q�z�� �ق�������9\x(B<�����+K��<Q�eL	y���8����o��2��?���?p�o�Q
:����b������'�x?~�S5_���G�n�uC	�=�^�O����M3+a�^ OO7���Q-}���������q��<�oÎѺ_4���Q���)�5��CT���(?�^Q@����K��+G��!�6 ���E���=��T��]b�n6�5	r7�}��ë�S�5yn2]�IB�¡LP
�^a�ھz�0f�p�|��eyQd�6c���[w'&��i	��i`�;f�3��%�^����uJ��s��9��̧���葖�h9J�,�Q�#�A���t-/'�8���@P��'��r������|**�v��I���9W���}6E�1`+��9o0UY����)P,���"Z�]�Sh�����D֟��������O	m�B�3�+�݌_�'�/s&dW�'��eұ��+���Y|f����<���^�����l��
cv���Ta�k����լ&uf��ǉ�����D�$@g���W�x��_���+�rI:ci;�Y�$�tX��ϔ��'<f��Å����t݇��Ja�y�C�֩��ƹx��:s*����ר���h}�HX�����5e�wl�O"�����L#�%[��c㨜���MB�t���*��2�x��u�����)'�C�K�+��_^F4�v6�y­G���#^�%	\xU-:���Y��]�3I"X^�Q�(6��1���8��+�Q�]1s�@:�g\�<��0��r_v>��4��6�_��,���^�����t+��={��OvC׾��G����
�_9f5����b�|���o��,vj��(>A�G�����?�<�_�M;Ȓ;����_�{;/����?�SXlw���S5ʹ�/<��q���s��j@�����b�	�����E�AD�oYJ�^AL���R���x(���k����d1����S�lF��Hײ��6$_�`�>&�pb�AJK����S��+5��ſvz���Kq��6X�b���5�p֏+a�"�9f�zWDS��Q�X�HX.>�=�C���1���r'�����]Wf�����O�U���5�.t�c�8���C��C��['��毗��0�"Хr���B?���H3�BwU\J #��,��#�b�1N�ŭ���}0��fEG��:�ZcR�E�͡����A��$[�^��B�5�M����v�%a|���&v�=��]`��}~Oɱ��d+Z��t��q߅�����=�;7
2���ϝ&G���-j|�g>�V�,��1si�n[�&[���ۯ@��4���	�PapMmN.�	��%��U��1��#�n�QĺA�����[���"Ƭ35�B�h���Y�_�;Xb^\V��Nm�MՆU�����=Z�(ދ��,u��:>r
��I� ��6�Bm��������lKC�w1��@86��6�6xR!�l6w��"��j��g+s���" '�O7�~gk�a�j�3J��bOȍQQS�-�}����	��U�Z�`����j�	L��Ï��'۸\�4�f%[�>��	�sN�U��yq&`E=i��BN���ѥ= �%��h��o�p�Q�t=��D�� ���ˎ#�چ�Z('�/d�p�0�'�:���_�ǟ�=�(R+xq�`ˬsGNA) ���!�1$����v�pf�T],ꕵ�|~V��j���h]a��c[�\�%i :2+�%}+��N��;X�����^����0	H�����������jQ$@ǘ[�aQ�HL�X�vrߜoeD��<v�����J!dC �����aNdr� ��z�f�����ܾUfQ4;c�0����C>΃�]4(u����FR��<Ru�&���'L#����<����;+5��'hHE��t���~��˂?^�S��_�&�	�A��&�}�̇*g�~p&O:��g������dߥ�e����N�1��H���ݹ���v <�$�Nq߃\-���N�>,^���w�tp�Vʮ�G���(q!^K�t��U�>�����Ӥ�a���.&8>��[�x(���/p�#��FkA��L�R�P�.�я�,����?,�L����B�
���h�z�5x`���P%J���^W�� A�14G��RK��cS�3zT?܏�t7�B�}70�Z&�J�h��t;Q ���'OJg�!Cݻ+&Ff��p�_��wg��X�����e�Q��Q {`�Ai 1Z||�&L��՟k�R�6�k�V��ԝ��y~���m��I�9�\��g�w��$)Gx�M�O�o�\���O>҇/������
��iK�3A�{S(z�iu�\[{FJm^`�r���z.�<�^��@�2�|d���%���8w�;&b�ydr���Q���%0U����Zug3*���<(' ��žAeߒ�'��:���C�^��Q ���>M��oR����g9���5P�}����/�Y�te�"��9�c����6&���Dg*����N�i*�4=1"�^���؅��Lkl��ௌgml�쵁�2H�ȟ�����Z9����9�{�\Z���r���t�"��ΖYA�S� �m:���B��R�:�h�J@;FrR)���`ekP>i�uK�ϱ�t�^�N�!4�;|�3;';ca��y�Onx��j�?V���aNx��qr�@G'��CJ8.;5A��V�,N\��HyfSo
��H�|�f[8F��'E1@���X��|�O�|8~s~�2��d��J�B����R@��=&ܠ�W��Re�CkZ�0��?�	����>Z�P;�'"��V�`=�g �Y��߄�\ �P��E����ڜ������o����ȂlQ+"ߣf(��$����}#ɉr��<0�>�����e|���I�ΰWD��c0��=���������pߪHu��l�J�mKƊ�uk�C4|qnmhB#�'ժ�!>3Q"����Qa_\�#���}�$�G�<��*��j��p���ɗ�<�8u⽙�x��x/�s�I��PR����9d�Ⅾ�QHxޟQ�F�$]5�-E��+;5�U��cM���4��c���C/���seu�����$[I���2�����Y�_��z<��R�c�i�-�s(HkPG�FdB�I{�����ʘZۋ��ۇ�^^^a��p׈~g����KPF�X���f�`�Z����B$���}k�'�_>���G��n-���
x��Jq-0����y��k~�B��~\C�u��Ҵ[;]���d�l�F˹�xlն�R'��Ш�:�5��.c��@A0� "{,%���0FtWq��WW.�<�,���L���ӹ����r����}�}�0K���փH`X��~`�HJpݴi�>t#��Z���}$' T�|���]�����n�w�<I�(�da�����f܈��s��䙼޹A ��9^NYօ�s/x�Ϲan����N3"�B��G���2!9�����OX���[_�:Q��F�N:\����"�t?_�4�B�y��;x���b��l�Jya�<�<:1cJ�V�0,~�Q�i���VU�[P������N���Q�E���N�j|����|ÆM����u�!�%@�
8[���Og;�����D54�d}�qr�|WN$0�����S���?a%d�K�UZ���r� ծ���E#cw-߇*)d/S�$%���7�ƹ���A��>�c���d��K4��2���L�3bD
��]~�5��S�4[�[��M��I����篏Z�n��Ժ�H_�F�3	"���^x]Nr4/����yt�7�ǮSw����Z����7���Fc�Ǻ/] D;���=BJ"R�ᬣ9w����8�2F�фW���z�/΁����ڑP88��t7��m��vTƘ�s&k	|��an���m^�WtE�L2*�L�@�h��8~C�b�C��
S�/12��R��I�� R��j���=J.����-�Tu
���5����-9q=���8�'=l��ɒxaM�3ݭ.�����M/��*�|�9U�A4֦7�S��*K)n�)y��z����(�#�0~NF/��	b�jim}�q 
�{,��^�k��'IXD�ܒ'ldCJ?f	��� -Q=u���*��x�_�r���Ү�i|'bI+�U�K�mTT��0m��.��E�Z�����1�`h,�$X�ؓn©yj���{E�93%�F���'�[qPzv��.���fîN�r����R�tC�����V�����M�������]95}c�Mr�\�|]�s}�_��s��_^��z�0�D?u����t+��`�r�Ύ4g�@ �T�iq ��l�M�w4.��tb�Pa����&Ɩ��d�(�[~�⤟�L~��]������nn�D����D nO���`Il"�R�|�Yr�n�V�M���ZZ��F���S����3�]x����!�}�M�dlT�	H�J��0���ĸ-ꑽ)��M��^,��?�&�p0󽼤� 9tWs.0��f�ٿ-��p��\/?-Sa��M���x�{��Tj�����Aa�kCs�n��Q�J�AK5�����隷�w1^��L�YD�9���Z)mf<Yìs׶�.���V����nP���y������Zx��#QÞ�
�`i�ua�Y%&g}���T�`bOr����Κ��S���}7��f�/&ū��ĸ��	q���A$��VW�L�r=�g+nY�:��q�۞:<�ož����R>���d��L,,��ve)?]|m�	~G[�u�b��J�溠��&_t<��u���Sp�Q�q���U���]唩�`�����}����y�yPRl�;l}2�a����0I�A�T�3�!�cH��,�;C�lo�mG��ZY,2�&u��߹�F@o���h�J�X�%�x�ֿ�S��5T�9�6�S��٤D2�߮Qp���0E�<6n~��\eODWyÓ*�,��{v���"q6�K�Jf�ս��u����q�� �
��� �~y*`��*��V�R@a��U����H[����^}�<#�vNm�H��`��9)�B�i�t�l��i~'�� �Yi@pB&�<o�B}�aG��hUmw�o~۸�d��<�!"�r&���<�}u�r<c�[�:ϛ��W������>�G����c��>�ow8K��� ��$ֿ�$���h<�9��Ɓ扗K���iK�4Ź(�tlM�Q���w7��S7�۝�{!Bxc�d�7J��fyl�!1״J����1��ӽa�;b��P��׌���uC���=<��\�\�H�3DÔ���]k��^���KKK
 ��9߼�h'YI�+"T�9�)j�1��(���,RV�p�s�mZ+?�Ȭ�9@��?pu� ?QE��AEM�=�����YC�	���W ߺ~ǟ�����#+�V7AC�8��p�*��	��u�o�4�K��槛������d�=��@���p���Y�r�;؆�7&�i�cIt1��rd��!��@V;yI5Ë�~h�cE�6x�Cp4�����cG�\\�2���É�]HL���2
��]6*�A檐X2v́��S���dmr��e�n%�����13O��x8o��$
��8љt�Me���oh����!O~��F�f�1WHΈ�$@�)H��}8d2��3c~���A,ƢoN	#?�����ؾR����nnB���Țˍ��N�D��j�z챑�w��Cn%� �ͧ�
�#�a�Y���;Y��s{�p����3kg�`?<���&� Tw=k��|�ubed�h5g:�����������~�p���}�N�wp��﨧��_�n8>���Q�>U�φ�?�����9P�����u�uk��ai-���b��L|��p����Y�#��NGD�W9���/i=H�An��¥���h�j�S65�;'皘I�6�w�NZ�e�CҸ�^U)��h޳����-	l����X9����B3��Kl�X��H=�nWxƝ����PayA�R�jP`���ǔV���A�v�/H�2 '��֎A��̠Q�t�]ix���4o�^E�7�:���������1<Ak�Z�7T�	Z黶�#;G.�����
HrP=��(�ɩ��nL��:��}��}uq��㔠��FJK��Z>�d��[����V�k�=�Mv�1�ɜl��m�l۶m{�d�\ӄ9��^��z���^X��� ��;�����ɹ�0�H���췿�i�1sa~��8�������;�^�]��=��Âݜ�3��= �Ƌ���_xxc�`�N�Y4��,;�'���#׽����֧�zU�+�� �,p�9Ϸ��\5*�� �1ZD!������!���&<hb����l�ڬ���gi����t#�&^y[I�c��&Q�R+�2ۈ�lJ�0&��[&��Aq���[���`l�Z�g�y����$�g��Gi���Ƨ*F���!��ԫ�Ur\c�lHs20b�|o����\o�u���tl��C��f�����-��-�N�b���Z��SD#�P�Ŧ��M �lԢ��w*[y�*��	F�*����Hg2o6�yb��&_��WfgJJ��ށ^6t�����]:w�zkr��(�~0��IA���|E�������Kb=7z�6-�����zs&W���.��f�#%�M�H��HB(7x����FF�$�U�R���:.�zS����~�o�����ݸ����Kޟ�&���g#řhh傍I�~�B5]dfd@%��323X�W�/T���g�%��E�#!|P؇Ɏm�eDK�q
'�L|��&���;���'�ܮ�^i�=���Á@�q���r��)#s�̮9@��yd� a� (6������q誉�����"k����F��\q�8?���� �8pN�[uv��?�����KY��瘹��ƛ����MXϕ��"_6+X�\#�9|3K����c_�t��dZ�7%f^�	�!����2����k~	�������U��;��#���mN�Ī�=����<+l�s �[�'Zb�V聢��Fra�A���6�LxM�ác���<1������������[�s�MчQ���пpy�qڳ���QO���vyRoYT1/ �*���e���r�P�rXj|��Ph-�c�X��ݹ�ݘ�ԫH�L���z�����..�H<DDD�����*s��DϹA�� }T�jׁ�R��*��pP��x���Ec�;t��R�8\�>�x:��aŔ5��j��!��ی<]� ��9)��R��7�"-J���G���I! �gd�ET�b��6�-&W����K��F �ā�����l'
��44�O��4���>@U�|�#��C_�#8�F:lsvT�@$;�����ټ�kg�H�d�X��^��j�>�ڂ{N��m|ˌ2��v���I��k��Ѱ:-x.#�]p����,4{��=�k�n��,�0nz�_�;�͙d~�a��~�h(�����=,�M�v]5������C�xqX��\:ə�B�`�BL��\�t�����07���U�&l�����K�yJ�RΕcnO؛���+�a�Pѻ�-��������g�7oD6/1� Xd2��ߩJW�_�8�d}���=�5AW�%�XF�a�V�y��-�0�Ԝ�*=��d���l�:lq8�t�4��%RZ�x�M'L9'�<�]�X�r}FEp`Sv�r�A����A)OǍXp�S�|�����\K�Q`E�aQ~��!�����j>m��j�38��A"��Ld-���5�f+�@Z�&�S�rzK>�Ħ�a�7�L�H�e�foS��ˣ�h�Hf7D�TJ	d�u��P-B�$����:>�y��'�Oo��@���#(?շ:��;5Dt177wT�읭�=����1��z��(0�����ڡ��3�{�αc���H}�(�/��`�2B�ulU�2��(��y�6�I�ck�� ����X�Y��~�\���lǞ����@Y���ۆ��@x�6y�T�ۻ��l�� �ɥ��$��Ċ ��1鴌��"kt�,����%��Z%F���Ĭ���	�8*S�p��S�/$#��E{�w������0�]ƗΦ�5{��e��Ѓ�)�0�_ �gY�C���Wt��Ѻ��=_dK`��溨h�H`"�;e ���2J�D���hf*�:��\6@d�d��q��(vɗdnQ�K����F�����"Tt9�^��TN/#�#��]�\�J�C��-J�w#�:��H�0U�>����4���+ ɓuUs�%�Jt��AC9= ��
��Pz��o!��_)��P������;0�g���P��|�a�n"�]wx�����N��r;�~��&��1S�d7���B��:��;����q&YNƷ�w��-��RP�ø���Q�th'Q�h{�jh]��}��~"��4o�!?�E�AZ�Y�t#M�2+ɕ_���,�c�����g,��+Ԁ��rp=�}�Sf�0�1��vi�#d�z�y�"���t#ە�Z�h���^e4]LԴPH�jќu�J�s�R4�:'��`���eE� ���#t�&Nt*�8R�M��L=�ʎ�'�������iΏ2`#�R�� �@�g�#^<]���Bng����1sR.�E��ҍ!!5����e旙�S�Jl5٥�L:��v��&���a����Ɂ�Nk�Dr@�ؤ ~���u�s+�[%`J⥠Rր�\�d1dI��7��i{��[�JgT��B���[�×h���+���QY����y��9ʅ���av�����?�H/0�b ��I}v+�=/��Γ�����[���)e����,V�rLf�耲tA����}�Zvu=�K�WH�E~��3cB�=Ff��]0��,E���3':�)\����'HX�Ycè���k�M��<7�b����u� �s��Ǯ�s�KƸ�����H0A� ���$~�����M5ݤ��s�5FFL?��">57���� ��6�E"D4��l�l��aN�>N�Vl~��Nk*��b�Wn��
J��zX�d�u��=�-��u�GY������4kd-�C
wQV�lD����� �|-z8&[5��鲩2XE�����{�Gk�{��9��o�5�k����������c��M����G
�|�\O�^%p���M�����Z{�x���|�l�uD��<<,�:J���s�j�"���m���fz�-�u�;�R�����#hK�F�k�%�gi���Nح9|Һi����(��UD3�g��CH+B݃�ja�++(�%B2�� !�8fu
އC��_�BLLL`�Wk�/$wyyzQ�(���R��}��N�_�^Ua����ߎ	n���kC�`�y�,E*�P�9AGcO;�� �YЌ���(^�W�ǥU�����^,1�葏�;B)0#����Ih&*=,l�Q\�l#Byzy��(��{�p��ȉoln���Hޥ0O���i���ɦ��'�Vn�ˏ+�2���q|�xb��k�w�J�c�;��T�2[�O@�!fѨ�`I�mF+�g���@R�^P��v��!�����6l������m����X*�z���AL�-h_*x�p���4����I7�{�"J�$3�R8��s־�;�쭀%�I�^r��*'�h�*7
��/cJ-6cDKm������R�) 0p ��V9��+��ZE16W��X��JK�!�|�z��
��A��8hb� ��ekx���V�<����2��t�P/��öyg�1��u��o�*J'�=���Ԃb�
��WTv���D�k�2�Sc8�f�s�����N%�!$��2�*�Uր�ɡ���|�I�#*�d��)��O
�lg�W/E#7 cB�����1�eX�����o\�*k�o�p�h'��'�R��YU�=5��z�{"�p�skɘmh�ߗ�D��trr�����z�--�-��Y�Qs�
#�����3��w�쪝��H��e��9��>��H��#B��`�$�oY7�J����komo
�$ڠ�u��P��a���1�y�l�F{���=���������,�ћNL/�%^RS4��U1��ᛪ_��T8��ݘӈ�r��Ї��oѾ�!��kK	W�L�u�S��)���4�x�Y�EX�ė-�ʨ$�~�qN�f�O����GH��&���V@�#JϯR�d;��'�&�C�>���`�\�����` �f�0���@24����OXu�*��E���gj�n���r���&c��VQ����G)5�h덂T�M��*ɓ�S�5�]m
�'2n����w�_	\���4I����Y�i�O��^F���ҲW�������i�ɲ�z�戬����XN���,��:������b%�F���y�G��k�Iu�J�ӨX�Q����l���A��FK$�-����zH�G˯A2R7��;/a��Z�Y�������G�!��mڻ�qv�9r2'���gc���0����7a|�"��nd!�Ƭ[�wڝ�k�wPq��E Sj�v
�oJXm00�U.��.�wΞ�xR�-���Yx��H��ѯ�\��5�`������H�1�o�R$�nM�\��NT6DR[Z�F0^>�:��1�������,���^z��"�:��8�z�j1�x5ioa�E�o�|�Wª��^|ڳ3����˝��=��*�/�*4�a�����W盅���b*Ɨ2���~ ����4�Q�3�4��iD�h睏���?6��5��-D ���EQTi��h�'~v<��2�� ��V/NVP�0,c�����24�����(N�`��pm
�eM�[��\~�2N���$)�Y��5��2[9�7��'�H�4�a)s�~��#�44dX���m����se����1�x�Z�����.��Gu���|,��c���X�p]�͹7�$�K�+"��\�����.zVP1fĀI{{*I�f�EE<�~;��n�鿾���ON���ֆ_`ZS� 4��~S*�ޫ�+��z{�ފ�c�]�T(v�#w���B��`�O�2�2:]p�#V��7�qF�o�[Bmm��� "���f���ݯg�5D��B�{Ź�3񒟠ʾ�jg݋�J4Μ���t
�=M+�^.�LGH#[��!)�ʫ��^]��m-�����T̆ao��]A�{g!�_Kl�(�6��́�E^�79�A�x�^ߜ�,�
��k�'@��h="�O������Da�w	�~����{��,~������"�E�'�H��Ͼ�,��)�wC�B?��d2�%��X�҈���I.�5*��NO��_�qm���7�x�C�P_gB�2��^2Ϛ�Ǿ�b�UO03<e�h����Ŷ+l�c�c�翃_(��[�������8듢��� �߻#��?}�q��C����M�(������V4:w��M��1�w�)��o��C���g�2���$����'���,��v�;����x�35W���7��_�����n5��YZG���[�?�_������v�
�/k�c���h�W>-�ey�/��zJ���.�.^M޽�����o1���#h��.Փ��/�4�--�ZQ3in
̠���Jv{� 4*�Uri�O��,~�c�&��SD��{�*O�:/�,3�c�_6�����-�e#������0�w��K�-��W_AqY�;esާ��Y��	\�sˌ{��0>���H��S�'���~�&i� �滔ʂb��Y�4�i����]�ǘ��'�0I��P����#w;Zh�k���q��Z�{�!Ӻ�=6<X%��)���r�\%�C�/$}�b���&�~�����8̂������OR:���aG������9��k=w\[N݀�Ѡ�y��O�!�츑�`aB�+�;"sh�I��!�ey8%������Ɏf�5+u#��%��;bc�;�^ ,�.9�����D�x��l�ZзpS=p�v�2ivU^��e�:L����`��Q[�|;�1�Y�^Q/�L,���ѯL/�ȹ/���4+��Fy4���aY&�����$��Z��}���_�A���3<����\��D�R{�V]�I�Һ�M�H�"o�{�����d�m�f��o]�U땯u����hJJu�'�������)d�����]ǔRG(��{����WokŠ+��vFa �Y�u����/Ep*9�V���P�9�7���z;���}TZO�_�E�c��+?�D�c/1cu
�#���&u]�͊f}��I���U����1�.Uw%��K[������*���ZM�jzb�B�̜w��/E\�0k�é妉^G�h ^�s�h�����s'�]Ȧk~>�O��tLLɞ wV���o�)�v_1RW�}(�Z�?V?�h�-T?R
d��ǘ���M��m]�q���bR>&S�����^
e�e�!W��'�W,����WІ-ʈ�ؿ�1G��S��h0+ti�!��{_���df��("\2]q]X�K�C�S�c�_�����oʈw ��욂B
r�1~���
9.�:�%EX�L� �/�hR��ڢ�{K!3��ϩ��r��D�7`����*���v%}BTb�!�ـB�oy튎"Ύk^�9	1(��� K#�� U1}�M�E=����fѬ֡n���^��,�1�+7�Z��Ж�a-K����b/��j����ң^�����W1('��GK��ޖ�r��23[���'����M�|J���G�Mq4����] MQ/Ӎ'�����o�w���s`�G$:��TXq ̓�}U�� %wj�y3֌���o!��ynͦ�9 Ȧ<�x�m5F�S�kiAE���[�|/����J7���/��\v���G�}5�y��K(Bў܎�K��F��Q}�Φ����'w3��_t�k�e4]�트�L>�w� �F�n�Sr�2(�e��;�yD�:d\�$�-9�B�%]�V�\<A��WM����"�xx��Q^���vnf��9|��!�/]�gή���>�WvC��e�F��D<�9h�k�<�!�ys���(�j��]]�Y�fz �&�����o!�׏�t�9��/�$�F}�,��A��!5��k���J�z�M����0�/����p"D���Z+����t�@b����`�\�:���7˘]܌�v�V�I��cҽʬ��{���ܵ��7`����7@���"K�П�X�C���$�WE!5�.ʎx&~G��Ig˘���
�1i��n�(��\2��Q9wo��[P�FA����n5o��Q}��3�R�E���& �*�o��$�'1#P���A���I�!��퉔m�y�?�
˖�#��ЈH�hN����>.���7�����V�rx�%j������n$nNK@H���C���XE�]VU��2q_
y�,�;e�SA+�X��=�NZ���)��Vyh�W[�,���������]H�x��8q4
�!n��ta�Eq����C#��_eۆ ӷ����"����+!@�v�r��;����J���:/#	���g��VG΋a�V�q>�-l�\�d���<�hC̸X�D�>Qt=���	�e<@��ӢoP��NY�O�l�$Aa����Q��� hE�){H�0b�1�u��̐�5)4��MGq�n�uJ׎�)m���4��̕|�Xϫ�'0DB-��k�+@�b�,Ei�Ԋ��~]]�w��	��m�+)��ɣ�^#J�M�v��O���Lr0��/?K��45FόY��>�X��~>*)����F1` 0�g,����Ao�`�ޭ�xݨ��G��h)KN��H�n�Զv���Q݀��'�~�%�QO���_�!�ݰ*G���.�s�*���u�7��c/�	�)22�c5>�e�wP���M�ZB�����U��SĎ..?�DEP6�4j:~���:���s;������迗h����L��P��cF�&��*�]�o�V���/�ՀC��F��ǌ:fy���MaϮbBޟFE
2站���c��v��l�1��f�rx��v����[�H.6����i����0��h0����e�,��R����\^�ef��)�Et���(�81o۷��%<�-H�<;ӏ��
3��e��o�L����
'�njį6=���\����'��Q�A-^8bI��5�jܝ�#����+(��T^�n�-'=���
׿�|1�aAsċ��n~�Y���g�&���An�e�Nb`��	���w����Y�_��x��_Z^�}��tt��.x���rK��C��hB�$*J3��h����N����lC¸%��Ii	SeOꧢv�ta��[�#u��*;�u�/vOG@un:�y���>WID�I��x�������S�9H�+<��p_��P��n˴�|$�j�����p�#��V�I*U�X���̟;H���ݬ=�!W��Û�3V�9�Ei�����*�`�=�z����C-lE�5T����rvJ��_�-v�?��9��d�1�Ľ=�,
�r��cFL<��}A���Z�7W�H����U����n{�Vѝe���'���&%��}v���Gʐn��ּ�e�Ю�+]�s��,Z 	���������E����y��H��丣{�2j֑}�oQ?���b�����j����I��;�ӫ;ʡ��_���T�lj�&�:5���l
s��M{����@�?5⫏G���P�#e}3M��B��vʑ��wD����A\���͌M�K��k���3rm"����֙�Tq^4&�z[���� �Z��X�>�zz�S���I��|C���Ff�	;��T�14�=���)�۱k�	2�����*ʋIX} ���}j�%n�:-3������tk�
}�j�V�Ɓ�K🄨:z7V���J[�.j�Ɇ�k߂6˧>�\9k���XVnf�!rpr¨W��U�p�p�o��L#�1�5'�1qOɾ(��tcx
��(%e�#���(�>U'%0y����0�z������jH��]�N] )sS��I�yk٣N�|~�	-EP)���'���P�h�n�VSY4[=-������$;аs�4*��σ�Oy%%�J���c7vԃt��C:��D�o����?ӟLa�'B� ����z�Ė�jf�ܔ�.ә[��C漾ݭ�_�m��������㇆�'��zX�a��
9V.pO�fN��F��v[El��c�6�椟�O�$��AX�>�	�fm&9�M���C�e^�ۄ��~���J�s��{���cz�ˌӔˎ�i��Rz�J���$�+*�����o�c4|S�1sai���Z_N���̸U�[��)�m��jj�����b��>
Ǖ�"�!rn^��\fc��7�ݵf����w|�GE�F��/ԏ9��Wyf�8��χU�%��������<�$��vnr�g���n�o��=���o.b���Lf�̰�����
��3��jS�ƹu!¥r3aE�� ���f0��CI&�gt 7�_�\᩟�p�+E��.�����w��⟾[8�Ë�ֵ�}��ոsʾ���)�ߏQ��������?���v�׾�Fy�
��7h�j��W�>�~%���/�ڿ����g�/z�.\��3�����
���Ph&&'���qS�U+˚��m3�O��,�W�E-���Y`�Zt/(]F�dn���ml��cyX-��V�5�*^�	^��N(������>��y&��铟��LLK�8���ב��O��i��[O�W9c��se?b�S�L�.��C�����:?�
t�7����\(�,�����>��u�U��0TV�`��w\��M�X��W}
qH
���u�!^Y% Q�8��#ucs��Q1�Zj}��Ϳ9�OsW^l)�FϹ���0|\ŰCy��l}޳N-�&c�	u�h�j�H�n7O���Uđ��|�ㆄ��.דyJ��~ �({�ͨ�2�0-N�ERe���:[�x!�"{��;hƝ$�/�8wsz��|*鉨i��E��ҫu�,��%� �s�Մ��e�>_x��-(h��l����#��W��^��-=�2���~�
�z�q �=�ǑT���F�b�QQA����U	��Jm%������+���)�{�7I��q�tǫ�s�E�сɣ>����A��#%�.T�\�mȐ�|��s^"olHJ{�!�Rɵ�!nj�w�rLԈɭ�lI�N�{Q��?xe#n����@WT��+�E@�Q,��oF,�( ��of�&��Q�)uT�����ksM�C�Hob��nzV�e�8}�r!�Z�YtV�bNL�����j���YȬ:߉�rg��;IKs`u���x&�����^�0o�8�_0�o��m���gpZ�SK\���c_͍��%�*��-f�Ԯ�|��}�P%b�\7����M�h��H�����u�:f�c�A	�q����e��������	��|�x��Tl:=�t&:�� ��`�7��~�[���ӱ�uy�P��pⱯ�>�����64)%f$�K��%ʅ�^+7��y�ؾ�_�g�?��y� L�'��{�d����ctQ���3�hCL� ����IJ��f�x/o�)�t���K�Ĭ4�w����y���vuw��3� �K��ou1�{��W3��D&�A�g|��b{J����e*��d��ܜGQ���@\���֨�ghyMM.���
̜wI�u�V��e��VK��f8�����~k��ն�Mwp2���y�fQ҃!L
����
��M&�3�xo�0JC��l���}}b:X ��9��kͰ�C�XI�!�*g�>6�9��,q�-�Ml	r�����Gk'������-O�����m�ċ���w���.:�:2Y�k�r})5���|���g�x�rN���T�����y���S4����$P�c��]p�.M\���93�4�M4μ��M����J�<|�u�23^CV�<P{l�d���{me"ۼ��=�^����+��>�ۧ-,���^i/���UO�N�=3�x	�ac�����jT` ob*��g�	�F��[�����y#�z��D�tL�HZ�����t�X���d �a�U>�i���m0МP� �OK�)�7m�M��nm���P���Hj�(ฺ�����q"!���7EݺF;|��쐢��k�����t��@�T�̦]�Ne*ڕ�&���P$֋�����ͅsNo��_&�3i��K��̟4n�&�~�����[Nߑ�H;�j^���*]����N/<���[\�%G|�Eg/��q&R�(�}�5��*����no���0�=��:�\�A��}���mC����迿�Ж�(c��X�~�)�vV�����6��*]�[����QH�r%�Y.h{}���M�@?<��M{���mMd{j�X41%�iϗ�m�¬��=7|����W��UD ߩAb�z*����W������B�/��n��:���� ����L��J�s�eВ.~z��n�L� 5*�@Pp��0�邙B�V����zk9�YP{�[y9�Լ��k�cX��:|Z�ѨZ�pZ�(�hT��U�	?�I����'�۫�qyzKC�kS�.\T���+��>��)�s��+3���U'���W�߷_�dJ��)E��&ڗ��M�`9��Q�����8�_��X���F�kA�a���#ő��I�DN�h��9�'N;)�l-0�%�.��3K��/�UJ��5��q�.�.ƪ��#(�α�9�©��E�Mn*�H������p2�:�����c2'�j�@y]6kP���l곍�z+*��d�.����a͵ӫ�E��bjޭw�.�D�\W�餟����wlɴH�D��� r`rs�EX�gx�Η$��By���Y]�8v���/4� �Z��¥At9wn�c��{��N0,��[�o넽+�/?�!��RŸ�魳bA^/nv`��8��v)�ӹ{%�_a谄�sa
�Bm��\/\����H�&���iErs��!��*7�aK&�ܡ�͍����A'���ƍ�P}2��{"Ja����g6�J�$��y���R��D���0���
�5�`����E܉��>N8�;����7WD_�~���	����!@PR�Gc���B�Vxbߟ@�T_�h�T�vV��0�@e+z���Ŀ�c3��ll��z��oR<]q����=.�8�� ��|YT�5iA�X��ͣ�w-��;�b��s]�^L����'fϪ՘[Ύ���'!*7��:�/p�'�=��N�x����6:�%�Q�Z1G��4������Z+#3^zW����SݺQ�s� ��e�)�Y��Ȣ��%l�gfE7hENn�.W��K5���3��ʪ+[0�Nw�[I�"�63o���}�o��S׫Y�y��U�ti,������)o���Q�Ҟ?g���K��w��F���	���.1�����u������iO��nơº.3n7���@TGY9�,�������S��h�EtN:�I��=�ʀ�s��cG�
csPr�_NN�q�`�=׆ֿ&�U�&A<��z�D�)k��PRQ��p\�N���w,@�i?�Ԩ�w~����7V��DU�D�;�F�C�/��h�2�ΘS�`��|��#a�&��ǝ��v��9
�Sk����R^�)�����s�M��IÕq����fT��t����nٽ�DW��Z��G�Gqp2Nx��O9eV�P�k����1���Sy���'��AY�#SA�7@:ʐp�4t:�7T���~��v@�3�3P�_��J���$+�q�<��
�-�2�ņ��z�&_�0y�)�:[�"�,��9C�I}ב�F⮨�;{�	� H�dd_�f+9.�V�����&#J*�y�v4C%S�=rʊ��(�����ƻ����Hzډ�%nљgC�6<���O�j�[F��(���e �%�+#�*����G����Tc��-��6���Jp*T����b8�D�<P?���k}IrUC������C���%}u��Ì|��\���z݆i^q�@C�&�i�+�/~����J����`�RYl�>a_
�GƳ>�K�Ŋ��?bfC����o�x=p=�c�$���e��Yu{�aYMF�C�A��g���D�PRS�@Jg��D<.����X��]�Q���2�(�,�(3��x3��W�K�0�(0�vb��A�T{����#���r����-%�Լ���2��!:��+[�x��*7'�f�����]ֽ�y*G������I��P���J�[�0�V,�Xe,�ܿ��p4.(Ơ������K��5m����@�9��������ڄX$����	���b�� ��D�r[��Y[�iv6̙�gUU	}��tt�OG3;&
"d�X�?D>��Q�\�)�>T�pa����������V��X�Id1������}�sN�<J��u�+㣞oG��sF�#(.��t�vYc�{<7�]�q���K6��� -|F�nOW�r��`�¦V���~��{�n����c~xp?��Y��ǯ����NYS/ՔD���&UX����'�|s�/7QFD2�/�TW���
i7N9dʨl�J������
ڥݵ{�w��Υ~��XG��̷�L��Q�a&���-ߗK�.��`!�:��	H�_���q���b�LD�������Jo3΍Fl�0��47��:2�L5���jpŷ�����i,(ȹӤ���L���6�8 ȉUZ��4���"��&)��"�.�/w�/�H�$�
	x�qg���D%M%�H���,٤^�C�>ҵ�8)��Z�>��]� #<i���#�{�G�_���W�u��,��ѡK��o�1(e�ǣk,:�����;2>��a��]��i?Mg��b]��8��o�����'a��#�px��YF�diRӧ��?̰�w̽���Hf@&�01k5��s���MH&3@�i�5�I
y�]���C�6.b|@.|
�S�C�d�=�F�����GSZ��6�G2k���U�� �
���!�zϭU��RLnˡ�a����1�KA�6�����{�����
�|||���:�{х��ԧ���~n�W��8�ea�K�R��v�v6fH�E�E��堄a٨� q>L�����A����ѩzR5ۍ�ӭ0R�� 8{��������gZ��
n8�h+��h�-3��,>�m�Î6"1�� ��߳t����u��\U:BY"}P`H���y��̩��JS���^���Ke<���(�a�KW�Pln��1d��q����1�z-�l(C�,"��l�K�M���Qy@�wx,N��?�M�o7��+�u��E�u���z�d��u����֡ݿM�zE�-�z�ٵx�8�r䏳�9���~$"Y�\��Y�h>]º9�����b�<1�9*M�j��"����d��Y�j���~�T�X��|��u�7�]�<�����n��:{b��������4�ΰK0��S�t��I�Q�����ꦲ��-��ুj� ����p1Թ?�Ig�#�d1¦�Tݲ����"n�g#쎑��=>9��4�rs����?��p��(Ȅ�zɣ��O��ORN7g���2K�U׿'W&��P�#���ӑr՝��+�� |�˨(.?��("��:�B��U̫@H׿���� 3��զ�B���M�7�{�Q���9^���L�U���!W��u��&�hg��}�]랅��ڹ�����t��>l��Q�]�g1�ٮ�w2�����$8�vca
tH�S'bv%^}]����~�G�0�"w�*�îj|�����K`�)���_�`U�Z���5!(��;�ǈ�z;��V!}܁K��q��yY�G�e&j������U��� >��h����M.�ĵu!ZDFױ����j�1�d���^q��t������0_��/J��[���xB@�49�3�Į~1St_~���'!F�\C;^�b̫�
��!.xޫ����Y|V�����1ǐ��{[�"�!��"ȚG4c��,&����'O��E�;�Z�u�U8�ҟ��[{Cj� eix���t:�� �W݅ ��j���{�QT2n���������P�u(�>��0�9mh��ާF�:�$��9M�Hy�B�k�m\�AQ�{���.,,/=��pbk�0M�{?r���쥽:��S����>��D1�:j#�⃵����a1�R�ZߒT@;|c���?r�\���ZQbe%�Wi�����9����\�����`�t�#��h$ ��C�^M�~�4MK1���|Q�?���:Hqt��Mk��?�೙��#�'ӊH.M���[#Q�[i42���l����<"�B���^"�35
_Ԣ'	{>�z+% D���h$9`���!A��E4VgY������?硔l��BK��+���N RW�EHx�X�D�E&b��dɘP
�T�(/YGe�O|_�{�q�.�"�T�ͧ��?1����~2B.@�M����.-$��/V8�{N��v�sS3���S]]� ����Ъ�b�Y#vn�g[5Bv硗>����l ��.�I����1����2䭤� �.-g��c�iQ�~a��ODn���S��5�⽖,̺�\X��sa�����;7������PF�7y�2�1�V����X�I��~>m�������?��K<�ٶW���A]m�J�5Q�z�u�CTdG��b��.��_"�m�gJW�ɵ\~4��o����@;)p2�3��:rO�l)��T^�(=���O�*�)�Ix>�e��h`��:Tu���eP��K�u�PK�V��A�o,!5�O=��o;JF"��;��}j��L�-��M�:���zε<�	r�-�Vn��~�3%�&�����a鱅+A������ci��������<3ј`J�����,�-w_X<��R�}�.�.�χ�����O�PC�b����x����3�'�g��*�(/��)���7*&�[�C_�!xs��+OD�Լ�� \'H�E$c|��fL�;*�����Y���N��tC3ҒMu��V�\"�4[�����c?�U���L��/�H,�{~���ǣe�Hև~h%J1�iz��R
q�	b'���qG׋�{:�nn&�����DpAd?K^��&�:<.(Ƶ����e!7�O���fb�K�m���7F�q�����1y� �l��l�����I@�*��>�y����+U��%r5����T��˘�p��?���h;\�BE�,���3�j�k�@m��_�*~ASF--�>�m����#a���B)$u�8�K�V��}�6��� 'XsJ����j**���Ū�R�� @���d��j�������	u)�����M�!��8���V���`������!����y��V�Ra��$=��}{�@,M^i�%�a��p�U�>�n�AHi�K�� W��o��AyҞ`=�癩��v@C�' ��&~u~�:�޼Ö�qN��@'��_�xL	_i�N��`c�y�r��6l�s�j
L�RAxh��/������	=�QvQq���yt5h1���pFrD?u���MB���Α>�9��9L�B�9�g�a`6cdd����@m� �+� ׼.�"���θn"���V[YeA����2@Ϳ�!�2M��q?�$:|���pa������m�JKK�j'�F�;�'��K
�"<�@#j0{�Z����ʊ��ډ-�--��MME�i�q��#&U�r��i]]�a��������x���$$�E�C(%��ꅋ��*�h�D�ÖK?���pQ��������+��{�O8VRT/).�=��#1յ�0�D��@V���V�����r"���1N˙���b���|ik��|-���r�ͷ����/<����DO��uQ�����8��Og�93�I��0�e!��e�wuu�Z_;/cv�Ztg�˘�����5�'9���-N����HҊ��a�=l4�<`���� ��b�I|��K��"��O�;�fX��� ��/�����"#�m �`�K��ׁ���/�����ӵ@��ZA�8�����G�$`�Qd�����X7��,J�C���&G�lN�41���[H�p6�T�l�QFa���Dz���*�����6nܠ3:�1`����W����X��f��]@��8;�t��%%t��R2�{��Eʐz���,�G1S���w�T����ܬ������SW�G,kyqQ�
�]n��g?��f_D��0����$�սte�2��-[mc���\��*��wiKٖ#XS��w�?g`�7�ҫ���o�u�՚n9n��g	��o|6��i�dZP��)xÅ�g�f�;U�����9�扖�^���I�\W���^�o���s�~�-��'5P"��&��%�l>�9���XN�ǳ���E�'�ee�H�;�����_�݉�k�?��sG<��?ƌ�@\�2��Hr�i�-��R�0P��ٜ�}Jjf�֋� �B�}m�'79���v�H��V��{ICƝ�@ 7Un�X�����p��}�����e��&Y��@z�ѣ��c��Lҷ�r�`֍����B��NZ�c�a�jk�6q�3��mD��3���?��.]�M@�MC�W����͎bTR���S}~�;[~�.��0;(�$����R�F�#�~��\�7?�f@M�k�.쿞��ٹH"�<��|��wx��wb6�Ld[A�2N�ñh����l&��q���������>��Nd�xq{2��v]S�`�^4���(�Y"��l�RZZ�:y~��ǘ�6��`P�lzz>��ԕ+WRI�����-H?K~����jg��d<I5�4�43�9�S��D�Ӳ�W��\8C��"V��F^(�t������W �������y������N�H�w���MH���}Ό3K8|I�h����]^���M�%���N,�P4�����!l��Xg�Ï<<�;?���������t ��5}�������y؁�{�͞R��!0��vz���ѓ�����>ʔ4��ly���Ľ�P��x����Ʀ�>��/L��/�8���{�=��c��U�˗�2/�JR%��������ط{֥	]�,�؜�{�$7��M�Z��#)�Q�3����^T&+*�6�<>����b1ʡ�	�uu���I����y �)�;;�ѣ�I���˖�ᣍ��d�[�w�qG�K��x�_����6.�Ŝ�|���1KBR\��>�KEXj@�_�2�_��U�����h�̋��$nw�+pŌZ�,����٪�ᦘ3��G��+��H�.kS�WBO/�S	]M}O�*g8p�����(q��H"�ȡ�ˆ�k�Ác��N�P�\�?j�U'/X��P$~��}`oyiY�7�{���K���!����{��@�].�DwgW*��݇����'����1�l��{���������R���a&g>��˿��P�c\�|S7�>'�_���/�7ސй�ډ�-]�쓡�|�YKǡ�s�ǔ�x���ɌY�%��c%�Q�S�w/��e
�0�-Bw=�˘�/��3��az +�=�����%ɑ��@ss��:r�Dp���!�!~����pnD�0��G�`���ّ���d��|衪o���W�>��j�F6����
�N7fI��M�p����IfG�EltGf�o�dq+�3]�b��X��6`�����w�� T���ܹ�;r�y��JU��-nH΀ڐ�I�mB�k}�|s�&*t06�_</�(�(n�����9�d���8�~1*�e�R0����]�H��W�[����1��.++�B�^~~A3�ַ�;c٬Y���=��-�zH����X��ش6F/xVE�T����ٓD3�בH��"�+���r(���p�K�pM�Q�����~�?�;���7:sx��/^��Y��O��#�.�?���0�+%	j4N�Y.V7�ǿ%����Z;?����L$kq����B�[���1tˇ�-��0�����\���Q�,��[��'�m
^�`P�]��0���y�<�o��O�vP�	c_��y�]��>��t�`&6�П��}a-����=��e7Ľ��ڽHJ�]FB��	z��@��#�и��3�ce�zI�Y�+fz�z��4��2ױ��z�`@�л�Ur���Aڌ��LP80���@о��I�	�7�K�0�R������H,��I��9{��wM��oPߡ�q"�H�n(�L��N�� ���M��2騨������-ܲx��U�{���%8fkNNVD6���F�L��1cF��G�5k~�>�md{x.��}ǜ���hl�$�~�9��=~�y��
���Z23]�nؓ$�x�Aw�y����Ay��G��y�]ka엢
�0)%cF;'i�8d=S��2(x���9>o��"��2<�m�3����Ƴ�*q�J"�(�?*�Ac��(�T%���\YJ��Z�fM`����'8==�����g����WZ�o�7c���e��~[��[BG���U?��<�^�ГEIR%0[�Ygi$#�����L&�r��8c�h����H}�D/��~������+	���\�7gp�p'J�%3ݬ8m�c;����;җ�1��W]�8�$e����|pf-����_ �E��B<'q�s{����I3	fob��d\T��9��36�)��J�0�gيeg�Dz:1�����G��`��:�n�ү��N�<ySaa8OJ_�8JC��;���=�Yj�j�8x~��,�W��2�>+ݓr�~6��;_��|�xe��>�d�b�5<婧����������C�F�=}(MB�
��
�4Z�a�*Z�.��Ǻ��]=�w��:s��1z8���쐿9F�kS���y9�x&-755����m��~����(-+E�Zb댹��3�7�.p��q���3>�������U�q����\���tXgGw0K\��Aʸh�pZք1�	��Tj��,��w�ћS����AD�oV7��t�|��eZ�Y$jf4BD��:�$��7'~v'��K1I%�2Ȇ.���f�>]O' ��p�	����1=
�1_�=z�>_C'8��s�[�����z����7��;'��%k���9s�u�8��
L���ۛ��)ō^��f
q|Q��ڴ��U�מ�L�N�ģ�P����:���pɥ��9g�����y�?	m ��8@ ߻a�hӺ�����
#���@2�p�~�j�}�p۝w�����e<�*��d�0��AE�0���������/g���?��`Yv�c1� t&�Q��tI�!��J��>�PG�e�U��3>����<~��z���׭[�!F����H�e�@�x4!�i��&C%.
���?���೭�{�7m�8~>2�yl��"�璊z�
	��P5T!y�+W�<��-<�l�755��9�?,�\�Kr�0��[n�ܜ�ЭBO�I�Q�O�pk	Y�*#�����$~���	������v�����n)_�� �~cg��+o�I\�'s�9�I�Kh#ao}�=	ˌ�����C�8�p�������^��X� ����z�0�c���|O���_r�����H-Rs�m/q6'��ē �����R�c!�a�2&�.[zx����8ԍýv��!`����- td�dz��D�xvH�نc�9��\��է�;����},�3�%/.wY4�}�π��7�x��3��o�xܱ�ͧ�3�Ĕ�E��)���{��0!���S������>�$׉/zni);/e�KZ�'�8�ˀ��[F���GR�=k�L����%�$��������Y��]��Թ��,9�˅X��sW���>sr�Ȑ?��G	�vʩ�9�)�?���%���qW]���cFQ9a�F;Pr�f�t?��Cm��k�C7�
�!����?EI�TAa�K�Da8�$�G:p��2P
3�J�Č�C%;EftѢE���ղ~�^���Y�f����E���GͶ�_�L��������~?�Um���]�bkgX�>n=x�>f�+�{&j`̬WD܉/w��x��H��Y�~�1�2���D�F���ae���A�������w����N�Ap�[�{��p/\$�x�l����9���EH.a�E��H<�O|ab$���\�Al��ǟ�����p\��O��!`<ga|&��`)!M��)�6����N�={v'��я~tŲ������Ix.��J�3[��H��`����.��u6���1!s��M������r2X�x3+][�"oHD�����e�#�(i��t��m�c���\!WZܙ��p�E�6&��t�NG|eUe`��)�U�V�9�D��>΍�=�K7�������M��h�F��?NxD4'����k���ƭ�xCB_�a]�/��s�׃_N%Sp"ŧ�rj���2�DZj�� ��:z�b -�1'�BAkW���<�:�3'd�I֕0�,Lզo#�Cs-
�>��=hX��!+��l0�8�n�~���������y��+(��|bx�G!Ћ�ٽd�)_��W?`��vae$���g�������W��m��)�T dX��k��F_�ͻP�0�決�U����,���.�����)�		Ϗ�f����}&<=.��;ݏG��l�@rA�h���`��Q1oL��^�=g�b���|���������=3�IҗD|14�������!��bd����> ]E��d��7bZ���&1��X">8v�����oo	������k>"fZc��V�?��ݕ�UbY"��w�Y�|�駟Y���>��q��>�]�x�1��5�G��>��ϝw�9/#��uZ�z��_|���"<3�����U�2N)ؤS�t�?!z���>xq=Y�������#�S��'��3L)��ں ¾����yͲ�����Hܜ\�܋K�%<A�Ú��95��=��s5Xax��|���?����߿� �b��_sK�,�0����02A�_��д�3"���M�����h|��e9�(����<����.I��i���q7A6~�㺤�@x} �8ƃ��LO���X^V����a֪U+O`�d�)�3G�[��̥N/�ֺ�m�n�drV�q���A�"�Hz�<*��D�"UM�3��&'$,~&��о�{L�.-����a�j������۾�vį313J�6��H��%#�Ɣ���-&dl,_�m,^eI��%�ObV5%����Y����)� 	wxy� ��x�Z�ɧ�&�pq}��w����"�m%oۼ:��!�s@���Ϸ�]Bn�ӶFIOyyY�{y饗.Bө�c��d<]�c�p���s�ψ���co��}�';���?��ŧ�zj�ŗ\(%mS&O�k�{���]��5}�">?��I��q������H"�+��w�]�Z;�0!%�q�PH��0i�q�S�[��������z"�O���<Ȳ8hs8	Zr�>�Dm@��ѐ�\l���W�-�'�?1u��u3hiuvQ�6�u"��c�>���%�#2�@���@����]���j	���s�y8YZ��~��L1�@fB��UP�����-���<uz �-[6��&� ���b�P��^.�S�I�׹�^g���}�-K[��Z�b2r.�,V��olO�3��r��F�ei����� ���&����&�,w��W�S7�������a������ak�;��eR����d��������Nx��U�N ��*��cg����+4���|�{,�����\ǹ�\��@��T87��D�P*��Z�7����!`� H��aU���h��.L��{��%P����-����W������_o��|/�f�,|��,5~c�8d6J���A��|p�}�W�Qs�S���G=DW%4����r	TszX9���d�,[s�=����p�*��:n�j��heh���b���^}�����8Q8	�fx��c wv"�u.t*r�����`�<Y�ۂ,y�����l<?A����_O���P��b�������K�N�õF��񈮬(��78�����us`Ŋ8	�2��"&$Qd�������;;�_�0$���kl�d-	O���Z�Ztj_B w��H�W	�ǣ+�V�9�V�߼�����pQH��EB��,�m�O������2)pW�'��ӗ=}ʍA���?����+��ۈy����5R��E|��w��Z�-RN��[�Qu��ӕ�g�3����b���n��4���J��{l�y���%������Ip�e�����N-j��;��q[��%�tN�>�8��Y4��'>#����ʅN��H�y�R��ڧ��~1��� ������{��P<�ᙋ��EsNa�A:�?��/��W�z�����;�����,���3	"����D�vӦ��U�W���� s	�c�Ԧ)�ǅ�K���(/O�z�p�q���|fj�9Es����ˁG���E��C�(�_	zA�B�����vt��7�6m�d�S��|BNcF<
�v~�>�����\������YX\T��-[&`���K/-(��G?vDV��p����U�I�k�gOŠ�l�8(gEtgH��Ą���V9�2qs;P�7OИe����T(M�?h�/cǌ=�Z����J-��7:�uw���BbL&��JF;6��l�w�	��v`���˽tV7@�ba�1j)ۀ��oCR�$3&u����,��t<��~�(	|��P��Ju!^D�.Ē'�K�Kϐ���L�8Il���X��&���3=
���5E�HO�v�v�e>� X�{��Zk+A-�p!��=cU
,hͺ�#����5�K��e�,���"2k]&z�i���6e�<ב8�����}�/���?�_��<��&�S�	�ň"�����)�"$
PÎ�9����DiYy��8�����-ԟ���C`�F �M<��r.l1*�
�{��@T	�y�a���\��������:��*����G�y��q�g �\1����|��a�O����A��s�h������^٪A��(9�g|V2����g:�\ZM$�Dz2���-ə���z�ט��<�^i�:iR�V���p�Pn��7>�i����(��:u���=��|�r=�ڵ����x�bP��v-�e˖WttvN�'�����,++	�"�o���XLf�협��������tS4!�4�_�����0@�T&cv��̉�{��G"�Ij�[h���T�Xղ��Ǘ7)�:w�=cv �0R�2����+=P�5P��G-VN���H�Xُqs2��A@�V�����X{{�AvH���̙��ؑĴ��	�fE��!(�wb`4h����Sq�̼��QW�1!a�<�&�aH�ºd<��I�����K�a�.�4r�脃xh��~�G��3]诬���n�ZT���K6��^���N��B|���d<��d�>`��}P����rb[��M��`�Fxw��u�j�=�\TT����rMiyy{Q�����4��X~&?�����<�����������O�ӧ+dGA|?a5'������q�����|��?�����>ϵ|>?F��c���{��(�<>���g�x�]B3�4
�a4���K0�D\f�c;
b�9TC�K3,%������C넺�A��
���k����f�bfރ؅p5�vh�,��'&�r�k�q8��D����f��Blʘڠ��1�,NP
��ۏ��C���w�C��%t�ӮB��2fP����κPDq�c�x���J� �-�p��mװ]���RW�z�Y����V�r�+X-7�F_�\�\U}rc��2sV+�����k�����d�.����}/r=��RR/���hi�9M$����F��f�^�����*���5�s��gRoX�`\�[��EE���R�+o&�B:���P(�p{�@LZdN\X:��I�mE0Aභp<�w�p~&��.>�I���ZS��ft��zb��7��4h�&�6~�E�\���s�.3׭.�E�yIkDwme����"`_Ŀ�E��@gAp���4����p2�݄����ɜdg5t�^���rη3�^Lf�9�`���Oh��sMIi��-���������?���[,�w�}0 �cQ���Lu�^� >V�੻�D՟��g�����'f�|�Z��(B�.����01`�W$T�g�#ao��A��u�`����M����g2�|�q��8Y���[�%�b]���&'�Tz%&-k�<φ�|�H��r2����&�H�C[��3m)�����.)*AR]���JB��G���}u�-�%���:�{
*�*	
I!�$3�Z�C�~��ʵ
ш6��d�;2�u�䑮y�@tF�4|^ �K0$-��Ze�ޘ�@�e��=t��b_��K�=P"Ⱥ/�9�d�)�9&�����.c�B���M�/����u�/�����I�3���n�A����_�MMiS��ݤS7��D>��N�T��Z��=ޜ�X0˱��=E�ޑdJ��.nJ!j��r�%%$$Ƅ�P/�zE���FAs�����f�ѻ�$���+p�b;2՘���=/�-*֌�����}	�3\�߮���S��J��}iod�Ty93%O�C�-�ɂ��7�����%���\=j��/j�kM��0����� ���s�{���$�'F��y��tU��m���S/�����t�ǳ���2u:�}f��Gw\=�ݚpQ�K�5�N����{��(f����Rk';m?�X/r���f�7����"�U<7]�4�q�%y#��򕯼����+V]���,?��F��)���2c@]6��i�H^Cx�����i��o���W^���E>�%���K7��r&���g�� �p� �%�|�#\��>"]�WfL���8��[�����9��+w�w4D��*��Iy�$��K&p�����KUxΑ�cL�CX���H����Z�vu8��Z���x"V$�D�)/�� �馛-͍��t!����$��i	:��t�r��0���
7}�\WI��,?���;pO"��0\�}P<���ʘ�ħ�����p�K���������.�'�	�yT��ttEt&�-U��:�u!�� >���+AL�Α��a��<?w.���J�������9�y�ii��nU��rʼBٸ��ɠ:���7ryE����U*O���ꗄBzJ8Y��3?��k20�4	�e㌒7�U-h�Ǡ�R\LL4q����"�/�'2�v�{�ny������d.b�3���q��I֜U�����&n�T��É���u6������_ �|d��<�e/���i�˗�'ݯ<;d=u����f�|[�[	�cTb���!�������F57;ջnm��ů����RZR��B�)��}KIq�k�	xb�̙�h:�u��X��N�c����X�c~�ȶ:��~]�G�)����I'����w=��og_�g�쨔�_�!�J��w�"a�|��$�#q��ə��t���v|��)��?7#���z��L*�Qń�^��/�/�'s��.�vx����埸�w���ʟ�����\3F�L�D�ڜ��͡W�OĐu9W���A���/���o��bN�J(��b�k���]B��
�^99��cZ�7��)����0�C0V���#�pP9�BPz�=!f�.Q�W��)��I�����	Vw��
hq�$Q@jԱ��n�U7/'�]K=�X�?���	.X���:,Œ��+�k�x�;{��O�^��q��}�et|p;7�'�m^��$�m��e{���`�_�tW3aC,T��xk|�.pƄ�c�c�$j�]�����l�1v���p��f�+��y7;��F.ښ��=3t�.��8����2dB�ٯ��(G�-P�{�"�E����V4 	����Dy�"͘�&nn�@�\\�XG�9��z�Q�=����q���BiF~|���T�[�M�|G<�5ɘ]�kÒ?^u�KhFn�D������d�{�_:��$nן��+�q�����6�T��������_xa=�vk�v\�R��̘1s�A���3���ʃn �c�F �b<o0������s�_3>��O� {�\���}^�7���?��w�������.e�v�.l*%���G0轋Cp�a�C��j&��h�m�	����]���V#��Tz99���tѿpM�<B�;�ţ�]�g�=�ܿ��y�_��;Ϲ��ۖ-[v�p�q|ѣ�ך�R7�ls��<1N4୐�Mu��T��*(�՗����՟�7�v	B, ^G^(����֯� =�S��W�;H{8Z���X� 	���jxA�1^h����g��1�{����H��������+�{�º�a�~����k7J�zIq9 q)�c7���br�Ȏ.�1.L'�������Ru5��9��w�V_���}z&�K}"�n �*����]��tP�D
�ˈ�	--�K�̒�_��>���P�X��B6�+=F�2܈�^&�QdE��[��-.�[o~�1�k�uV�3_u�3�A��De��f)�\iR�8k/5���
�-z��+��uĕ���"��H������Ǎ�t�Iz��g��)�$��='qlX�/U���#>\<��\~q
�����].�ܒ������p�E�9�%W�'�H��Oq�I��(A��a=)0��O�K�l���
'������$��-�[��"�B,������3c�rmo�|Ϧ�[�^~�����{��K?��ێ<���s��m�{��q�����yP6[��&��ԩ玮��e�02�Jr��E��y�M�|�/����z���+��ށgi��h����Q�B�'�B��c�nu��bO���|�37&�
r8n}I@s�u���o3W0 MUX�P3���1���[�g,y�Kcc�3g�����e����[o]}�1��1����	�8�먱rT����KQW��C�}�W�f�w�b��m̄'����)���/d΃|��en���}	�����s��.L�k�j��Ƃyf2�Jq�����24!tU(�Pk�5AN�����{ᩆ$�t,^3�t�Eb��cx0#��-ؠ+����s�4��#��B�C�?`���!s����nD���zXw�w��3��κ��uH��^���6�s��mP�\n(:�$1I�sV)�M��yuwG$���~���,x��EހX]�o�N4�L��������ږ�M���%,�e�
K(a�8g�����_�|x8#�rC�.�g�w^=��|$	o�I��,Z��	�ˣ���C�<J�bH����y]�.�uB�|��eϐ�s�{<�:�F�n�-��鳳?�>�3g�('&��GE��r|���L�J����c�t�쟓G�C��qF��:q(�d����%N|���s_|��5�_ݲ3�u���;l������s�n��]i��<g�}B`I2��	�E�{0`���'KK˨i:�妛������5X�Ѷ���P�&��|����d���]JZa�"ܚ��4=j�ۂ�$���m��=�d�?I�|�J^�����,_�.���g0����&�1����I�'���O��O|�ï;�w�����{o���
�%H".�s	^>�0�:L���1�EY�Ao
����PC�u�m�U���p͗b�f�{{�x�A�fϞ��ם_O�2eJ������U��~�Pr1
���&	��x%ሃj�\e�9�aJZ?\I�g� ��@�<�A��iT<\)? �j�u��&P�|/� V��(y�]&�PY�t����M��vc�n!����&�L�FZ��S����B���Ar�Ĉ�a�!	�8�&�;�?����V���Pt��@��Q	K����	M�(,�B/A$5��5f��S��s�K����Lc�Z2�������{��T�qX6�P��Q���������#�C��H�^t'�� g���h�
���k��ϊ�d����}a;�ϟ����,�k�!��!���xn�Dp̶/�EH(��c���/dc�}�Lc�2OQO��`B�1�^t�9o��k>1�Nx�mai"]hF�-U�2�����'�|���r��5k7���{ֿ��s���Ϝ{�Ϙ��8-hD�Sm�`��C �c%x���~����0>CX���_���ћo��/��W����Ճ�ùУ(�w�=Ƀ o~����4�fz�y��D���yJ��K���[
�1�{|��4��K�Y55|tL��Ǖ�19�4��1�/_�F��W|�� �ma��}��=_�?+W�<4���6����8���y�@�U��Ti�����\��ҲbI�+*���N_�v���g��O�[y�"ۺz��g�Y�ھB�Z2*E�����/��,��܋� ��|X�y�.�X�G��|�$o!\\������*��:e-ZB���2&��I�M��	�$�%�/���.n�x��׸8ף���P���s� ��]O��~��LO��,80���(�X�襮O
|�')�����9?nFf:ϗ�)�axG�BV�6���X�1HP�!	Z'��&M�(p3O�����w�g깋�;{��_�cӥ%nx�S�$���/��\� ��/,��K �\M�ć���0��Ϗ��H�	�)����zޝ��N�$�E+Z��Jz��s�����5��{����2y@)��q5�E��ᗔ�N�ekB��H��P�����Q3�zE�e�{=��J)Ӥ�?�tC���B&4nR�@X�w�xi��L��K602�$H.�'���pEP"��BRae_"^	�ȃ^[���K�}֗��-��}�Μ}�?�����}λ�˜��nC n�,��f{CȳD�X��#a7��s��U?YR�:�^S�sA�eo�+�]tZ����فv<ǘ��ۙ+y*Ո?3јdLCP\۷���]D!�V��k�nK�/���olX�^&�|O�I�m�w��+>u�O?��On��ޟ�7ߴf�q���ON�\!	x0���AW:?.�bl��j�*HXϰ��2	g�S �mk'b�U��a{����"ٮ�d��5A����Q�"vy���!<��łHt�U��s�R�Z��:�&�Y��f-,�R�O¸
W��ú'V2Í+��zp�:"9@gy�h�Ei�C��E�6׷�s1�I��8��J��|7�������o�r͸�2�[�����x_��:���b���ū9����#D�5领�-ऴ�c"`d��[��
�#���nOX�	���'E-�Q����g�K�$!/cL�����T���2�A���QA��>��M�S�t�z��D(5��f$���cN�8A�9I`q�nՠ�<io�J^�Be؄�;mҧN-7�I���u�{@�9���z��*�/�p�g�0� ��}��P���s�dn.��A����r@�P�K��1��1t���3P4�o6�C酰>f�@3���A2����p��ɛ,�=�X�x�'�����z�	5��B�*s��;���_r����>P��?����8�'�Z����w�}��s/�p>2����{�%�g��Û}��sC`(���^q���&�JN�xAy�:%4�H�>|7w(���+h���㏯�w�����ӟHd�
GVz\��+��#��x~� �^C��u6�A�Ⱦ�݈�0���!N��qR�E�>'��w�Ir�yu�&p�=����}���4�.��G����?���<��U#NJ8��禪���|�M�����\ /t�����{��I�8']�����f��X7�ӊa�Q�����x��B�S�uww�����`�a�����5Z�	B�U����T
�)������A�]6o�tƂ��xa4+o�>�������+�"Z��P�R�Y�b���1p֙�W�MW8��H:�Ə����+ȳZ�e��|��\�p��m{p��aA"-RZ�$6Z�L
��L� As@�d.z���X�AE=�j�=;�q��a�ɜ���̐��9��HV��" �(I����$�}ބ�oL�dh�*c~�s��$g�h>n�	���2Q���q���cẙ�_�.�z���Ӄ��-�����nL?���k�1�\�������ߑ� dNvwt`���m�ǃ�$'�Ԇ��$���$���ᘅ��øf��n-���c(�k� ��g�����}��s���[�86����ޟĠɎ<�MB�|`-�#|���3Q����j��rȒ�KN{�W?����^|���w�Yg�����!=|��;o����fr)n[�!������x:$;���\�p�-���^�_X��x`��H%�H�|���(īfB�4��3��DTgk�s�
�R�+�TU��A�	uKk��6B�^C$���+�&��<��u�o�3�/xϏ�ӫ6�N�ܧ����׿q��?<����È�1[��LN�d���XI�!y�x����aULR�E=���޸�L�C=��׫���'��죹q�(X�� ^!�X2Y�!����a>/Z�b�;��+��\��>��<�h�t+Xf��L��� ��7��Ck1���i!M������-b����e,ĺ�k��W��<\,l�RI��-�����_��qC�7ԋ�;o_
!=y�'�Iӕ-1�� �s{!Θ��\lF�W��%qq`��Սx0���\�t�8GN��3���L�B'A	�t�;W=�H<��+g��{]X��=A�ƕ���}����a=?u�s���u�M������~�P��s�M��`���ɁFsnK[K^O$Z�Y~p*��Έ�11���X�{�׫�2��tJJ�S��1iB��>J)�Ck\,wu�����C9ϸN�D�
�.�^��]����$D�W��f㞘��]�|��w��=O��޷�p�	�;�̦᜷�kl'=��x�e�gN�x�S�����}݋2�&t�㢋D�aѕW��s������X��
x3�w�����uI����U�D]:�8�9I/�E���0�|��ۍ�#&a�� O��~ͥ�����ַ[�{G��G?l��}����U+��� �����#��'�x\��"[D����gwS��$���lK�ݳ��֏e�}�`T�L����7�c|��/����l����&H(��J����$&�`���q(��-�\DH���7ez�^l���	2�3/�8�IZB8g�ޥD��d5 �	H�a�!�M-|����b��#>t�c������0H|8>����u���:�����m����omxH�9Ȥ�D/ƚ�2�.W �E�K8A��f�k��b�>I�T�SB繐���B7:�������L�s)g����M�A
<��P+��$�����^���p�~+����ý��t�\�A>P��3���QRz�7ea�8]^SsSbz ��0��҆��ٍM��F{z�0��T_�D��<4J��5Q��:�r�,��� f2��D�r���1���t�����`<3;�����z���G-Y������?�λ��ǧO�z�	'����w�%��;� ��\���\ͷ)�=�5�[Ҏ��a{s�5��}�mx�֋�{�����{�}z;���Å^��g��a�����j�&��+ߗ�L��(�!;���{FMI4��Y����ԇm둯���Y�{��/z�����&`�9��E���������B�k&�pb�3B����B⛐��W�_��%�n�n�T�KA@��;�a@��a�[��[:�shr���߳�:�����ys��k�{_��Z�����}���3�3u��"]����W�������}sg]?�6��K�}?��T�M`"�(��l��8���s�ɷ�PE1�<?s��}Y>�x�eJ�8�C�d��x�w������;ų�|�r(.Y4`������o�N�qS����z�spG*��H���*��"��G�@K�����o��{L����6iA��qO-@�#w9fZ��˔&jQ��D��HϽX�B�̹o��x�\x�W��+,�G�Ӧ��o��<�@�|������ތ�x\���՛EsL��S1Z����=��U�s�#��\��v(���s婊r?�&�[�?��
���C!�=�Z����ZM��K��#��l�0M�D���n����X ���f��i�N��mu�w"�k�b8�����vk�u��؃�q�Q���%H0V�vi�s�-�(&����#���@x����?m 0�e����������IJ3Y/<���iD��W��):e�2���75/��~�%zu�����,/����Q�%%\��A�x����E:�����hŹ�^��I>����f̚[V#X4�v����f�M�����ã󱡤c�O��,�nZ+�=��dO�����T���o�:�]�����J=�<4s`�-p˺�7	��qh.j�͑a��E)�B�N�,� ��ϊ�z��r�EU'�_����yשz&�4�����h��s5d)j���%���'p
F�J��x�����>��S�8o��	�L#E]�s��Vi�N,�Q��"��kF��(If��ٝ�+�_�)��d�]�Ps�/���J������/��J��Z��
��ejk���F��!��v ���TP�:z�"�'��6<���ׄ�lu�l=��(A�����Ih��{�5 �!35M~��bW^�v��T���������0:J=T�f����P���/[�~�L�m���ذ��.u�b�7�[�O�\$��DS�(�]�X�߇b�䔥�l ����A� ���l�\в谺�1���ӻ"�US#O��#�JI���P�rSQp�Ơӿ��[�.��Ha�n�6�9OG%���ea�S��}�P,PUkg�Խ�}k�A>����ܑ���+懤�t�\����7�?5g����2
_]�Q���@H'�A�Չ"�˿1D��/Zx��	�Z>�]q<5�2�&������:k"�&��w����2l)�)Et������|#ҭK ��>?���;��_�u=�'Mvuc�qXf�B�V�\�/��d�L�Yo]�EJ�;�*�$���eB-Ea�+ޮ3��+��9D �������=)��?���Z�7crR���A�wW��'{�vm��N�	
�XF~��`=e�@�C ��&��E���V�o��f~X��[!�	��P�ҕjxn&SUX���*�5���]W�
"��O������/1�o7~%g�:u?k�D=�-8�P�P_p���i;�^�ϓ�>�a�����O ��̣�r�p¶2KH������8}�]��I�#ۖ��1ǳ�w/ۤO�o=���ƕ�ʂ/��*���F<���(��Y�2��t������|����%�vQ����i�n��#�'U>�CܺQ���t�<|YZg�0���ћ"�g�D����޷ˎ���3�#����j58Bk)!p�9���-�2~�b"�ן|mU��D��8��f��ņ۾ea|!�e�co]W@Z<z�+D}��GK�������ݔ�|�F派��{2��%�jc�
�M8Vl�*X2u���(��@߼g �������|V�Qִ�HW�)����bO�GH�E�aT�E�N
���6�W��X5$��+7lY�<2D�K�8��YI�W�b�`��|C�{,�y��Խ�Z~j h\���ik��z,�C�5�\@��߀*�`�0���>2xq'}71�� ƿv��T?��Dz��,}UYD�5�d����o��'����4���5��P����Іc��qx�|;��+��.�L0�>?p���{н�K9eM 0�U�:�HnE�v�;aܰ��b���q\!�;��f gm������|�ΙN���ˊw3��cm��9���8S�)���(^H망by̡�F���̕�S��|�'�ض�zvT�[�"-�W�/��.�5�����4��R����5�Z3H�/<ırwB�I�jXnr�.�%�kH)�{�I�����5��s���*��O������yy9�O�"{g�����/�Lu����1����k���k��~Y��;<���������EAĈ�;q G��/���C{}R�$m�$K����I�I�&�8����O�>,���,�Ksפ���o�x}��դHSF ���s�1�7��F��E{�=�F���Q�Χs�'f ͥ�� ���ՄLi�=��r�q��aK�� }6�伈|�;h����"�x�_C3�u~+�ݓ�~�����Ա���l����`����k���p�i{`�ɓ*~Y�X����J�D�0y5��&�%�&Ss���lu�}�/]�@��:/�k���tE��%�V�~2Z�t�3�G�ŉK���6:U��U*��d�S��
�C\�'~���sjZ�ͧ�].�yN3�k���u6qE&��	�GT>Vj���t���ei����̵�!����n�W�5�H��و��E�Y�S
{�y�#��H��Qr_��[�zY����N�n*T�i���xUԯ[��G��yj,�\�G%�o� ���?�g �K��5�1�;uA��2.��)#��?��)�T���.Zq�3=�,h���o�&H�?�jI}��S�Z���+�)�,ZaP �?IS�ɷe�3D.E��r�B�G�㝨����r2��S�u������j
�x�X�����F��)����~b���W=��������5��$�kE.���G˥fx�~j���.z�أ?�5�E-��YdT��%�뇖��WD�KHA�Y�CO��l�ca�Q��w���p�b�}&���[��.A�Em���Љ�nm���ܺ�ZR��2����g�G�B��W�k�Tp}�tC�䲒��r�w=�*�YK�l������{�d�Y�8ȫ0�-��wu��,��$�7��0t�6_�����T��M���ε1�;[��>6����2ՒG]�o"I�w��u���Ys��Tȭ�_�ic� ��nu�X�9�L*�k�� ڰ�N�t���M����^Φi�r�WոW�vǸ/�Ҷ~��
G����aj�q~���6��_��~�}�'E��L�B�1��E)E}9�lܪ��ؠ�[�ݎƁ ����Y���?�#EqF �	�,�"vv�M�r��/ �����ɔ3�s�
<N�K�ks��l�:����ig9�uܼ�ޞs��������h��i1�<�=�$vמ�.Xg��]�ݕ%&�Ǔ�+�Mg7��-g���W@!�$�d6�2g�k���A;7�O�h5Ѱ�������K�Mu��]u2&��+ ��ѽ�O**8�����k�/�+��H���%�N�i�;���<I���������a@���(F2�ѫg��¿_KSmb:@�x���,�����֜�Ԋ���Tzɏ%�"$I䏭F������,��i~1���c:A6����d��"���F_S�����o_s����ύ���&	�wI"�
f2�k�����
&D!���ë�%�*�ܻ��o���<?�J�'T�&y%�&}�_eBR�x������WK������<�Fb�r�z�����-]���P�����\�Va���c_��x����%��0]��/����oU��]�֕D>�E����KMU�Ғ�v�Ҧ<z}Ӌ-������S�I'ZF�v��N��~���&����Dܑ���3D�p��U.QI��[�+��#���f����$��2��\�-�&P��]2�޸��{;*i���J� ��\;y
����q��|����Moܳ^��O?�>���%h��됔�E6�'�\����w����JN���ђy�/�(yF	�34�+�O�_��բ�#�UG��Y���̙�N�oS�L�BG����vgXEq��nqG�p���o>��8{fy�⧊�x����0�69Լ�;�Y��ʂQ=p_x�@>�@>�Ɣ�ޚ�Z�-�&nD��Y��m��4�}2Sl�t�'*h�WrXT*7
Da�]S���Z�33�w9�+#c�VI�B+�o�p�%Ǭ��X=.GK�:]�g66��J#���-�c�M�Ὀ�p �s#�	�Z��w<*+�w[���(`v;w;f����F����]ւ�+��Z�1���2͗�7�����,dOwi�$���ӉG��
*96���Tid!Pw�L!.BY��I�P�]�/���jkh�S�#[z��4Y������_�0�t ۳Nj��ߴ�_�^����x�p�]�ts���^?Ǘ�\}�����AS�H��$�q@Lq��~�����M��@7������}7��d�����X����,�`��֊���ӲgU/tV-"��uSNS[L� ��Q�����T"u7�+����������N��L��k���`*bo�� �>���)�	#DL�y���̤M��$kA�ק/
cQՈqK�>�ˍ5�U��f����qM�@iI�lKQEV���膞���?�k�[�����TER0�=~l�q��Y��((���J��{r�;�e��u)���us$����������(���_D�B�gv�I��9H�~+K�(c�A8�b^����ESբ���o������Gt�Ź�w�Е'ˎ�9����?șq�H�_�U�GGN����/�Dؾst�AST�SuǮt�(y��l���b��D�B�1��;B��a��=w%1-�q��;&�v��bS��L�g�!J��A�`>�5i�u?�Ɣ���[h��j��O
�Gѵ���N�jxK��.�Y�A1�,�Q�����]<�uh�"�\��Ӊ'�*p��ϟ!e_E*{R{�%�5 ��9�FsI7Kk���}B���/�#Rv�'�K���-P����-���z�ァ6��/u��O���"�c����m�� g(�I�)Y�����$��'���Q��D���S<�4�;܄��+�_�8�ߐ�/�<˞�����ބ;澂-n<�/����6^`F=z(spj�.ٛ{���Ы�h�Vwv�rޯ�z�<;��<jI�]�i7���Cs~��q���!��9��Ynm�����"K�;�/�������u뷇�N�MiEZA�ٙ�#I:�����$�I��}��ѱ#$x��'��,���v�Ӱ�����~�i�0�|����KT*�)�9���;3�}�Ï��c����mv��Y��C�9��ydo��&B����y�����ȶ�s�<�X���&���QD��ܑc��q��������wt�^/�	� ��13<�ׇ�����������]yL���K?����B�+�#��W�Q� sȒ5-�ǰ�q�T�-�!B�M�$'�M�5>rS�0��|[� >gzYܢL��rL4vy?�
�M�ӯK�X�d�K)���l8��8���%b����y���2�Γ׸������2}K��	�	�=��ܳ�����r���k�Q2����k�M;q
�ה��UW�]��o�YԆ�ӣ[�#)Z�;��"{ϔ7#M���K��}���
KG�z�0G.2�0�����D��y�_%ֲ�]��#BAE`��8n �c�@�@�j���a�`��K���y����.�yP�4́���%j�^�층�x��D���[��D�2gn~��~(/�Z��Mã�]x>�X�� n0i����Q��*�5�V��o�u����6 �ϘaE���!gDª�ٍ:��j{�V_&T�n-Y��fU������ mfS@� ���N%Q:��C���RJv���V��Ϛ���Y�h�-�x����Tc�--��m��D�)m	��T��"(�n�ݦ]���%�\:k;��(�Z�⺒J\�<�;���e>$'���S�v^�pԶz]�������i��
yM+��m����d� ����v��2�'�	=���Le4��R��:!pރ����8��/�q�
E��&�Ƌo|���0��6�߈8d�a_
�4�?��l+�p�g��'%�l4k�ٔsEO��^3o`��gVVb�'��,rB2�T�>u������=�͆�"KA8��2����X��h��)�ԑD8�]Jd���T���_���S��$d��Y����Ş�{�6�F,�_�Zױtj��k;�*^�w�僓^�+~6�>=��}ڧYY�5�쳬�T�p\UYY�݋Czw�1)�Lʖ�{@D��,�:,>���;�: ��S������B��N)!���v������6 �,�ݶ���M�v��oN��Yn�|��ɫ��������$�pp�pJ��Z��~,�Q+) ���kp�_P�+^�%�-P�m��^'�t#N�3��hu��
������[N�c��T�}���8lE����35_��˞f�X���O�1y�����V<Q�i��R�릸�k�:D����m�z�]�>2�6��n��.�
 ��"�WR�K�����:+�]0��@�J��OM�f�V�~�jre���gH�\�v��%����In~:���8*#M�m�}�����/��:.a�Ido^u�[�D��\N.�ïN1V�^�֓K�J���s���G4�#v�]�~k�~_8n��U�m�����x�ԅ�h0�vn/���'�x�Z^���N0��,��7���ʳ)^@-g�LE�j�ؐ#�L��ا �B��i�ɭ��i�����r�Y�_��;���fK%��W��ݖ����Բ�2��u��ߔ��>�����Ԡ%���?9jo��?���.Y��<�=5�&{0i�)r�gC�^��eXt�`دk;��⤚vUU~��[�A����W�e#a��g��'�5��0{�������cO_~*�39ZaX��Y#��Qek��z*u��D����to��T�t=xoC�A��jl��f���-o��r�)�����5�A����=���v�J��ӳT���#�o�����n��1Si���-�>l�t��P�(���U7�a\�+j���u8�����1���f~��I���2kK,t����d�_��m�:_\XX@#BQd�4��$,�ר��=zV[��o��F�_��2tZg�
I*�䷀#����s��yb�B�G��F��mމ�� 𦞩��y�T�U����_�G���	d����ff>��z�>*�a��M����� �����l�z�'ʃ�pԹ���f���CW�pt�B��B�.���m�A�[��zH��?�ݟ0�"2�2!����&��O�g�.+I`Z�~�@��fp\�>\��2`���Մ�T��$AyM΋��#�������ʓg:y�Ttb_���m�U]N5V��h�s�h�\!""��Ζ������^�2�h���#�b����y�~d؃t��Z�^�q�d�3Sߗ�������^��6���9���L���{Y��7�;������t��Q�����@U�0@A��������(Ia%I�	��@xl.Q�Q�W�K�����_WS�M�?٬Ǫ]���$ZJ;Nf�f���>����IÐZ@�ٌ��N2	�����(
�r�T�.��>'����kx�yJZ�b�2��F�2Aȅp�H���m*�)Y��ű��G�;&
�)����Y��w��~G�^�'uqO�XA���^�f3�Ut��|O;����-��3W�בo	����������뾋[�5 �,lpKeP���c�ɕ�wɗ��!u�@�����J���(sę��s��G�O�U�P�������.�*m.�ܿ����h���(m�ọ#aNK͑Ū�#��iF?~�(C�n��{������  Ȋ��R��X�\}?�ʣ�MKś(�=��-�i���4,�u3!<\PQ���Y믣��~	�llP�yV�3�I󜗟H�2�_������o�o�%a�/���*�s�>fx�%ȝ<�E#�-g���5����u;V_���+VNN��ۓՏ������%��F�g� [4&[�����yyl�������`�P�8�y�_��<�E����{���@��j���)��m���� ���Qb%*b�V���	-���ڶ�@_�?-̭0��߾A����۾���=�S��C(�؜"�Ϯ���̬���*[~6ivj��hsO&��I�TQ����p*5Z���Ŀ��-�b~xnv�?��'�nW+�?>mї��ӣ��π7����ƪ��I�8K$ r�?�A����_R�)\>7�(/O�X��0�ay����i���'U��bA����iտ���ArFX�Gy��k�S����Iڿ��7DH���	�f�ޭ��$f�s��i�ovV@�*���^V�񰩌s��MKK{́w�0���/�o ;E�"���&u����"n�y���Md�]B�/6�<I��_S����|��QB�t�И$ɸLSI�8Տ|3�e{���� �ɛ-2���oC'~ڟe�����=|3t�6��� ������K��8�O���Q_��x�ɅǸ7�O�W�Z 2��_@pR��ۭon�y�C�F���aͽ�=���>��XXX@L���y	��Xgut��Z�U�VMs��3�������x��|ƺM!�T�./b����n��6.M[�*�3;|�PHG�\�E['֩�h�['��$!�����0�U�5�B_��7�ց!Z� �ad���KC��@ ��\W�����p�)	��Շh��Ɠ�|~׸�����f��z\P�67[>OynM��� iA�Dl`�hA���8�0n�\O�w��bs^M��HJ�z��(n�[@b��]�����Q�m�ᓤ��᲏��R$��ɰ�j^1�麐�֛��m��a����	'.��v��\���qw8��~-��,�����z�����[e~,(���u*+(�Z���H�L�v1�����,�G��H61Ƚ\20_eo�ԪTј�_�"��5�'Ka�>Y��0��[��LA��sjR�X�����`-��|Ǎ
*$x�E�/{\��$==�K6mL�/7��*~|#ƨ������a���	Y��Z\�v�����C)�ן�o1N�?ӂ`X��7���'U���^
&5�mj�4V�<�%R_��5fʪ;���>�.~9��m�w�����g�c�CTr�@��,�kJ"�"[K��Q���
���ʓ ��	����@f����*}�z�ڞ���B^����6j��4�����es���ߖ�p��V��ۗ����V�H�4��8�C$Ժ��(�_�p��J1Y��
�&d�	�v�pK0\��|a_�~$�A(��!`|�?��!�>�s,T&o�$=$\��ej�����ʹ�,'�#@����m;ȫ)K���T@�j�;h���-t��B��*ⳅ.�h����-�q���~?��2>C�T`�ax�T��=F�"�����֠�d'� /x�=O�~E�?�ɻ�3,��Z����e����C�X��\� 6o�� h�J�������As����a �Q����Q�H��;�8C���v-�;��������OX9���y��W_J��f�i�h�M���>�
̫|��e�DK?0�vCAq ����zT��m�&���*�x�N����&dQ3��e�
Kk��o�P�,��~i\g�B�n��d%���5;7'BPlB
�1��W3��3lx#�+.ky����|��Df��43�1�5��@HP�2��U0�ń�Z��E#N[�?l]�3�ݭ㟷T��e�7��aS�EO���U7��,i�|а�SV��Uı�<����S�.��P-HW&���a���q��3O�Cɾ92���z�����-��^j��=J<����a���#�ȑn9Dl ��+�{\BJ\�+Z��y���� �j��^�=\N��1%L��M�{�
),�T�����Є��[������m'f*�/�k��@���)W!+%�U���M�?������e)	�qʘ���y��SW�zS�d��PK   �cW�Q9lpz g~ /   images/b53b9fe2-18b9-4e15-8ac2-a2240bce23fb.png�UW\��-\��;$��]���$�{�.��Ipwww	nU���]N���������\����jk�1����75YTRT  �!/'� �\�� #�]�Xڌ P+m���䥤��\�,m�-  `vJ���Q���J��La�,,�
�rp���W��hd�h�h�VB��h�f�:�%��(����� �֧����<~��i�7��% �I��|d�k�[�6���J+���Dz� C���j�.������q���}{}鉎�H�B�J	�'N�H�p��Α�:p:�w��Z�+��Cy��==�$�3�/O��6y�1`kL$����W���0&G^���l,[o:��/��'�M�-"�|�!0�Q5�K�te��#�P��V|�ٽ���-K �d��D���w��	t�Z�#�x�W��wh��f|��"�&Cׂ4��.�v��ߗ覟q�M:��k`�F{�{Xب��F'VD��p��:���!�9P_)�w�y�t	��n�����G�����K����*��+d�Y��?xv�i�^a�}�B��VK�m��tyh�|OReC3۔���>�k��W9�0j�n�r�^�SX�m�Ǫ\8J�!��<x	t�Ӊ�D���Y�����~9=lAՅ
0�
�w�m�(����5�l ��R9���a(�a�L�'�j��{)�p���?D���P��2�ň�`\AnQPø���@��ct�4�]�Uv&�w��21=����e�Ƙ��6ŭ��M��C
��V#O�J��!�F.I��|F9���%?i��u�����5ɧ���'�t��!���(�AI�,Xla��~Ȏ!3�[��(	���0��kum��PT���j
�Q�ɵBm%�~	����.`��#�)��a��(,�M~P�0���d6���]����H4�5�I#g*1?:^��0�0��8gS:^zLzGz��/�Do��Qm���=�'�'�'}3�/�z��@����r6�4Q��L�Y�TkC�Ak���JMd����L7y v b �x��0<�$�G	]��Yk��k�Oߘ�5!q�HW0T����fǥ���!������8�Vb|"[��|�h�W4�H�<��5�P�����=Ejt�N
"�����mޒ�Қ��;L(�ڌZ��� �"%5>mKf��Ӛl:b�~R�Q
��j��)=h��}~�$��Ԭ�D�S�+qUۏw��.�V�W.Ѥ�Q�aQ�4�Rnw����ѿ1�1@(�Q�pN��z�Z�6�<�@�q���i��1ڴ�k���X�;�G菽�O�:��G�,Rn�N�0RZ�8R/^1;.��y~>;�%I;=�E��&œ_K���w$�$�����|;�H;�yp����������Ð�D6�e~-�	�hfnI��SX��H��.+c�Ҥ�;�������Z�FC	�:*:)%.�^�|��:zd�u�%+9����%I	�7�����׼~�pu��,�q�g�|��dhr�e�r�4^p)�"ײ{���~��w3u��f�f|=H�i淌c!M��Q�z�u��rp�r�)���	��e|x�l��9�o@���ߌu��,��T��b�ruVq
P#��l��lt���������?Y8�^\����%rd��c�~`�2fռ���s�����Ut�qlj�u�t�DbA��p��f79i�E#͘'Dn$gl��kB��CW�>�Xϫo(M�4W#Wj������Ĝ7��Իa�i�s��RT�1��^N^"�aS����Q;G�/�<6����	>���mEm�o����%.����fY�g��Ȋ�⇹J�G�arcL�>y�y:�l�������EzIϾ#�!�R��\�&�%������]Go��{W*�F�ع��jM���9<���x��xe~���>�E�fY�O�>�~�/�)3�ˁ���}.����]�q'~�T,�'�Mc�u�1��D�<����L��~z�b`Qr	�7�_
�Oz�,`���y��3�#�>'A!�*��q�-v<�1����P�݌��Z&/F꒥�*Z��둜���%��ǥ����'��s�ϩQi�_l��������ى�����/]�^�C�)��)�:�f�F�k3[�n��,�K��6����O4[�������j��UJ�1<�5���^��~[�X���c?�?�~�z�9�j~�������{�Y 4���QF�<~9��7�ho+�:�Q�l���R��A�NW�\f����{˞�U�WN�ee _���V�;H�=�+ġ�g�U�ڒ���b?vO'���ם���c[�vEs��I�E�C�9ܙ��R�ci��Mh�U��ʝ�b��@�O��8�Ҟ{C�(=�Tbk���ۭ���
���E�S�S�����I���A�϶/'���%�*9`�`����jg������yP;���s��p�3�uav�/�~cosᘞ#��i�F.��L'�W��v��9�y�S�-x9�9������]�k�'��5�NO�n�H��5��WG{A�/d���s-ғ�v��T�uEeJ�"R,������j�l�r���k9����A����#Z�zn
�ƂhK`��l��A�7���xL�����x˚���������es���E����ݎ������� ��҇�^�����<�OD�}�e���M7�-��$�渹���Q�a�ia�-�� k~���z��g�t��<`�a.��6���*H�	P���Q�d�"�a��3�s�I��x7D�U�3�.)��Y��Y���z�Z���N�'~�0��;��{��  ��?�O���-_�'o��>P���0�o�;<�Giux�_�
�j�!As�>Gܑ�=|����OyW]��O�(��(�m��~�?�����^A�ؒ�M
��Q�ͅ��W,4�Ê���nj�(000�l9F��/Y��t���&%r�������<||l���X�Ư�'5y����b�ν*$��"ߐ�����?��KE u��ݓ///�k9>��V(�U��P���tiU�B��I�ull�A�?�A<��i%���|�G�������uWUY�	�/V�D� MV36v���spTVP�fg}�om����r����,~"���J��ֱ�����_[[����lw�fccӵ�����v����|V;���Zk:@%����
���+"�	���OOP>��2x���������Tm��i�R[������J�Y����>�c��:��&���tț\+�Wn�nG�����@ ��鮧$U1��{�߱�}
�VRR:�����v��I!�~�n������5��k��_�|1��[!��)�Ƅj�a������z�&�����w��819I�~�0�����~�^)��)99��ݶwЫE�:���߿��.Q[���;��T��m�����>7�G�{銽I���ն�Ѝ�5ۢ����r`P3�>�kū���n��y/��c@�p�4D?����c����k<l���U��KW`G�K���YUU���X{Uyu���%�g���98�-����aF�j�>A�R�I�Bk�Y��ҠRV�q�O𷊛���L-��ϗ�V���?�j�{L"�?ő����tE?�_^]9�L"m�n-�n�:U{���\+9��$�{"�3�1����	1�J��:��5-� ��Ak�u��ݠ�1�(��^�پ�إ��y�������Sg�Ǌ���힨1 �
V4��?���?=_��$ҧ���CSt�t}���Lf�<koB�����.)�y�;,zbM�ջ�� ����EMoʵ�� ��9B��R�ƹ=�+/�LM�I���;�ýCo���zx��rW�*�UU�M�o��S��&ׇK�Zy9�~nl�����oP#��:p�ɗ��"ZtL1�>�i�VM5�/��V��.6��l��>��~_ϥ�޲����O���Ty�ɣ.���YWS���_������Z���#Ɲm�ܻ�&��W�vq�u��4���E���m�߿�\Iv���\O;d���4y�O�pK�˧�vg@������̕��Ɣ��PHP^wo���ݕ����_�(�}\�f���1��}��$x��LM�׉M��B�6.�.��u��G26����~��]ԝ�����UrB*gG)z1���[�:����	;2�9B{�Q���f���\]�]t�싃��D_��o.���^�;���Fne���ഥHܲi�27���Z�/������^Y��W.m���̰��3*6�Gm���/9s	��%𻪪J^xw���HXj,�?�J�$�`����緟E�m��;�d٦^َ�zM?�N�i��C�
�p7ƶ\�d��0������'���UEƙ���!33�����Q��@��Jָ �HX�\�o��N�����]��3S��� ����t�2)��X7��X�1I�ï9ѯ��� -`��S6��}we1��}�<י���%`O/����g�t�ԥ�`F���%���`bzw���C����� V`bg���� ��6~܉a�\�(vc���%s�"1�}e���\��e��̞}�]k��ҩ�o,�Z7>���sV��	"m倖�RC�E1��N��/`��E��w��9����W��I�
�*(耹4��������W�*~�V~=��c�Sɾzcc` v�^!�}��v���X�r�^��>�7���nm�#�]h��Lr����*��%d+�k%�)3�7 rU�ꄀG�,++�}�+��(ᕼllդy�����w����{{{=���*�����l�,���~�
�:�2'##��ۼȥ�%̊�*��pB����wK�����J���x��4;�-�p�FFF��ж�0��g/m��`^kq8�#~,2>{����˚x��a�S��a���?�T|N�U�����	�����)P/5"=Ӊ�N-*�0���s�+,+���:�3�]bw5ހ�9o&��x*���H������8��V�1�"av���ݵ��y�1d+! !d
j�p�⽟�x:�;�²l�ۇ��ء��ξ�U4�}�#�G�sㅵQgP;}�� �b�Qp	d�d=u|yf��X�{�?�uJ�B��~.t;��.��J�4?�n�X�D�¿��s�vcfsk=F��d$bq��ׇ�=7պ^�\�N�(#���zΉ�aZ��9����&����r3%9YI��.Oꮥ �PO�uoT1�^4�i���}������xr�|�Fa*�O���h0�;o�ch��maq�-d��9?���� ��a`��U]X<:�7����Y@����Ϭ	�2�OG�;(�F�3=Hj��Ю� ���fϰD��sNL�~=䗄�o��� ��Û�}`�t|.yN:L�(��������'W	�.��#�Bt{�S+}m��p	rZRRR8{�(�m��.������N`�R�[z�ŲM�|L�-!	j�C�嬒_��8��2��T[Yİ���)`��X���lo��*�� �c�^3��<�3�����<�����4�ha�K��)��)��aG�p��ا�<g��y�O��W���W����Nhz��S.B��+��C%%E�nI�T��O�G/�>py@�]�7ǡ�	���_-���N�;s8<�����@<���/�X�x�˹�[qowD��3J//��{��/��5�p�w}]�Ч&���m~�W�t#B��5��.���޼���m�4�C��W�eX8�˃�x�	8#8�[������-��`smI���b�\�����Q׸ϖ�4�r��H�e6ڣ��]|��fff��]#� �GϜ��!�#�nzQX_��7!����M��[.��&_�Kr=ǝٍ�kf��y_�_=�r�N��8}�k*�T~�x~ E%���K�_1�m�[���~��3����N�_�4TC]力��݄�`��������]�˖Hy�D��Q�8>u.CaS����,�Bx�jÔ6����-���^��%.�FtE�v9^��d��EF�k����0M���5���h�Q	���ذ2��w/�:D�}||�Gm��xXYYq$R��_SG
�)������fn�N�:դ�Q��R�_L#)<��s}G�7F(�27+J��k��,a�>��r��������eu�3�v%�a�y6�0�������SP�h?;��듊�� �s� �gT�U@�L&��#������3ݎG߿�tCq>�Ǭ�X�;���ۧ���>ĕ(�YCX�`�c\���%���^b�3ݮ�ȷ�`6/��IU�{B�����6V�����,�Ȧ�7�4���Ry�N�>D$�c��+��_ob���\���ړ�U�~�G�}��A�j���]��W1�YY*��y���e=�ח)$�rM��oS�0+����XD�����
��*�UU�M�Wc�	�?j oY�~�^[0�H�,��`0-��x9	��e!��3�צ����7A��������G��Oѿ�����?u�N��r����>7-�PǷz:Z�H��~:O%`ii�j���gn��`49����������6ӂ��l��N¿r�L�ߗZ�Ս|���3��7:G9�vˊa�]��� ��i'���gC���Jr\=bO�����Oc_����}�~p�����=ZZ���o�Dq�tK'������R�FWx�Y���|���b�9��K���M=?'��%+�$��{-��x����ىyy�����0�?�,'��>}�NY�"��wR����G�"�.F��wn���S"Z�ъF��:#�{m�:*���l�++W;��c� �􎶩Z�t��<.6�\���Ӻ\��C>��0�[�+B�hj�[*�CD�A��Kl$���ݢ:�g���{?ľ�_n� �<�>��,| �Z�=�ʓl��*�����fA6?�1������?˨�g�^n��[]g	_8��	�ck�D?\h���b�N��H�n�o�E��L`n0T��8�@.�,^�Ϩ��g_��� �1������M�W��}��{ˎ�ʤOKI��9F���~�!)鷂q��o��atm_Փ�^�JX��9��ޞ��4n�);���C��atH�΅�PGSM�~�JUP*�ʂ �m�&�����J�g�����頿����̈́���Xw	.��,�W\�aa\�b�w��1�7K[�3U�)�`�I���(}���-m��c����y�{@aj�l��$�	��F��q� �쎭Ḯ��;#Q�cI������kqt�9u��q�o3���r�����YXN�����	��6�ܠM��Y�0���}oP�h���?��-�0�?����jR�v���_$*���z���t�B��w�;�����:��T����:�,	�t��n#n1�%�h�M��� �[�^�>���_���L�I>Q�-���q@�����ž�y�Z]Et�m���7:̞ЏNf��lL���� N��Vo����J�N�(��	����0%K�a�hb�]�e��3��o,�6z�_��j2�L�={.�\{��D��n���N�T�3f�6���u�-_®v�>g)=ڋ�C>+�:f��>G?#��C$�,���-^�$@�!JY���[
��T�ֵ�����������ľ�i3�z�zlWϙj�@�Z>X��DOԉUK |}��h_�lXԡ!{��V��O(נ�t�y���C?%�}��b�`����,X�s̓܍J�C�q�`<CQ��e�%)��k��f�B�UqaaF�HE��C4��HQ�J�5�[��Y70�֬";���f�)�*��+�f���;BnL_���}\a��^2sb0���U��x��=R��_�| �)x�R��U]��$�.�4ͱk1Z$�ҿ�[�*p��W��f9���S��އ���~����Z��9s��k>�/k+;e����?�'vr�o�ܾ<���m��=�ce�Ay �iI�Д�^���A�����Cǉ�����̢je6/��J׃D�|V�{oB�%�a��P������N��pp'mH	8�P��ߘmco_�$� ��y�[����"�dG�p�=��=�6�c��09�M�����=黖=if���"`/u ��H֛S���Οq��r���׹|z1 ����4����u������\�+�[���e�N�{1��)}nz\�Gc�t��z�+��Qv�N�fJ�7��я2�Gx+g3�7M�/� G%y��9R��]˫"3j[���6�c3{���6�^��Z��F�#�8H��'��	��؈�fcc��%��Qo�鸜�qz�$�`�~�E��H���*p�Yx�}Y�hv|�;Ş
����Ǚ��V�i�W�i;�D�{�fcR�/�g��_�g������ �����+�#Z�>6N�\ 级vv߾BZ{>�K��i��q���$�M���z�Y�� =�
DҜ�.�F/F��v�ո�.I�u2�g�m��J�`$�c�$������R�D~c�u��J�HM�7Z���*�O�|AF[,1;��G����o�!d2
��z��]R�)V�_�$��DS0��NS^���-�*.�%rAj��^�hD�K�VQ؏��n��#I�R�Ԉ��3�,ߓ3����-}"��p�L�ZB����F�d� �9P����+�jp_q�Q�\�⁌�3�<�8f%[Ք�s��ѩ1����e#�����%V����f/��X��DA%�}�ݴӈ5`�$=zZ_�ô^����G��U�����;������?����d�t z?+�6�N���M0�҅k
e�[�̎�3ZR��5���$n6����DZ����2�PҺ��=L~A�{/}bq�`"�+򭴌�Lm�0AI��^��7D���Pyv�!�*�X�	�*�8��2r�t�����������X�e�tb3��� a�hD�(�&Hk}Ϊ<�&Ew��F?38N�48&�	�K[��K*�n���H�uړ�/�<ch�4���������mXr�e�O���%����_.x�8���H��g�zW�C�`�����N\d���cZZK���/���<�#H�#aw�Ү��Y��·�I��0qG��i���߫��.�rj�[ZY��~s`�<�j�G(c��t�Kj|$�	�*
�61��'4�����3�O`��b�v/-U�T�L���=(&��O�cԡ�[Q��̍�L���*{�0��n&g�m�a��>/�i����w]���9uFn�_��s��M��7��@7"�=��>��u�3N�e_�(ߜ.���!%1d�|��K<<�fcތ>�$\���K�F2�݅ݜ�]��O���m�D��.�1���.�q��ư�
mGH��W.�Ow�RAA�?�/.�񷚮���)�l/���`^���]�90��~CJ*����b���xUV��rf��}���H�ժ���Մ��Z�]�~�M7֨�-Gb�/��Ca�JnJ{svp�r-��8�L���?o-�w\f��`fu�G�TN�^�7�´�~8
�B_�06�7rP�����l^+�j��;����r��o=��w�&��U��
3�-�XMRZB1���l�ԏY1i��[���[��j`\�ǥ=�9,�:���)��M�m�!ᰣ� 6/�{`�|�Kʱ�0y��y���g��g߄pO��c���]N.���6�[���rQ�J��D�P������+%���&��j��L[I����ѷ����{��*��T�������&x�;�8"�ê�T�'֥�O�S6��l��������eŶ���J�u�^mH���	�'F)S�͝�Ï�M��̤i�lx��'\`��Ú�1Kd�RN �:կ�OZ��;�CRC��ȳ�+�)F�w��Q�"rf&u���fn���#�?��o՘�Y���_)�ac������ڕ�����?������8��
�S���?Q]��ܖ������t�K����)�]�	�m0��%7�am�r�j?m�v�4Ek1cAl�S!1����;.la����gkqt$�2^�����Rb��/_!�bjH���X���O��W��]���Jn�anO�4��i�TT,���5=���]��;"�Ѧi/�v�N����"-H�EkK���Y��0���Ȏl�΢���.KP��J���f,��qGH���-~�6���A�0a��5֗Ǳ�eT��+��c�RK+�o6U�:�5vE��$�����b�#���)��<ԁ��\�[pwσ��da��_���82lO��L�_fH�%a� K��I�	�-9i�M胴����:��(e�U�IM�k>����s��X;��ťAW���G��-��E�")Fdjx�"����uD�U�t�b�ٓ<��o��F��
_�}�L�T�@���J�Y=}p0C����EA������ �<L�2�@jBǤ4���H��)B�M�G;���Vfh����}�}xp&_Ѩ�g�L��x0a����⾡��+��{ty����� ޒ�WBV-Jo�V�2�תw���/���3a�INxl.��p�m�M�om��vX{�	�0�uue��V�br���&�����o
8�_|�;�E����Y��"Q] ��]u]L���|��-ER��7][{NݧD�����t�g�U:�ⱙ���z}�F@����t�}rb�8��-Iu0��|�+=ZH����J�)�+q(;LE�|��o�[&�)f�)�Y5���y� V��Y���Oރy�h'늠�F����*���^�sEN9kk�2߳6N���M껫(���F/��J������7�T:T�8��C\?}J�m�ѵ�cfsdua�'Mؙ磣<�HQq.\�(����M��}�X��V�����p�KQ���՛�ω���4P�Hyy'ʬ�$�;<�o_����2������Ԛ��C���M�"�./keBR�x4��ʬ�3b�	t$��"�W��~�w{^ �尼�5�v[d�HEfDף6� V䯞l�1aK[�����8��k�n�@�����o��6�\�m�J+[�W�LJ��I����$);��v���B�v�@�ua�U2ϟX�Bd�{���o�D$���#uH������+niEY���wYvH��4+##�
���wtÒS�!�ДY��[rG~�����W�ڙcɂ=1);,�7��>=9ӝd&��Р���N�����2��O��2{����}���T���C���������M� �L>>�=�}���i�1���V�U� R��	����F-0K]���������^Af��yʱ��ݳEMF�A�
9��oo�Ѱ/�#u��>����H���O4�g]{<���)kd̈́�s�P���*���K�d����|�D��" �i8ʏ�"4�okh4�zK�w�1�ڄ��hzX�!�_>Mg~C�B'0_�� �%s�-I�"�t������L�r�<�z��,eS�/��fJ�M�� �����,�g�	ߜX-��ٴ?)��˵��|�P�H��[�ߡ�B��6�rU�v�p�<���B�V��;����d�M���l�K{C�`�t���X
p����n���[n�e>��Wl"�������̻Q�1Y���e5�ϱa�]��鿽��jk@Ƹu�e��g�s$DL}T��,���<2𨢬ȉ��F��b�s�J⺚4����A��9|o����Rz`�$��n��s�б]�d���NY8FKW��s5�����s� �D)��=����zh]��o9�N������	���nj�g=�n�Z�G+��?&���ii78�D	��7T/<�_X�Ps��_��褃�S��J�.0����P;y)'�K\���s"���K��dd n#9��G�v��[֒�'�#����J�����`@���c�	pF��}WWL�l᳣��g6�3�i�h#���G�#/��J��M�b�+��[�����}ۺ���I�b�Zb���~,c�u�K	��T�eh��)�Õ�sK���w��?��+�w����:��$��h䝳�����%g�z���l�kY��oK���R�e�'֘t%�F��-Зn���������F+��s_�D5E���b��q5�8�5�+��5D t��1r�}Y
�247Z��)���x+fI�v�&�~ �<x�:�]ʩ����(H!��Y&]Q	|1P�9V�A����l�}X�`��>6ذ��"��\f?��=k~M�W��>���J���}�ߐ�����Q�ʫ��L"�\H�=�^"��X�`��w
��Pzo[#�T��	G��z�������3yy�i��.nS���·�Q{���Da)(ss��r&!b�	��e:��ñŭR����K���}P�1QzsT�D*���q�t��q����9�1�R8����|01��=kp�=��������\�-8u�� .��j��s�����'
�ߨ��9�t�=�,���9��ϓ��#���,B�/𮩌�.�/��P�p��vI��X�<t����ȘF�� ��J��:a���OGV�������'��b:NG�jw
�u�#���hEX瑬�ӝ蹭56���r�3~������a��1��ޜU>%'cg���<�޲��S��)��.�>h+�Ye>;L�ǗRQ�4��k,H9�� >�zN�sC��!�.>r�)��f"\y�Q���NK���RT[�yi����3��ŷg��q´������1�oh
�?�XJꅰ���#��y�]�w;��M����;�)|ȇځ���z�&D�u�b���,��r��BxG�������ߴ$G㳷�x�(#(rm���y�+;�i�	\�X��^��*I7ZoWu*�3
r<)C�=S}�� ��ےJL�M���=�d*������/+�|�X��i��S/��x�=�V&� �s�o�ao�F�Ԟig�l`	���{E�>�ઉ �ں��%��%}��lNO��mN{k^<B_� ||x��$�L|h���/eUBh�5�?~�J69�I�B0q�C.B����Z��"}n��ֽ�X;p/�@�+��<_qFD�;�����)󱮅��f�z�{1�7��x�"q����Ti�Ǜ�+�!�Kz����B�2�Ů�A�a-���ES��~ku���u�+�F'���YYdg�G*Dn�o7���7��E�z��rS=T��nP<���B���\-��A)qZ�'YZg�㭎U�Fofݰ�9nל`F}B��2�ԛ�@�3�m��M��N[U�z1�\��7�D~�jQtB78�=�3#:TG���r7���'��ѱ~��Θ];�"`�7���h+�����	t
���A�����]���Ba
*1�<Ǳ|ݶTrD����I�3�J.���
� 0(����C#����~斞V���f�5�H��	Z.^@�~On�O��:L���%� ՞��7�=:.�i���2��� rv��H��3��)57�]�&!u^,S���Qxc�]Z�I�TL�oKw��h:��LV�y��Yo���B�a��t�=��6�nʆk��Зl&m���S6�Lw���C-�����H����۫\�(��H�A�uy��ƒ ~Dv�|>�ҤxN����f���2#�3#�@�L퀗�C��������9N�r�q<��F�Ri��m��Lh�IF�{g�@�都�9�����~�<��tu��l~�	��̨E���G�����,�S�pGX,�+b�c\`fP2� ne����J%Q	J���)�+�P�'��dHx�>�:��#�̰2q Q��:,�>F�=��n�<Z᧷t��j�z�<�Z =o�8�3�J���*�a�;��,bH��v~v6֎?%J���X酗�Z��W6�j�G0j�03-��7�n�!�9DtiR��e��*#�U�;rƾ/�o9�$NU�� �z̚�ëE�9O)$�~mg;����QWmѿ[�\)�\ɀ��ܳ!8:�"��5���8(#zL-V(���X$���p�dS��]/7��6MU墊l������8?����b0qy���Q.� �|�?��L����aX?�( �S���l¨�fX�f�a�Q�͍=~Z�U�+�f̀c
\�X᜛�#�ڭ���*���K��u�ʹ�+k�/iC�#&���Cmm�#��^w?P���S�����GQh`G��vަr��U֖���� ��e�ɫ��a:� ֠}Yo1��RM@[;'1߳-�^3�B�;,���Kt��a�R�̨$9�inZ���k�suo���"1랴��L��t��:��ph��nR��}�� ���m_%����6]�d���]V��G�2D�\�%"����)S�禤8phY�������q�p���:��ݡ�P��t*��:��B���Q���]S�@*dx���{������'����O�C���"�h������'(��hѹ������uv	��'b]��9�p�F5ɘ��^)έqg�;c�T�{)��� ��e�wpZWr�O�j��%w���P+�_�&^V]M�'�(����\9`�3�v�<��ϔ�R�?��O�a��gj��uf|��N;بkP�h5��7�r���,h�1�pE�B�܂a�OpR��@�s�_k���TY�$dz�`�	hn
aI5���J�2F�]_������#������%��Pl��]��n/�>�3Y����ؘ1-1��^S��B誩�aS�g*�G��{��vP��HeoHY���b� ]�WC����_����:�(_c�A��_ՌL����NKK&5�Љ��ArO�W����ʛ�'ޫ��7��S�i�ԟL�I�VL��%���'�#utb�qnQ~Q���j������ǵ���x�Z���'P��Zm�]ϰqC�r�=}Q*����[z� ��iT�A	M�ǰ%)��h�B'��j9�<C�?>�!+C<FP�\��.�X�~+�l�4�ܠ<]�}����^�ϔj,��]yN�t}��՛�wf�aA��8��L���O|P���:� �� J�����T�P�aҋ�f�7��RԍT�{w��'o�H\%���B�LDU���6:����MB�D=q����T!|�2�o�$|��w
���zȳ;�n�UrD���q� ~��`(�@'���p����;x�?��ߤ"�OUZ!���F�InQ�g �[!$��hO�}��lŅe���Y7q�ߍ%|N�u�ҥ�i�t��nx��?�h����o��6%+2K�A�p�<oH5JW��zG(�Xz�#�u���J��z�vM�s��oN3�y�Z\�z�s�+���X���g\b���5��j������5�I��{�ҿ��k+��e��FaNp�ً�j��'����z�jN��f�Z��JZD����l�8�n��5�i����%qvD���c5�HK���URS�a#M����d��̟`��J�klJ'�p�8�F��.@���M>�&�Up`�+�\�rG�[�H̳9X|P Dq�G���bƢ�����d��F�Tf���Y����>�yl�I����ŬrlR�_����P����~#1ۋ�w8=�'v��Rv�ZǨ��!y>C�G�<mL���U��������Tz1�gw)�/��P�����B�0��<�k�%¤�
�W@�A�!��,ƍ�?x��v�䋇C��Ya\_ZJZfk�}W���X��`VH�]mFrS>�VeW�DG1��[�Ou�a107�� *�'%��e}��I�G1��#?&�؝�_Өm~��T��uwOD,PQ篛�w	��A���
��jp�¦>Q	�uY�0��B9�dQ�)-+�3�&��H2�q��&��մ7$l��ٵ��@��}ǖ$cJA$C��>��Ӧv� 	�t��ſ8h�u,u���.���.�\�$��K���b;{ЈI	� Ժ���5�Z�sq��Z'��,3y,p����]A��p�� 2e�$O�<\Tɻ8V̮9�-��i�k $��/�p�~I-���F��ύ���.Abh��PP&��b���5����\v�m���X��ī���M�h���':��v0}�]\ޅ��T�'ǧv�J4���(���?Vf��=HG�k7�#I��jm�w�k:/�23I�uqV�R���m�>�18�e6B�}�s���D��������|?�Cρ��q�p�#}�UU��a�3�,{ș,V�b+B�v 0>1�̫Q"=�ֱ
�����4�:bU.T��Ǆ*B��0>��Rw�A.�PC�ڪIօ�u&�bw*Ѯ;L�M<d��-���G�;��"ݲt����n9�:q�Zh�a�<�ҩ��<v`�d\�{r"�=mK<��ݹ��=+��9I^�}��t��g�2J���9���,��;Y�Q��=�7ϢZ�̓v���W7,�Ӵ3������ E@��j{(��Nr8g4��x����|�[h���?��z����A�9��c(u��O��>̼�����d�]���,\��=��~�\��O�ޑ<	H	���+���t7,�a��2�+�zo�f�5��-6�ӑ̩�qM���Kֳ\Ҵb���+�M�r� eB���4,軻��x6ܺ�W�� �_Z�7n4�>D�{l��A��T�@��H�V9���Jur��q�	b�P2:��E �l���BBR[Cw�I-�i�&/2ٓ`�g���ej+P���^ k,��q�FSQ�ML�Lk�j��&l�l�BM�*@����Q�y�S��2#wNK��)jt������u� �����w����PHup���f�����l��3��[L<� ��w9B#A���5�Qt�C9�w7���V�e+u&O�l�,���	c�Y�A���s�q~�����*\�g�6�n�<���g�y��W�Bߎ���I` I k���~㫯�z&�8�rR"��"��.[e-7᪖�l?g�v�o�t4��N�#��{���9�F���R�NYW�5/��ǵn[�`�d&+|РAV!�oeee���1�T��n�;�b�	���`g�8F6��p���XR@B(�� �-�@�߉\��v��;b����B�q �v4L�L���w��δD?s�i�\e��6 7���vW�4 �d�'�>�LBzWqFz���X��h��ay�_@���� �Rα���q� �6��k-��LyS�i@�� �1��� q�7���/�;�2�P<�I�C\<��8L�)��
��iiS+W��|i���Q^6�N��[���;�l��yփSZZZy�wN?~|�@znv�x��|���{�/@ny�%�\�8,�9=.�Wr�	��TQͩ}`3��F�V8x�c	��e�`'�B�E�A����9(��������w1-^����[�F��(
<�������t~C�� H;�\�r�F�cEF,��>3#ۆh�s����l*<�壋!�o״�L>@|�ܓL\� ��Gь�x#�=�mn�6�%������LT�&cj>4q�Z�w��I��A�f���ĳ ۑ�J7
�t���":��` �Yn��MnlyY��z��[�s �֡<kI]�)�m@��od�'���x��.H����~�[= CB�;Y������l�w�CQ@FڴR�UUU��g͚K�#�Y�<P������+R��3}�B�M� �q�� o	x����wOF���c����6�7�%KK9.\ZX��%�Ȱ�hpن��8i^�i�-Mݹ�.����n��>]2��y@�`��s���V,�i��0*�Ҏ�c�$,]� �6���,፥D�2�>�Ț��;%�qy3o9į63!8�Y�����B�`�����C:��fw��Bm̗5�m��zM��x*Z�&����0=���}{W�c/��"��ކ���ZY����Qŭ%�`��/4�gm���a��n�~-����@.@4�з"��j�5���`��_G��]mrC�f��B�`�h3��Ȥ3��4:����ߋ�+��Ϛ�(D��D',qzL@vZ�~r�Yek��`?Vnk���?�$ ��q�$�ʃJ�-D��N�[�{F@g�S�θ~zfl�<���
�\�,S�4A�uF�������˗;u�qLʘE�O�GĒ(9G�dP! I���lͽ��;���(<��c�[ĳ�w���ړ��%p�}�w��]{[G2-ovEs:���`#(�Ũ:���gNЦ�Z��|��m\�@�/an9�@0b�pk��joFL��[����bv�v
� ֌�2F�+�#\i��c���1�;@B��>���;�+��֭��W��Y�Rѯ �q6a��)^�뎃��c�"��a�Pb8�v?Ҭ�� �:�� ��S0I����[h�8�t�;�\RM��H�� ൢ�i=�,
l�ë�ĵo6�p�O�6f��
͢���\�ԅg�a�_yG�J������S�B�U��{p=]$�!,�E�l�&�}]U�����Ѓ� ��>�庐��8���P��8{ͼߡd��A���V��w��7���ޘ�D�q��>|�W2����7 �a_zG؈'j��r�h�"��k�E*B;�������ԡ�P���Ќ6���#�.]����/�3�Gd惌�����L��fE��J.Y��s�,�O����'��@UU5	w�u��{��m�V`A��3�)���hN�p�ָ�2g�ַܦ�צ��&%N�P��+��e->k塠,6���0f��	"�����&���p�8Z̹�*�������⭴q}Y�ֽ����Cl#8:1\;����`I��"p9���I+J����|��N��Z��� �*+ViG�u��9f��cM~�L��Q����h���R�f?\��M�&��lB-�~�Rf��%fJn�9`�X3�����AJ/ ��2��̔�[��|�!��a�w�5)���[o�"T�{%�h%p�7�K��w������(��V1<T��T�����
�_
C���p웞��m� ��ߊ,�9�3�A�2�kŊ�E�����ݺ�my^GA��ƌcF�u�O�����1��!���a~�C��h<KIP��anĿ�A,<�z����|�x.ұ�d��^�wq�y�܏y�Y=}�A���}з�y;z�x饗����~WQQ1��I.�(�I눋���ց�h'�Y�>�XV?��X�p���ۊoNmwZ�\�U�� .��#�{�U�:�Z��}{�	�<���yy�����?��2���p-ww9YKn[�#6�m����x��8Mf2�(%�c"k��yK3� i����Y'���n{�1ӎ1�E�L\r>���� wm]��.pȴ���Mg�j�VfF%w��F�y㆚�4x �\g7�� G�5ޅ��`�Y%�
_t��������`b����"�@R[�������p�[gYY�� ,�9J��^�ŋ�oX�֩jgr@H��\��(Zݔ�' �Ly��1��(jjMKPokk�s���2gYߒ��ʘ���V�j�s,��y/�t�{R�򫯹zzAa�G��]�v.�����bΎ�2!��͛7σE�.��C�m�c:��	�I�[o�uhqq�K����Q yVBYA-8�߅�� ��b���Rt"|�o�4�x��i��$0�%p��w^���_	�t�
�XK�ø9no���.���Z��nۍ��ߌo��r���C0C�˜<��Dn�Nk�/-�����	r,v��\$�E��7,71�	 ���g�}ӦM�	.���!��k��f�eq;9�
T5c?��`��t�6g� �3���inw#�ߍt�[��ZZt�H���sMְ�d1�&�FO�z�m̘�����r�l41�%��j��3�LZ��(HD��(^�}i�+��3t�Đ� 0oA�?,�F��q����ĿR�Ïk�AU8�G��2l��~;�0��e��I��U��<|B�$������+w*�9� �/eOYp�P.̑F�zu��Y0�[�/��F���Q,���#F�0U5�棏>��潴�w����(���0HQQQ�����IG}�#�Qø��S�����|2E�`̩ �7�]��aÆ}�y��z�ꡰ�W���K�q�˖-+�<l�=����\�zȣ
J�Z�{%���w��5{��=��˓�N� ��<��?~�Řq�ܦ��҉j��K���ú��~&З�]}�eY����b&\� �u�ז�ޜjnr�v���{�u�}��Ph5�L=���{]`�(T6��nzE@<��,lV���3�q	�RLl�9����k\t�`NҲbл`˯v�d��3�0��: �c�e�&0�`�77���l���^[e:�^�E���VS�`�lf�D>r�C �hia�Z7e�`2Zp�`������&�y,�����Y;��5��]\�@.��%�l͊O,�1�ٍma��9���~�I l�$�I����~�<�F-�S�Ԣ���[OO8<B�*���QA��H�e��z��E 0��b4j�Cŀ�`Y�]�������Y3�������ȩp��@#��L�آA���%m�ر~��ǯ�{�?��<����o����J��r��4i���6��� ���]E��u�}g]��;K��y<	lG	\|�wz���O"��-�d�ÝR���4��rv�r��3.N;��k�)��X������� /FA6U�Bύ�� ݉�:�l���sQ�Cl.[뛬�X 9 77q֬�X��eG����,�����UP�@�uL�/ƶ��
w��o�^��qϓ�����w~I� ��q7��m�O4C�F籸�X�m#�?x��w�7PDe�I���h3� ���ֵ�t.+�y�&�_e�֚�f��@�r�ʰ�Ŝp����k���'-����y��Enx�Y_]iւ�W���Q)�G�9z�����A��b�K�9鼿=V����En���V"}��,O���9�nN�8��;�q�ȅ��Vz2�,<b]9<%$$�5�xϳ�d����y�2#��޹� b⸩�)���3V�s�R�p}�s.��lfFdee���Ǉ-�gђ����C=��s���}�_�r�P0%B񸮘�ںK[���B~�& t��ިW68y��>��?x�(�C˺߽��kp��gn �k{����c��y��$��%�|��a7�tӭ���!+ƍmmt,Ќ�:.vX��W��1t��ש�F g��0���<#��q���ئ���H���	v���<X�y\Zx��,�H��\���w$K�x<�m)
Ы�(��I$ޑ|&���n�sG�P�Kx�=���i��c:��p6U����
�m��e-s�{��Mn&x���ʴ��9����2��:���p���oG�ض��Ymf��i�N5c� �u&�plx�ߎ��.�aI_��P�~��_�@���5�IE�)i@s�lE|�&{xQ@.������0{b��
x��5�# ���� �1u,�!�!�v{3z� ���P�!(5� �r!O��g�.((B���WX�js�(՚n��t���O���z�S����^ıQ��RQh�n�ǵ���R�7v����&׉�ic�h�0��Q�s�>ˆ-_�?x���p��0>�i?��'���DM�0����xCVNnegWp8��a��U�lޔ�����toX�Mp��Z�BZ�s��}	Z�>�/�n'/I��<	x�<�瞿~��G��6C����"6ш��9 F��#&�8��݀i��߈�kl���iAQPyUZ�Mw�������s�'����'X�o�9c�Xl-Z�'�;�-������6�c�;�eѽ��Ў�}6n.�C#Bd���{{x�nc�zg�u�w��f�&6� @g�
�U���} z[����?����h�6��$!%��7\��MS� ^�`v�k�5^��d:���Fgd�����2b����):�܂�ҡC���t�O���޻�.@���@�����{)��oYG�|Y�L��=�A�����|R����G8<>-lZ���u���9��(�{�n��P�V�qpU?�����s��ܜ;lɚ������~���6o��QYQ�n���P�E��pTG�9����s~H��|�LK����z�?ڸ�����ڴ��Ƹ9�g�OO9��'�Uxc[�=��,�xW�1y�'�����E��{�upƫ�*E.�N:�CrS��nXr�tk�e�)�g�9�WZ��yv�炬*_���0*�MP�
,;�0�`>�ST�k4� ��s.ܬ0F���Z	s��s�����X�$ө��n$\%�9}=չh[Kܶxu��<i]�3�
�6 mr�cL��9f���7	��\Zڐ��{�i����5�"�2Q�`5�7��5��c�S�Pj�	�Pc���88� ���ՓA8�Bӕ��TUmb�3���+~>��c��<�z⤉��ݿ�/��k���g���W_ۇrq*���e�$n�9y�YY�VA��Y��~�J��c�p��)�[��߈�r�T���e�X<�5[JI���~&Lp���t) N��x��c�z�7N��~��d����^�də��9��3G��Y<�8NJ��o���c5���TU���`�}������_��h������?�S��Ɠ�N� ,�8��nX���C�7��-�b�8MU�x��Nw�,sY���.S�ޕ�ҭH����f+˅c�R�H��s�U셋�j}�;������ N0wwBs3�Y�TֹW��+ے���ؒ�����cK�r�
R���h�:�?ۤ 2���f�����1�L�,8S��m*k�M+R��p-�!`�M*���Ӄ�	Ef�X�TH#G��Ӎ�P6mTQ�Ղ{5b�5�����㟞}���y�q�ѩR�isꞏ��9���w�}��y;Vs�I�N�c.8?�����0ġ�*���������[%�aÃ��<�і� k��YY�k��f{�;y�Jw�}imA`8�s���Jޒ�_�����C��Y���'.����kX�fm��Y�v�Ĳ���G0��L�\�"�9�g��_� ���l@XaҸQ�\~ż�&��E��@�����x���K ���+���)�\]]kL��m�/X���*�[��lV���p-|�<� �:"q�����W9r.�*שEZ�B��mƫ� P	�5N�z�\�	L]E����׻���B��y�ybR�m�I K�z#l}s'VN��픰�U�w��V#b��@�1�x3��lO7�Y�ltכ͛ZMM������Yї<���LΪ7�.o&e�:MZF
,r�3`a�B7���XcYj�����#�yҷ/�l��Y�>�^�juʊO>�L��!������Ȅ n^W��Nv�Cx���aIua� ���~{�U� ����QFR~�'�
�P	�1c慣�a.Z`g�9�ͦ.*$O
�]
��-�G4���Z�d��;�oI���=;;�������`|s ��K�xN1�h;��I���������"����	�i�7��G�����ޛ��;���������eoO��o�uӦ�s��U��Jy���v�J��l�/0�8]p��j��(H�pcզe��Ŕ�0���"Y�6�m1ñu�U,�$��}m�i��X�-M�'#>�]�X{��a�R�Y���)��MޢR"w=߹xt�d��@�⠹��k��� ܴt3���`���Ջ��ZX�]]�"S���Ռu��IJ�5�9������Ԃ�\�����0���9�s͌b0�Q�%6�t��.�n�u`�Ԇ5BWb��h	ZWߞ9r��=��iG|v����^܋ �|�'�6���n�o��o	YŸK�2s���f@���� �ܺ���P�fH|T1~HO�r��4h�m �n�:0���q���Rg��6� �L�8�:��է�^W[g�����U,k��k1c296�`�n6�h�"�c�%�TPQ'�	�/3X_�v�+�Q�t<(ˋ�@F��@
�c������C5��ւ{M���/�^Vv���n��7ջ��[�=���t�Ý:��X����թh�:���.7���ח�
^)�nXű	�)h�����0��E����nk<A�V-rZY�Z|�7o�EbT�L ���]Fw� �E��7�qzx,y!�O!ࡘ�-a˖����T;�)�)hTF:Y�.1�L]t�1�p�4E�|���:�#ݯVyWS�In�dffu�ç�	�~��0ac6G���}�}h���c] ���S��Y5j���{�M��Tnˬ��O
~��{!��Q��u��ͮ���I��Z'������{HM�q��ȅL;n�u������w����+�*{����6��� ��ޛ�=&Y�Z��x�<)}qy�a{_��j~I�SiX��9Ǚ�H뛛�GO�=,���܏m]5W�<�`� 5���>}�[���0eʔ�1GQAh��<@���w������=��� ����s��\�,�H,tZ��6INU��\P���|u)
\P�z� �0^�����j�Dl�/4� ��[�)����ZP�2#�:�4���@�M�%^?O��ǡ�@����r�,�w�[�������+ !�B���%�XK�)��{��&!{�����ִ��T�6!�E]�Qw��L	�7'�k�����`=,:T׌�i6] ��Wnѭ��ެ��1S��w�e?�0{�H���؞���@�:��Px� |
�F�Kn6̀p�\ɒ����j����S;�9r�5ot�x���>n�8+s���v���ga�-�,O�6�)��>}�LS\4�*xTJJ6[K܂/�%���@��V����	̜C$�q~2���@Q�cz��9���'��=O<�q��z���"����˞���{�]��i���/���Q��b�أ�h��K�����[�U����n�i �s�bK�U��UJߝ�' ��.�J�JA4c��E	�l�9z�(�7����U�V�	�	9�[�"fh�C��{>��AŃ��@5���o�HFz'��CH?�B�u����B1�/g�p_�;�D3j��&:%���)���
/Z�M�I�Tfr[י�G��#&�UkHZ� !� �4.��02n���k� l��X�C�Խ����o�p���ބ��)����5��LxZ�a�QNv \����`n�vsxo�B�r$�����ĵpu7݇(xD��M�%�u�{-�Ӷ���m��>�c��eja%��=h�3u�^��/���ڵli[t�W��W���-�9�q�ĝ�l����0o�)�*_�qr���ͼy���k�iON�6m����X��K�y�������	�������|���V�d���b1�^��q���.�ҟ�.�F�9���^X,�.�\��ƅ�~��v�|d;)H8bƎ[>��H�.������Gpwb�1Mʆd̸�̹(3���ػw���~�fu��^�8���߸�NE��h0�&o�L3y�saI�D���3��hlR�cjQ��4l6	��ʹ�nsּ�fdB,r� �{>�4��9]�(Ԓ�km½�D)֍�SG�x�ċ��f��k�6g�}��/.Y�����
���G�؎<3w��[;x���y���MJ�,g���օU��9�;�񾒫F��o3�B`܍�6�x��"#=��C~����j������w��q?������
��l�>���ps��� g�I�t+�6��� l�����I'����	�Z�E������{O_@`����x�a-��H��§�4��H�uWc�;[�Rה^ƅ��(�r2��OFo�ܹ�ˢ�� b�HE�5,;��J͂+��*ŷc�ߴi�z�Y��w:�/�9-^���7�%�3�{3��q�&!��.�/�q#V�]�n�΃�YJ�2��dFM=ڄ�
����^�q��y#�䡆frL�9~R��14�$Fw�9��m���3����6�U�rVZWk�s�?��+'�b�1_y�}�7mܘ��[K�}����WVN��l���)oy(\�Wt7���)�E ��t�©�Hل�����d4C^d���A�@��T�c����B|��q�W_�T�����O�S^حd�ڔ6�p���q�pޒ�N@�&�*����%�K�ёGq�����ĉ6}�Gr��������;K���ߜ�2��!9���mOQb5�V��ÜE�a����$��-_���IIW[�P�@[��v;ӱѳܺ�Yl�)�j�vbc�Věa�[k�g�����a#F�4Y�YvQ�B����KJ7��1n֍���}��mS���X��s\�o�Z�d�+͏k#�\G/뻳�-7Zr #�CɈar0d��-4S���I�	{�-�R��0��&Ђ����L~W�9ez��?
I�D%���䰳�:�cc����jB���k��fą�����������x�׷j��̕��,���|��{���T�ohjJoA���s0���܎�/���V�MƳ��k;�me��?}���]����6*��H�k';޺��H�@�ڰbE�txN�9C�	-��A��b�VX�d��;�����
#�@\�w�O2"hs^�'2dHf/��������P>׹GF�S�9����N�l?~�#�8����_PR�	�%�>}�|I�]�'��)�G��Q;�z�����q�cC�T��B��J�l�݄�Tv-��v����1��ʭ�zxl��]�Y�r��� ��u1�E�+**� L6;C;�:� WbALV����]�N%3�4�!�J��M���vt�b����?��g�u�z�EI7������B	f�~�����_�`��Ae%��T;ygc�	V�4�涛����ȁ�\�Vh/�ȶ1HN����jAtۀ�n�Q��+�|�	��<ˊ.[���_~�x��x�5Ëº����X8�kk��#�;��M ��S'��Z�9�V��L�@��S���TN)p��0��sB�T�w������#9p��ra�w*t;�����+W������5�yY���s-\�f�w��K�>�ȧv��ұ=@Hw�˗B��z��?����M�u������Z�$;�m�I�x8���b�֊E/mnZ�IP#��=I@�b�z�$8�x��ȝ�*Xm����i9�XLm��̰`KW,�m�{����I^-�Z|�e��ī, 	���yn�[��ң���n��9�z/Z����B;Үn��ʙh&���;Ϻ��l��%FKJM7r���5fD�z�x��̃U��Tk,v�������F�s?5�6���(����~�-�=��e�V����s��=�2J��\�		3����y�.���Bߑ�?�]�8Z������m#X�1>+g���'�*�K�bs�m��x`�R��>dm���I��B�|�E�9�q1�a��fJ�r�d�s�����A�rH�"�)�Bqx)�v)rǃ#��	'�p����������z��$�_$���7�x�[M�-���"�9nQ�N� ��^�L��w��u��)R5B!+mH�h��:V4�j ��/"�MU�K��~�sZlt��H˷*o�Ra��;&,P����`��� s�y>*)���)�
g��U��s?>@�7:`Zq�æ/6S�f��
`�'�z�|7��U� U��6��)u�[7��&%�y\ZSM��!�n���,�C����2�@2l��5u�u�.y����Y��n_}MM�-"�0�QLt�ض%���L�g�/�C�۶�"�J U%A���7x��Z�|罓+ܶ�e�9���-�y����j��Om,���{)x"F�A��a~�E���T�8�:��k#y�uY���]�Ga$����-��K.���Yv��<@�#o�wQQ�]w��<��w�s��H.pr{r�akLZ��6R�8�Bn�I@��m� �c4���d�+-M�w��V�S6Uy�vF,> ���t�ع���lkx� 8�N�<s-���tɒD'�B�%X]�JD1��L��b�v���,�ޘ\3f�b3l�I&%=q�ӌc��W�vx97�6��5昑Qf�p�;4�T�M�֥]-5����,���%��Z{Vי*���&'�:��ށf����30�K$&9),�̷�*�@ ���ۅ�X�@J���*�J�I��	��)��6�A����(�@W�/+���Ђ�`�2 "����q��ʅw{qx�=^����'�By�l����^T��n��(�EuT(@π��I�X��������N;���S�n�����_Dz�o=	l�`��_����e} ;^��Mxr�,�@KkX�i�E�ɸrQ�s���c���gYe\ܵ��o�Щ4hq�E�����d�sQDC��߷y�����wt��B����U��S1P,��]�@��+~nY� sM�q	�TnP��tG��?l��~�yƗ:
��)fMX�Q��PZk�Mlc�9tXZ�v�qY�CKN������1X�;�g���H�B���6S�㗡t��'&ކb8VAB؁�ud���4b�n�oh��i�=+�[<*jl�R�P)�]5����Y���a�.)s�i�+�z�����xX �t��ߜ��!_�g����O���T��oz50��q��h����ڵ�"�*w���˭�c�s)R�Ҩ3_Õ��̙�~���E}���"nã=�v� }��o@{��/_^7��/���[.�)ɩx�YEnB.8���1�\�b��G;Y��
\�i�E�K\��*w]�N.j�-g�n��Y������aAe�:����?4�ne�jZ�E�sG���b�\Hy~.�J��5���k��M���-r�.�q'u��W'�m��S��)'�X��1��[K�L3����7�hm����E���(1�mO!C��{�l�JJ�V�U�հ�75����j�&�F=,r��Yc�y��:X����G�3>1���~	D5W���o�Z�V��x��í 3=�O^�l	�j������ǹ@w;-a~oCT��ܼV"Y����Jh\��v����ޅf8�r�UW����v��d'�%^c!<LT�ȵ�w,+K��l���XRtt?8v:���TU�c�t�Q����:�NF��x�'�������{º���p�k�&	<��?�C�`X̳�&��� V�'�S��	'��zV����������n�8V�D��GV�Hb]a뙟;nx��@=q���p�
&��h	F���~r���
7����Z칹9N�IX����my� �0���ƿ��j��;G2�9�{U�!�!F�8��s�b��nN 7��'o�jB�x��e&�s�>~((ɦ�;�Ҥ�X�L{r7���I��11f^a,H��`���v4 (m\qJ4a�5����˫V�� t?�����1�F'�:�[�C'Т7+�1��5�8V'�<���r����}ܩ[����mL٫����&8Q��M�R�t���� �c���u��NPV���n���s.�3�1ʝO�����������������Lɿ2���)bc� �	�Q�˶��Ʉ���`�Q@S"[3����˖F����X�Md�r��_�uH��Sikog�Z�{±��G�ٳg>p�y�]5m����%o�����;X���w�^~��7�xӵh@1x���V\�}�����eg�q�m��~�ED>���ʘ�\�ӧQ{d.Z\XUU�����ֈ��aEp?[ ��>���/'yH�U��V�M����$1E��W��:A��6Ps܂���H~��v��;�S�)}��q�������K�>��8J$j[�:�MC 뮞��k���+6s���d��n2Ps�n�Z4U�TUi���m(7��	c���L��eμ��t�5�R���~$�f�uJM���uk͒��M,v?{���MЈ�@\�ն��P6�`-W/��'�-[}/9Yk'Q���k@ T}~�ʞ��g�lG�Q�j:����u�y.YӼ'<�M�/U�S(D^ṿG����9�8FՕ'r\|�ژ)��=� � 3��S58�%�-�r���=�=3�sȆ�S�Td[O�ѡj"�{(;����� �x>�=p+7�N^Y�|�c�G"�����ZB�g���.��-���� } �o;D7�x�EO=��|q��咣��`n ҿL*�2d�s ��v�������g�=�l�5u#�3�ӂH�Ղb[L�%w(-���\���z���j\��rW.����	t<��HӵI a̜[YY�u���5�G@p�(,�|a|���<���c�# ;�'�1SZ���bc㠸 �Ob,&WM%W��ef��Jl�H��>֍��/����KMQ{�9zl�9ķ!9Ѧ��ڄ���EHk;!=�D��X0/G��'�X��G���:�D� ������^���6���4q��	"����X�<�������x��y�w��	~����!Y�<V"
����-�c��`8��@��=��{-�ق������C�)��,=��k��p��HY�|�qUj��Le���p�V>Cuίd �X����6��,t[8-R��><nfv��l4*�\Pৼ-Z,�r��E� �-t�^ʊ���9GH�龜�|��`��l���;�����xw$�y��yVl�7^�<�ȱ���o��a������ɲn���c	>pr1�����S�Ǣ��{���/�m7m����3 ��X�S,��:�dfbĪ��z�����AN��ܬ���2���<1H�/����6���T@�}�p�LXQ��9..����`�˵��on�&*r�r�
��XbXۅ��S �lw Ӛ1nZ��%��0S�;��?�h&�Մ>�d�7����mfj�9mB�L)B�ׄ���rT���֔��PS�i��B��/�ؼZ�Jv��cl;�r��Vܵ�w.�n+RӚs��E����R�X�n��o�G q��+�͝7M�Ku����$w~f[�☲�[N�[�mA����,����0i������ץ��6fdf61�l?}>|��J�|���yI@��1��&�SU�8&��b�BH�����E���8��1�s�P�� "]J*ȏ�wP�n�Y�D�Eſ\?HqkV�㉃�C5t��yܛ�Gjpd=qγ"�]�3+2m҉��]kKW~�쳮>�so�t)�=<@8���v� ,�'�As,�\`�N�;@�@�m����"��p���|�p�;�������]|������}�DSA:��`-�0�)�,f�+��Um�Q.�-�fe�D*�)UI�b���sk�c��~>��:���a�|r����"�:g�"PQ!b�.����]�=k�AΪo��	�t�G[%*�,��U&6g�Ʌ��[o6���Ғ��5���Rsp���=ʌ��������mt h��M 6�ʵ�M�'^~ˬ�g$��lO��3@+�z+���X92��6B��w�j��Wh�fy�8p[��ϔ��&�O�N�
�;]�5�'��m8$�\��c��q����:��ۥ���{/�{����O���ߙx�.W�9�\�r�s,���Z�ᒰd��Y�
��=��	�gn@w���T0��
GD��SR��$��0�׍7��R� �s#�HNzN���#3n���6����B��5DB(�b8"����D3y����ڳ0�w���ڬ��߭$����FO�#z�+���U�m�A2�MaM��`���b�����ґiN��E+���)S�<|�\3s��5[X�A�3��g��
�B�x�I�\W�;\��HZ�ղ^h1��AE8.:\<�o,��!����Wav6��l�ȑ6�Y�kn���^ۻ�`��9J�S�F�s`�"�EJyq�'����y�5����ml2���"�c2K������壵gB��~�%&s��&��v�����7��r��Rkw4��E���&?x�c�ֶF�@�	�N[ ڔ����5��+M#�Y�6�- ��׋����E�8��y؅�fO�b�#�B	� \�r��)[���u?)�>��h�4( wg;`�jܧ� j�F��U3g�xs	�7�i:�7�X������N7�\�w�}p�t���E�kAe>��+�T��.��e�#�b	�8�ʹby H�K��=���C���ic�U4��3�JT
�;s3\����:�#@	P�M*%"�ɳ%���%�Tp�	Hu���1s㹋.�������Q�;�P���z������h,B�q�����6�8JSs���Š�7�و�N0o���	x}��]��e�	6��MA��8�;+�9�_\x�7���+~|���)�H�_2t�X��R��wb�rEr��)[�v�#�2�-K�LcUS�����NF"c� ,(/:]��/�՘���\�6m�,Y�	��1�91^X� <.�cQ�SiSt����r��!��MZh��UJ9&�5ޅe��ĵ��D������7s����J�7�q�����)E�4
n�Iћ��Cb̬6u�F;Tp�����bL�P�Q�ԛ�*�S��/���p�R��LgC�(X��ę8 d@��g����¥�;.��2P�8ʀe�{AْI�ڣPw���#��� �p��0����	9�/��:�ǡ49�Iv�_؂��r�N�q�������g��'8�
�5r��Bo�s�ϸ)�nCC�㜧�W����5֊FV�i�Ń�;`,J�n����dɦu�����1�M����p��0�����<��:�Ȉ��Rد�o�v�)����������"����7/]������8n^�߰��s��� ��Ï0'�t"`�4�]�L�)/�����.�e�,,D=���m��η/����_��n�>=^.�p�
{$ҚPL[�h���Sq�H�l[-��q��B���8�93�&�$8�:Y�rs���d��-]�ws��oV�Z	����(No�H�"�M�S�Ƙb4h!ى��\�TJ:���M�`��
G��}r�[ڑ� �Fβ��3G�o����U��DHV��4���LBg��0'3ft6�M��pq��I�uŦd�J\�Y�w��fX����Ŕ�X݈�ˣ!����jw�7?S|�2( (��*�u;�d���]���8G�U�%�y����@�zw֬YK�����=��s�:��פ�9)4�
l�)���8'�97��+����S^;Ă;"�)�B���@����C�JNNɲ�L�2ͬY�Ɣ��~K3����'H��M�R)���*��Y� ����x��W��Bl[����c8֯�:�c����7�u��gݻ��׶���m���߀��m��v�����U�Xԥ�s�f���K�bܓ/.��0ɰ�C>q�Ds�Yg݄Jn�-[61#=+މ+;��E�	�)6��mmm�;�J����Z�<�&�B2t������7����e��_R���P�f�8�P)�n-s�E����C�1��Ea��r`�O@#G���]$8�����L��1�Q�&��N؀E@h%�\�cڔ!�����Rx����k�.o��v�������|��K7��{H_���_b��oX�X�/oEJZÞnX���ᾬ����M�?0�4ɣQ��Y(��_�,/�.@�����s��Pփ*��*��Tcs��R溯N�T���N9�1	\8�q�1��[�`�KӦM[e�mW?L���૯����Y�v79�s\$1빀��P��7eQ�e��u��-HC�H��q:��N�n�斐�h2Q�n��E���:ʾ��q������裏���O�O�|UOwʒ犀:P�z��ro�>y��I�^���($ ��m�rYY�&���+|<{M��>�?���x��L��w����x�V	h�j	*V[gn7Z>�j4as|�z8��n8�E�yǟoX��	�Z0��#੅��=�����H:�RqR��)h�NZ����/����"��s.4t튔���ʧ�$�O���2��9��	���[}+a ���1�o�1� ��R��-vZcښ,R^��F����x��_ZY�^�X@�beJZ�4b��$3-O���j�a�u�ׁ-]�l{ih4EQ��М
sP~�dB!��1-(���<1�T�45���ac�������7�N��BE9i7A�GE�7��y-��h��T�T����7�Z�����{J���V(�����}	P~�+G�r��a�6����W���G�0H��4([EEe���S �>�=�=��x�	�n�������\ʋ�U[_��}9�,a:���b�KV�\���<�����NzZ��w��A�|߲�?���3)�G���~����ӟn������/Ld�	eR�: ��p�*�l���<��?!PO��1b��g���?�ub@��<@(O�7��,�����v�A�[vk"���Ȅтbc�NP�.B�b�B+j-�rOlkm/�%��`	�ڶ�օ���<��_*�A���������V������zܗ�%x@�N�tO�s���"*��]}ͺ���| �ؑ�d��E��/�-]�4R�+ �5�e�(�K�@4@��c�K�r1&����H|:?"���]P���66Mi4ݝy�c�Q1l�e����7f����1��m�̫MEsr�f��7��U���]&D��(��E58k7�����|�����j��{��������k�El>���A$�'�J�%��al��V�NZؼ�S�4	��)?*P
-p)G\1_e���YC(��f޼�K<���	���Nb������g�s��?q.�CL�o
M��S6�Ӽ6�w�znB��ok(�K�R~�p.���>׳�p��\��\�&�
`����pᾶ&B-���%mo��JZn^n��׵a���'�xr�}��w�<�a	�8�X����f»	�b�k�"�q���˳Ń�+X�/#���y���^����/*A���L?����Z�s���/�(.F�l�w`�`��u�5�.vwb
����J�ꪫ��4q�+ �r�߿��c�}Vo4΃�Xj�b���P�%�*�Lł`�Jk�4gQ`��(���0݇�c?p��ݮ{
���uυP��]��U�BDr-j^��BL�Eb�|�M���\-e5g�eo�ń��Ѻ'K����F�(����X��W���l;�o ��c:cM�Ժ}pM���}�����o��s@rZc���Ms+��m�t���o5��ZL��P��ף�	� ���T�*͆�Rsϋ��
jhI 3� t�0N��c��u`�k1�uĩ�Ģ���=���]Ff��j�Z��[�:e�+v�c���̙*A�YT�s�}�����pb�F�͟�`%+����;��k��n��e��ЎR�x:���~�'�g���%J�+�CJ����;ޟ8��f�$�͢E��������5��o�����7�]����Z��q܏��MϨ���\J��?��y�����
%97�CC%�!�sh�wܱ/���pvخN ��<	� )�����k�_�x�f�������w�5L�؏���\a�I��R������߼�9�lnn,�4i��h������WcƎ�����[O�;XkY��˚9��\���:r���ǎ�:/7�Z�<
G�:���e��=�>.��'7����4{�tsR���@ke͚U��w�qJ�bg�e12�9*"��qNŧ���6�`��耕�� ʅ�<��إ�9�H�O�2�)hAZ0羐Kʦ�z�f�?*e��w��&� e\��u�(�g�:��h&Ƶ�#2͔l�SaE���3�E��{���ܼ�v�y�|�op��v�c�*D=�T?*��b�J�������AH����Tz����e��p��������F�t�"����i���/p�O#��IȬ��;o�m��?����ڥ�*���v��{7!4�"�*;Â>K�R��|d%<�<p�wL^)d����c������b>���N��20�32�+?M���������=��?��G��s:��h�á8x�	���|�\�-"�\��Zʀ�}�hI�a˽�z��&���?���1uꌒO����-a��;L�l?������V�̻,q� ��^-(�.֡�Әp�H; X�Q�>Ǭ	�c�3���QI-� ���csֹ��ݖ) �rā	��0�ٺ�m:XXy�e�ࢅ������.���΅E�n�]��w��7	��uƱ�d�R�E6��Z� Ál^{�US^ZIR��r�KW{ܜ�F��nD����a����kh`�<�T�kHM�0흭H/*3=h�d�cCae��k�q�)6ͺ��M��Jӄt����Ob�9���IG��J:�Ւ�Y0��X�l>A���N���.�G�]U�/�(O��x�N����-!1�*,Txĳ`��VX�Z�e�iQ�;�ߋ��1� ?��<>o���?Y����� ���KsO:�3�a�τ�dJ咗B��gFs�'z�4K���0g�q����#���%[��u��	�2Ȑ���Y)�it���aCֽ�ڧ/!�b,�*x�~��������w�|���5���"��ǨbR╈ۢ��-���OE��eKS�Y�n���W�z�__;��c_����=<@�q�����%����_{���Ag�S�W�[k����9]��J��c�5.���U�X��ASC��NG�̔�s�>��|7�|�d�t��=��6טǱ���+����TEk���[nF��3����� O����	?�����g�Rk����ff�8Ÿ���������آ�nz-N�:��h.vT���W��b�}eI�]����r�Ғ�8x#�����O�y�����jB�3���������`]��*��!��5�S��A9~3$?F컭�q�n��EBV��|�n�y���x'����F�"a��.w��S���P��<P��ޛ̬t{h������[l�G\�y|\c5b�Ϟ�կ�v�!��6������c��W��nb^� ���VQ�K�DD0���:�ox��]n{�,c��-0/A�6�y���1�G��,R�\�d������+.��O��y�s�Xz��j<�x;����Bb�,����)á��կ�Y���c@�{ﳌy{������w��*<P=�ȣ�t�
T�Y�w4j�v����p�>�xq.:�'�п�'?���^x�S ����*:�)ϝEVx<���͍�xZ�|�x�;��֡�#��"�Ϩ�+��4$@u,$�ղp+�1昍�pz���u"�2�1���r���b h)���J�ʎc��=g���C�q�*I�6�-^W_gA����D�	a|#�3�}�$�0]��W�WA�91�̨zshZ��7��dgLb�Mkc�iC�(	I�٦u ��_g]������ ,��}����eџD��B���=⵫v<e��=�	zkTz�2�X�S8k�9^:��w���5zT�}ܿS��:�&� �s�7�g[p'�J�T�`��E2���46�OV�@M
!����t�D�ʒ�ou_�'�2�s���/�g��w���%�^�!x5SĪ�xںN=�r��y"�Ze��R��\vv"T~A�lЕ?��#�?���t��;�^���z��]!u��E��6��_���X�sk�c�>p�u�{.��(ī�r�"����t�H�ZU�h��	xTD�!�ۜܰk�����jī[P���Av8�y�|-V�b	���� v3��fW	UYC���srrMNv<y���M��A��z86���o��e���G�ʋZ��M����$>UEӹG���Z����+�uA	�H�fg�@���L���P\F��^�5���<��4y(��wr�9"��$%D���Af��OЈ�ˤ�K@0_�z�Y�½��d���܍X}7��l��c2S�L�i289�GT�xo��y���8��H�b��fy(]��Sv衇������ìٳ�n��9�b��m�4���-��G�S�w)/ʅ �9Ap�3"��gH����"�Q��;Z�8��P�<�X�W��s��s"�Rl�Ǐ7�����?�>v����8k�kb�������9c���xw[��Y#7 ܤŖ��r��
7v�<�s�	�Y'
�amr,22lv�'���栌�N�t� ���ﷻ\�\s��񯃰6��7Y��lw1 ��Q�Z����D�Q�X@��n�ȳ����-��98`ύ%dŪ�BG�� �B$t�%�Ϸ\�<��)wYS���Bb������@����,{����0_!��iH�c	�yM��xN�������gmA=�);�C�0!)Ҁ�
A�y�!��Y����;C1�h�1f��SLF��Q�V��$�J/�i1����i3(���Y��)q�&5��D�R�Z�� ��O�����v0�{a���ݞ��j[l���{c��Z'�S�+�����]��2��֦�#Kp����B�љ��v�~�������?��m�=�q�G~�9=�!7��N�ܙ�*�C@�$w<%�� �߉|���K��� H��7G����9��<��(Ϫ����Ri�q�K�6:�^��v��}�u���;��s[��yR�� �+_�a�X�-�8z�.m��:��w������;N���L�� �3���y J ES&���?��{�w8�d�%��  l���hU�=��᾵�3�S��%ښ�Ȼw��Ap��a����࠸c<��w�>��c�x�l��I�bq?ܜ<��V3e��Xyl\��E@��8�e:��!I[;��XeS�x�!p��7����%-\��Js~�hw��Q����U"0�p^�%�����O@�NUU���r0�[a��*���&*�Y�f���؅g�삡��:�XSe6�Ԙ̸X3)����fƤ��dTr!��� N����yk�z��G+���t��Oiw��y&#�]�@V�:`1�P����`T���	 �u�J��I�:�G@��[\	`*p��Ay��Cy�c��wʔ��q>o�1�YШ�;�U�@V�C�s���c� �SV��X�Ҷbc���R	�����6����˱�����|��1���l� �M>9P��j��$�q_0�M	�:��'�|��%y�7?������Vʮ�L#�|
|���uL#��F�C�)[][l ��`�g����ݏ%�SS��i���������;�R� }{��x�L���#P9�&��p�m	n'M6�F���P�Ÿ�sQS읋[Z9��+Z.��S�Pq5�[�o-^t��1
�u
�p!TS�m��#���&.W)���$|���M�<]�UU���;�����*>�")��vE�P��zXh�8aM������˗��o� ��#[FL��=
9�Q�f��#�轎B���Yc**�͆�&��}�M�5����4��{:,�~�� �t�W��1���R���2���q�yH�L7��Y�el*z�sL��:y/�P�n��QV���	�^��)!X���:&O��*�p���O~|�MНxb�ϣ<���&���ͅ�弡)/w}�Vil6�O�*Z
��󷽣͆<T�My���Anyy�� td���e�����V��Xi� �Eoݺ5��.��ٟw��@v=�?��𜧶C9W���y�a���	*9N�%֯wJ1w#Ã�V]PVi��svN��={�_�xӭ_�װ�cz���$�g�H�tsI�W=���'��8�-����n�j���)iJ0����+�G`��[.l�ߨj����?�@�"GA���v�Z�`�ߍ߫�]�<���&92�YE�q~n�xMؕ!;)w�7;ʉM��E��gtw��gr.����y9�u�ט�jt���<D�9/=,�j����a�N7��:��b��Zo��z����$�(7/���^b���9���'Z 갼��2Mo,_�ʼ�j�Y��{����c�R��O���H���F2T�.`�xB��TFT%�r�Ti�X|�-Z��q����G��N���$�����/��tC˩��{�9�yE��F˜
�Ȟ"@Rt��9��Y�����p�Q�U�.��ʘ�6�e��]HKĘ��)7��2�:��cC@w�=��7�=���A>�a���{n楗^zKue�L�кr�-y슧K~N<�U��VH����ˏa�gx�������2��~�e߽���v��� }gH�;�.��m��z&������vL����B���c=���t��ݵ�is���8���?���\3rT�P�խ����}U���ZV>����J˅�DU�Jȱ����a���
pp�)^���$���	��u^Y���'%�v:d��܏Vq+�����d�4��ɺۻzRʹ}�4yc6���l��5k7���Y�Ro�N�1c2�A��X��-+7�X����ކ�f٦S	K?s�h����@�h�Q^�
��ڝ~ٔ+�#*"6ޏE��V�9e___��)��SO=�N��e���w��ۅ'=����[�dɩX葼p�Wy|8���9������fΜiಷ��2�A����	�h��{ �'����n*L�yi�0��tI�#��58���NT�k�yH��}������o���b#��_;����{�8yt-�J��αp|t�b� ��"D�kb�%��N�!���FS��}���kG_�����%��I���W�����r��<���Xx������Y��)I���J-��h](��A� �:�z5���Fp! s#���$cs$��"��]�u����z�g�WVd�O�
3����d�x�F�%a��8�0�t�\|����g.o���c��F�e�J���zPծ� ��E�Jcu�R�&�E��q��>Դ4��k��֙|�}�/���I�B�9+�!�9׵5��A#`�Ś� �}��χ9�KGEE��*{�1mp�Yo�F���8��O�e7y?��ϰ���|�����g���wΝ?o�5?��.�{���P"cr�d���+�#ƶ���ܨ9�,�6��C�Us�>/�6��C�_$T�c�KD���*�W
����x�`�ű�N:Ƕ���o �w���,/+?������{�E�e��8'፟�l��xt�;�U}��^Jk�V�D]���� ���o�MYYɋ`�;-!w��Y�;H��a�^}��9W_}Ϳ�p��c	V>�|(	�rE�a�@Һ��=r�����>MZ�d�;ֿ��*l����ӱ�/�<��i��A���	Z<{C�Y��.X0R�Ĵp����C��4��y��hWa**g�e��87K��%��òo�h �6���cf/6�g�e�1X̸�r(��Q���LΨ�!�������B�=��5���>�b6ĥ�ެ<S��|%����@2
�?���IOMO�2���?L�\*�1�J~����?���{/\���-�z�i�CF��/��ַ�u?�Qʷg\�c���U\Gb���RFQ%�r��Hx�&)��)����TUW��"��TH�S���X�}���t���!C��[�:��3��c�����o�i�c�9�"��r��xŏ��׿��G�%�?�����g�W���IK��*�Dǲ�\S�������b	r$�9�Z�����X�#���C��<�wlO@��6aa��+��]m>i@֓@Xw �z,d���̅�1q>�	��q�=l�pk�Ӣu
v8��	�Yٙ������$�y	�q$�ѝGmR±FX;���`�ׁ��ڞ�DN.ݔ<'�7TD����@[�:]�P��~�&L�cg�� I�w;܁����F�:��k>|<C,�x��f��Ֆ�܁���.���$���`�.8�O<�$�e���ëŔ��ƶ�R���`�g$����n@cX�H�1�V�[���k�L��[�̪����o�mJ6lĵ`_��A�7q�%��R�@C����v��ԗ_��cȰ�{��y�����-~���O]|�IO~Y��'�qƙOc6�b��8�ݠ�H��sS�R���h:Ja��k�tX�~���d�X|��a�SMK�yH��N�N�~��EY0_�,�	��N���sX��<�~���s��ߩ�/u�/.����Ȼ���gӲ�m)�z���a�'0����M]�{����p��B�o�eK�9�w����yQ��}GJ�;���@CC��{��裏���,Z�L�b�]��@B���̌,�"��"R��ÊPa�.H]9v?.vH���b�q3�!����$�<����$���[Ak��apHq%�׳XL�P��n���p&k�nX\o����`^�~�h�x@Y�`C��]�C�?�-z�fc�o��C�cL��i�C`�C&	qP&z�`��bc�Y�E����4�v�?y���d�՚	�Xؐ��女d��d�;h�i�b�^����'��@��7 G�´:r
��q5��Ny5"&N��K�R`Ѣ�O}������~��b��A���y ���Skk�'�&e�Z	��� �:lm�ȓ3f�h��t��l�8��v��΂;�CV8�߄�����n'e���=��{  w�fs��v�a�D�}�C�N�~���x��׷�t�M�w�S-�[?�ӀƲVmJ��Z��"��L*��a^�s}N��ɻ��1��G~�G/<��x�!iz.��<a���\	��T��g�_�<���}Ԫ� t$�0���+���(/'ߺ��p���E9y��W��K�2��1J�R%������6\!�)��u�k>.�Xq�D�&!M���{V�R�T�2��
�XX�����qqd[K�Д{^.�I�<�.�W_}��WׂS���p��e/�޽QA���3=�If���L��CM1ܩ��jj���h�:6��`�O��������~��TiR����F��S���!-m��ʹ���$()�P�Z�|���>|8�?�J�w��ih�+��.d*����}�W'�t��Ï���<�Y�(4D�L1oY���W��	��D�t���e�6m/(��lZ��*����NT���4�@�9�9��t���D�9�V���9�&BTz��)-���^+���o�묅�^�sW�-�������]��(Ŋ ��Q@l������g*��0ߝ"F�n���{�r6�#a����G��#���!U�B7�x�%w�}������Pj�#8;��v�"���E.>�"A
�a$dq����{.d*�︐��(V��SN:]r|���SNӺ!a���
6�1Y�~�6~I�A�G��X׽�7/��E61��s��r�8�%<!&��s֦�}������R��g�,��6�],�� ��k��r�N7�f.��6���K6֚��(�\n�� �R�ZZjLBZ:�1���fMI�y��* N9��':������<�^X89�|�8��@���/eh�0mP
�u��}Gy�Æc��z{�����~-RgQNt�;�B���̹ƹ��h�)<$"��o8�gϞ�XvBG����-�J�T� ��ιEœ���*�|Ye����5�P�?�*�T�<�*u����y��s�=s�@�����E��E}dm������th]a�HB	�c�M�o�C[�����d���?�WW����~� } �o�U��{�i��r�� &0�����O�v�ňV��<*�V.�-M��Ō<��$��L�Br�ӲNAL��LNN*���"*7(Ϝ�<�̙ޖW3�ϱ�{�u�W�WF�{��l�����j�GP���b�Sa ���/8&ǧ��B����-`�-[q�w!t�{�_�c��4)��	f،��i'���[��V��}>����H�5����:��64�io4���ǧ�Һ*�
�i/yÔc-kE��$�,�x�bР|2�[D8a	�,�g����ϛ7����k7}�1�ٮd7=���k�����_~�4�*Y���0����/��T
i��X
�_�7���g̘a��ꙻ(��Z�3����,����E`�W�7�o�&�b���L�|�R1����2�fS�ӈ&=�����>����(��K��
2W���u�� 2DʑJ݆�p��7�t=�v&�X����Ғ{���t��ٞ���з�4�c�R	 ���U�+���d.0�V����C����U�b9Z��gαV9]���:��)`��)A����d����cFR���fIIg�uj<��[XD�|�%�pa(-��|�c)�@�{��$W�������2o�3��lZ�ل$�@�=r}s*+\Hy,Z�,N��(4�HLK��!�[jZ���M���`Q�aaj@�U4��۵��Sk��d&ܤ���&{�00~s�ƪR�1��=���k_(1�$�P�w|6ھ.0`�3At�3��c��׀�\t�E�������'���>����o��\�之�8ȉ`��r�~O��q�s.�J�x禹?y2��b�pNp.pq~)EK�7�<T܏�г$��"���@/��#�G�=���'"[�G��
c'��뮽朳��}��'���6[&�	����/��j?)L�G`�2;�3���&E�}��?��+�{,��89�S�8	<��#�/���%�2N��sX�|�h��v�]| f$��$�PlI�p~)����e˖Z��'9�+!�Km�9L� AY�K��CL�&I�@<8����4��Y���:�h��W(5�w�j��jj˺wX�Ѷ9�!��#�VRs���HHmڸhҽ΂:|�b��9eT�̵���Lˡz�TX��!3lڡ�`́&9���A�W�r4��u�}3P ȵ$��n�0\��f%B������KL�#&#�x(p��AE�`P���|E`�w�ܔ!�\������׿��?��l����-�ϑ�����7o޼'���������&;x2�I¢�I˙ ��B��K�n�m�~�Y��e���Axݺu��F���8��3k�g-N���*�B�@2,S�;����y#L���|�|d���犞$��"�s�S�,\�N������W_<uڔǘ{����w�rؗ�7Q*�s����ԃgZ,�I8
}
YqzA�Pt���r2�����R=�����w��.��e���u��'t�w�Pei�<�A�J���?��"'��?x��
���,Ɉ�:P-�l8�����6�6/�T�	�v��� $�{���V	��ېrD`�e��ɲ�%���UG��CQy���X$�npN1���$�SQ�V}���R�YԠ���l]>�Uu-�f��L���LA�������`̨��fJ|�Q�d�a����M<����5(���+��o���.�&:5Ց�����<���6&����l:����Y��)S�2�mpE�������~�k �$Z��4)�Be�� ����~������9�qc�Z�7�TD���UNWmsٲ��!���D�%sN�8����[2&��+���,Pz�HI\��m��=ǳ�����\}4�OĻ�C����a&+��9str< ��BY�P�b�ӓFy�����uF����|l���fз�$���t	�y睗��?���aL�b�t����R�����+e�z��J�6_�\�r+�=΍�7 ���mrS�s��"�'xh�T	d�Q�tÆ�va��{,�6
�,Y1�ݖy:ڇN�4�.b�;g��;Hm,$B��,�~"�r.��o���dj��rF��.[	]��+JN�ɟ|�)�z���-@����5��P���Y����YP���[�ͤ��\Y�h���G�T��J�A�=`za��K"��2�=���YN ��Ds�aC����s�v�y�8o�4������Vs1���b��1rI;y�H����`��Se5�1�v��99� �T(����s~q�*��1qr/�Z�3�>�J[#��8�	b�87m&2!����>�A�d�S^J2D�`�C�^���o����ۡ?����=���{
u�Q�͂5e��v�i�Q.���sn@1-�32��g��Ӌ.����c��o)z�ة��?�y*�o��YD ����`�u��L�@˺�[,L�~�"��E��16�X#�_��(3�׭A�2����7v� �S�Z��و�MM��o�``�&�8�����/��{m<��ظ����5����cĈ�P$����1�?;�G΂���ӳCT<,�dt����D�	� ��d �MV���Lz����^e�'���,a3�T��X�P].@�\��-}ǼU�ҬH���;8�UVv��ۿ�aE�ݨ�t1a�7/��ſ;���<�S'� =��{#�� ���\��,��Ls���"�){BJ��Ys�s\����$p�g^���w��(���C����3%eR�L~O �3�g�n�M�<�ȑ#�"���L�ٌg�uz�# �����?�0k�.NUۖ��삋QJ������[Z�tǫ�]��l@#/�Brtǧg$�������ζ����������&�����?�1`Z/1\��R��ۉk9���Z��Zw�|:�H&8J�Ǳ�L��L��2N9d9�SV:�����L���7���'[��I�)���z4ae,����4�&�T��w��U�E�ik"5�˿:6��$T���������D.��\TPı�:l�ϓ��lZI�KD���}̰�G�!y�MX�eu&���,H�43S�L��tv��^tע�6g�xӌ���7���zݼ��-]�-O�61i #�ӡ؏���VoCzeEE���ɵ�����촉3�O��� >�x|�`�%+u�s@�����P>��Nn�U�s���A�+���[����G
+Zu�\�¤GI�,��96~�����:
Q�%��J!l�����TWV�����������ߏ��i��-Z��S7l>\���2��nzP(?�Ii|b��_��"M���yp�}���}�Y_T�Q	z��)���[�BӉs���ނ8�"	NV�еh)7��Q���:Q.�]���򷅨�FB7�80�m��;����Μ5�P&Y+��n�z�uwd;,]�U�cڪo��k1�EC눋%��)�U����4+����y�2e]v��ʚ]x�H8%m��ʈFe��9t�)w���jB �JS�i��2���f��z4|pɳ�l
��u:��g�2�j��"v�OF.��ňD�vT��F��{M����_��E�.|w�L�z� s���������cnL�0�y���$}}��<9���:����ݽ|���^�P�#��N���)Tz>��&~�H���vftP�\�f}�9���j����S�{M���
y-����ǪB�7���fC0]����կ�;������|��NX�<c�,:C��й��2�ʒ�d�m(���/|:_�N�ה)��|9xik_Dz�ow�Sw�]w����?��mNuQ��Y����]�u-nZ��o�sKF.(A��̇����*a��2���S$�	x��������#������1���g,I����VH�����;����ƅ���&w����s���
�V�d�Z'y5��(uI�ǔ�|)���$��u�D�3t?X�,��/Uu&���L�.1S��L^~�����fr�Ơ�j�)�Yk|a�Y��ߝ��f2�w����<)
U�P|��B=ʑ�������w�r�=�̗�������_��:��pomE����Jo$��I�9�:���V�.�^qpek�9��2���R)�|��YX9P�Ws� C��s��@$���sP)��g�s�r?���k�q�<?���PoY��|>i��w'0�|ƌ�t�-w��?��Jݳ<|�p���G�Q�7P��@�
�sƚ�t�w\�C��EU�B�"��~��$�~��<���t����g�!�A��Mz�ūx��*Ң�\�d�p��qt1���Œ�4�m�jT�"�N�:5� �\��NW�8��^3��uʙ��K& ���K��b�9�r�y�n�ŉ�a���G����/^'c�����G�jYn�~.��Y��nb�M g����)�EE<����T��P�Y�TkF�
��� L��.���s���nS����1��(��;�%d ^g�ېn�q@�h>餓���%�\3x����m�<�̔G���K�,9 ���  [;UJ"��=I[5�E�Bj㵸Gnֺ��n+[<��	���$����G�����{�u�*���8�8߹��|>��|��s3Փ^&��ށҒM�
"s�QXi��7�iވ�whK�5�8��O9Y�A��gɟ�*j$*�_�<'��e���B����͌�s��y���畜��"XI����[o-;Zk��F��2O*樬-Rr#:�`�����|�TЂ�&$) *�b�Jw\RqKV���|@QW<���}��#���Kp�*7>��6�����x̢�B����xi�G�� V)(��Ɣ���4{///���R6p!YN��3�n{Yc��At�����!�\�Վ��Xl��7�}�JͰx�Wg�XR� �� Η��0U���������˦���f�U�d�R��c���	N�>����?�3g�r!�I���+�����_}o����g���H��-&K�8,�w!�;]s��R
t�#s�6SqJ�r��[�Z+2L�s��o[�K���[1c�*'춶5f�[`./��kKG^<z�x<�8H�d����j�~�s��g�vک���۱C]^^��OKJ����2��������� �@��H =@¿P����II	�'�cf͚����?��=@����~��%����z�+W����"�I��	#����%�o.f\P�Pq�!���|��^#7t$��u5d��?�-�)|��8�ƍ�@�җ,'�V��sX��~���#*q�/�˱�4��q���Ij"���y���s�Jv�5��-)Y�v�gw(K�������Z��}���?Ɲ��숷WT��P����lơkZb,΃Jv���:�ǚ��B����T�;��O���r"U�9�Rz�3fZ	e����7�x�)����>A��~�����gb��90�!���B�➋(���7�nX��yUt߬�
k^Iq��W@-�P���Ir�K	�8%6��`N���y�yF0�<�u.EU����ܧ ��9�S|�/_n߫*+p;�_|衿0@o�6��o=�׿��_��y�ć�3K@W�&~�6��J��g��S ����垱EEC��y�=@�<R�~�]%��[o�E���H�9�D��W�T���oG �K\P�)��pT/h��i�<� NI��b�e?sw��]j�r�sw��w����"餣����q*|�'L���Y�ͩ��,0,'�"���2�yi����+֒҂��|���*�BP'ܜ�&}�L��
n�NG�|H����k5��&�x�� ����`�R\Ee�Y����zs��Gw8�r5��ҎX�+�Jz��?�f��~8��ȩ/��n��ǜݏV8n���=��P�X�\��}˭NPלp��#$6���a�<U�<;?�Y��r��b���j��U���pϗ���,����[�LJ$�#�o�2�|I�9�+�����(�6���_�1�k(,̯���r�A;���Ξv3g�^�F9*�+9�8Ke(=-�:?sg�صi�d���I�߻���r���:<R�瑚���"�_�vnD���D�n3�!q����t1{�1H-$\|h	��"��Y�Ņ���j�ld��b��.~ȹ�"�ŋ�b�nr��VY;<��EN�rUmcr\4��M,v��m�o'��8���[�o=Xh�"��HZ@$ڽ��H+���-.ȱ��˭��!�/#����0�Afk�3�����SlD<,HXM�&M&3�d��٬D~��/-1� �2�4 �Δ�"�T9��ښ�����N9�+���o�.sc �f2,C��C@Ҝu�@�ɐ�O�A������IcyV���BC�}H��]!#�L)������a��d�t����n^�I.v�_��"1�W��R>5-s�s�Mr�O꺩8R����U��ǣB������ϿsOsރ�O>�ϨV9K9�7AN)]"<Z	Y'��f������?�{�@Z9�DcA%��A�6���ϥ�,6�8��~nқ��-y�9Y�\,��	�����l����'xҊfE��%NaY��=-�����s��M��Sy��f� ������v� �u#f�m].X�$�ECA~�yx���B��l�p�\�>^�/Ή�R>T&dau�AЋC)��LB]����dFf�m%##'���Eq�6���t�)A��>\n2�!����6X8f������<������U�:x����}��b�����F���p�F��d@�9x�J�ï�.��<A7�S*z�|x��Z��r�CLl��9�qh�U�o�?��V DԒk��s����3�+=������q���%�3v'de�$�[n�FG�(�1g�������k��lN�4e)���)P�w2BX\K���;>�T��r�ُE�[jj2֯���n�e�iӦ}������%ã����<��sᆛ��'w��b��Rd��ߊGr���`I���e�;\� Ŭ��.�a�V.2?%%�&[!&�I�0�ƶ�/�ؔ�[=j1V!��X#��ey��LSS�s��U�&;'��C��C��9�0;E�n�-�ِXD;��p�e�7��Tq
�g�9���"֦?�듻���Q�>��2�U �E8��T4G��1ñ�up�٦���l^�٬�,7/�]eZS��x�Ow1���5����˯�1s�S�n�o�oL�7aH]m]!�e0�a$HZ� 8�p�
+΄S0? r�tos�?w��E��A]�k�A|�m�1�T�@�Y�n0v[�[�H�����r��s���ЇPq0������r�#����S�U�W�3'&��}9W�b������;�B�	�#R!�O{��+~|<M�|�|��=��S�/��%�2���)�dSY�=mϝ�gk���=2��Dx�X�d҇��Ǜ��Y��g����� �1����E�0L�(�_8
���B؍�^и�
h�TE*�Z�K��K�ƺÅ�;�5ÿy5��9xQ�u����h�Z謟N�����G��Y�B�s��"��b��ժE�V� [��+��q���uӑ�
���7�.i��l��ꫯF�o����.r����$&�Rө'��$��u��b�p�������	f(< ,:U��Cqٰj��@ј76��z4a��eA�V��}�ٿ��~��&��rݣ �)x�UWWX[˺��dpuUu^eeUa]]Cd��W�@�bǊc�]�b":�	����,,��݀��d�+�#o�b���\�w�<��o��=��b��IϏ�E����"�����p������3T&9���}V��T����%�|�H��<��Y^Zf;2�d҂���W_��Cg͚�nL�q��=���+��uMJ��MD��p�եQ�Y4La�@�'�����9	���۸y1�m������5kG��_���W��u�ʮ���{1rz��n˙nb���gd���*U<�E�"�^\Y��P��ʶX����,hFz.,�,,ΌE��m����8-�*:�4Uq,m�/i�нFb�R���E�c�΂"��2��#��T(�t[rq�9�~�w�@�EҐ�Ȱ�,D�F�3��c�g\�)[�<��4�d-*u��4��,�C��<xV�^c�˜z��M�ɦg� E�Ӻ��)�Wv�a�}�ٰ�%� �$C��M����mmi���]d#�y���Ȁ���<����* `�@6�\���Y��,lyS��w�:�`EF�:�h�2צc�w�[**�\��-t���Vf5��τ��
h7��@ǰJ�kӼ�G� ���2W}۽�	��4�w��s^����-w�=H�k�N�V|Kk�u#�~�iW��`N#���\��
kh��ܢ	��D��y�{���c�.[��H�35-�,�m_c�=����f ]i(�gtee��2'�zf%�d|>�mj'ܹ\DZ�6�X",m���*�ՠ�ʭ%�Ea.8\ű9L���\,e5��N��"��	���󕒜a-��6��D���0�V[2������l��$kQ+�.��O@�I��VV���8� X�뒟�<\���%^������;n�C�-�@���2��#���)*ա#����1G/��5w�Y����p�++W�(��\4����U+�1��[n��;��!�|I��� �����ИMw8�0E��ߥ�E���g�EԽ��ߺ��X��I���5G$'�ce����rY�:�[!�}�����F��R�k_��-W��`9a��[�u�#�uK��ޣp'5���`�χ��34�����a]s��Q�ܧ%<t�6]/�����<A�~zqZ�Z�[
uΜ��v�m�n��3Џ1~�� ��|�d�Xe1,�=\�O�� �:�S�m����iio�.������,��Y�EZ_�}1)�����
*�u=VQ>����r�Y.^� �"�`�Qp���
l�V4犓�e9+����]���є#�;�Sk��3��m�k��Jq�B�ŏ,s�ީ�J2XK �7#Sʜ��P���:����c���h"���mƔ5�Bz�j��q��+%��HB�V>�#�LKO��O�U��(+K)1:'�!��oAN�緱O0gE��T:���Р�(Ѳ��ġ���k6�,(5U�fCjקe�|�
{L�;p�7��oϻ�?�m��q�a�$���Z3p�4|����&�&�����BOY�hQ*Ɣ��X#����&ݚE�}�r�~�v�qa]��Nƀb�:���=� o���厗�).�l�ѕi��x�����/-R64w4_�f�Km�Fc��(�Oig<>�5A�
-9}�����Y��nᰛ�I�t��lD�����1|����F�����u	 �K�z~��g�y�ͷܤ�.Z����rt�?�r��;��v���J�Ұ���,�m�����,�����
�!Xt���B�wp
���*#):pm3,�ablƑ�cީ۵n�Y��z�Xy�_�ۊ����x;�y��X�t���N���W��qGjq����S�]�SV�b�4�jM�M���k��:S�fg4[���E�1& t�	c���QW�k^S�x�|��9=��#��CF��/������S���0kٳ ^* \�U��Z�PVxn��J�v�0�V,�ԓ���Yf����
l>��=䦇�z��n�G�2�1mZYRR�jȚ�]<�������x4�K"d�K�
�B���:���ܹν������+�(�hgir[��]�n/��x��<g_U=�|��]��v��n�+Ḙ��q�c1��:���#������GK����h�)���w_���F�Ĭp�Jϒ��in��?��b����2I)7Y�Mq�fC	V<�dI6"�U1�̙�إ�^r�����8�����s�~|�i���yZ��f�x�==���b�Ef�iC���<�7o+�x��Jj7ܯ��.�dZը�>���z-)<xcO=��4,���sk�bpk�u����ʉ;�B���<�C�5�mI��5)�[�:�1�b�];�@�9Ӷܮ)Z�\x����x<�դI��wt�+6�p�:��	�:�m�����:و�2N���p!�n�E�硋���ֲs[pvP
ҕ�.M��m��Aȩ��Y �Q $� e"�X:�v&�_2�V������˵^*�`�Ӻތx�;�c�抹[� ėض�[���ܧ\X��7���V�
^�>vZ���u)b�EP�H�5{.s`�;�X�׃�~��pi|E,V�"�z��`6(�(����t8�̶Ly�}�f>>AG��l&b7K�$GЉ	[0d
c8�+�U�6eb��n�츁�$K~�l
[�cs+���g]��l���g��jv�� i̲��ˍ"��=���?���ܗsGU��%�J%�@�5�9��	>H�2H��D�;��9�y˺�	anH��������AFr������l`N�/\���Gyd��GIu8�/��H�xԢ|�&�}c�K�y��gN��<@w?{�ߛ7��7�5�u��Ԙ���ʊʡt�7��dASq��a��	0�m[��;���m�0&��!�8@LL��s�UA�NX�Z���UY�<�KY-܏ #�c͑�|GK���D���d��t��}' �b@/�_�*'Y7:�M{��ՠ�wg�S�����X<�@���"x���=�ő����b��D�cxB�92�W�Zi="FB�
]�W)ib�+m�c���j�Z�b�;���qzzU8V�#r6n\o�M�/~��>n(lY�5+�Z�Q��o���D�w��O wV?�_}P��`'���=5*�W��!�k޸���"�O�����f7���[����;��x��p�GV9��=���[��8(/�_�����9��}rR�͈���F���Q:�쳏�
'���&�AǦ+�̝
��PP�k~��˿�ԫU�&�=��#�8�|���[x5�^�{蔑P����I��� �ND�<��m��g�o��v�>(t��iS�d4z����8,�� �g�yV>*Je�a��AU�e�k��!0�̽�/��X�sZ��$sj�;�8į�s	���</JY�tUj���N�������.�J�[i\p����*�	\+�X	����' q�	X�x,.f��0�1���7�Y��N��<�䷞pg+�X����L���BH@��}��wcQ�B��k�U���F�����o��j[S�KG�wͰ��ܦ��x�q�O��ڑjG9r<<>�Ŋe) =Ѻ�"�ř�.�kq���?�c�o��#P�5L�C��}OŕP�E�#�W�.�[1Y)r3�����]/�UJ��\��a�u��pD*t�_�u��_�)�~�[*�[2��/!�?ױ�
��w�V�$ӭ���!�r�Q������ DJz�������3��RG��s�,� Q�c�A�E�K���5F��q���.���x���p�ܥ��w�E+�L��ᵩC��<������3��J������X�j�|\���rQ�o��v�>p����B�m���2�nf\����8v�`���4'�\�c�Z`�@J��X.;{��w�u���;nUi괔� ��,�t������oMhw^�\��T4Ŗ''k��!N��3-�V󅋊q\Y�RPhYd ���v3L�hȸU�a��?��9��1�:��H~��y^˩{�x8�\\�&{��%;�ٶ��Um�a�H�IK�7K^�b�R����0�M�as���ѳ��S\�99������([���c���ph�h^i�{C�S���e�q��B�9�v�x�y"��̼+oD��8�bu[��7��<\Ӡ�[��������ּU��z�u��{��y��kqw���+�n���m�5�C��U@�c�|S�a��=*��8׭7�V���IƁ�,��y|n<6CIr[�ǂ��y�q�]{�	��s.��šg̘�Z�N��=�s>��Ț�h���
�޸h�ʝP�c����=�桬V�8��c�=� 707�V��89�}�6�$�V��)`��.A�$���F�[�B!w����z��������v�z��m]���X�4�f��\Ծ���#\��M�:ϧ�W�\4� �-NW-t�B�nd���T\�����q6G��#['fN9��<�8��[�Z�����Nl��=O�T�rܞhe���?�r�5vt�j��<��\��R�e�IT�"@��.�ױh
���N+KZW�`����\-W;���쬔%��Zc���G@Z�syK8�{E|s��e��ik`-�
!����� �>���n�� �9r���7��ϵ5P�gn����-v�"���f�������^��w�s�Q޼�T��;�7UMT�\�TU��J^ �U�X`�����T8�68BJ����kTB	�H9���o�ַ�u�i�偁����qy���B������V�\)�n#Ak+��~H}�6�B�&1}��Pz*\�3��9��ŋ�A��MJ�C�v?��" ��鼳#�G��र�FW!����E�Z���U��l��ط���R�k]�p�G*�9V���!�v/PA�]���>wm����ⓛ��˶�ݤ��
��E^�,-t*>���GK�n�T������2G��U8�痫Q���/���Z���?�*+T�]�+��U@��k#7��Z�@$Y���a��U(F�T.u��o]�h�"ˊ23z���W<�c��Q3�2��@���M�����-:�O����Rr��wY�7�[���۹��Bױ�ρ}�^Y�[����������sF��z�fU���Y�[;�֮aŖ)v� r\��|W�ޥȺ�.(��� ���;Y`]b�~�ל�<����!������W��|��\�����3N8��?�J���={�����
�)�/Y��ͽvII���Æ7��������>81���y���]�\Uվ��f7�WR		���"Q�.��bA�
Ҕ"�?D:�	��@z�}������s�7swؐ&����y����)�9gmZ��('�M9�km���9s�C�\����z�4����b�E]����]ҧ��Aڻt�)M ��Z�	˄L��$1��4�59y�:���&�pa�H�&�Ɔl²�P9� �dX��ɇ�`�}e�JcS��l�����n!�q"�P&�H�V�u�ӥ��RѸ�&��� <"��뉬r���CK����] d��	��J,`$~����e"!,q�G)U�Q���
Y��
�����\m�[�i5��m',����Xy���B�`���m�G�;�~\�<���{~�����#,t��l����!lPW��FȌ�W}���O�:����|�n�S�Je�*XW�l��-3���Uȑ`��J��Ҙ>F�l��Vl�խ��w*A8��D��T
��o�~	�Y��ǡS��Pl����f��6�����ߡ���c��	�Sݫ:FG����*0����Ք�*�6��~��\�ێs�)P|�9�E��Қ�:�ܗ��F2!32����(Fq"+��s�c_ka%���1���s���w�	��΁m�|�e��[��}W�;�����P��/��C��:[���pڊ,>�X#J̟7�6ŀ�6	E�O�2�?Z'��{�6?�����J17xK�ba�@n�1A0�˶�6!2!�T������	5}�h���T�#��e����\��;�l@H�|��i�r�bIs� j1��ɂ �Ʃ�CV/S�Q��;��w��I�#��.�m��p�5�5 ��"�7��q�N�fM(�n�:�����X�\�tO\��Q��*n�ג	f���Yڒ�����~��C,%KVb`�񾔖����W�d����'��u�	ބ��#�[+���d�_T&�����4 d�}�G�%l�w�{���_8~3��ٝm���(e;;b2{��W�<�&�/���J��O�kMn�p��e���o:b��}��J@x�u�{��ݮX�|�6�`mG�����o�	+;vQ��4�h�*
���u��p�S�r){�<5@y�ϙ�/r��A-s=�\����0<�E�5l���/��A���k��o�����tͰ����kM�=H�lނm�k\_y�fΚ���N�����p�o1��MfΜ9���?�����R�f�|X���ǭרCp
�$m :����j'��X ���>Ս.6p��Ԃ���7˧��J#��ĵ-n��#͒���^y����@��grc��)�r�9�"��9�P	��[���d�SI"�w����*����6�+�%���<�1c�s�'>Xy��\\H�����yr}CC����k�լŔǦL�O�ʄ���%.���.�P�p
�\�n�B1l���Eٸ�]�W��������z���Νe��tP#Y��_�iAxoKG��?ɧ�#@n������ν&���ud��_�{M�@*sb����|=��zR�=��-�����
s����&@z��9��Ȝ�|�i��o���؋ ��O�=���c0_�L�����馛��=+���xɈ�|R�0�
��~�����2c���p��6/����y��Xt���%��b7q�!����tg-Z�U,����Z�����mAη,��C�����*���`�ߡ��\ϑ�\��&�����4qxL��4���^�u��<$Ņ�#y���O &σ�и����eTԫ\���!#Z瑂����M�fV2��v��g�g���,ؾ���\��=�
��g��Uq~j�Rt�
�46�;+�Ǘ���e��R�IU:�r"O��5]�|�ɱ�z��<�<$����Q�B����D�T6��ڥ��Kz�`g��V�����A���fU����Z���v1�k{�.�5-@��*��'U�]W��Ї�[W%cM�_�q���l�z�PN�!�Rs��d�xW:�*���b�9��K��O��j:(��^�PQ�r�TW=C���c4�=�1��d�v���_���?�ѳ�Zc�k�o��C���{��'L�>cW�2��I��o>�"7+u-�	�'�W��f�շ�aqw�'0�;e��1G}L/L��l�طz�$�0�jOҘys� I�ҾX�T7-��C�9au��do��b�QJZ��-h�� ���뢕�T�����@$���B��u�'��\���C9���PU�	�-��� �@+S .b�GB��5�{�(@{�h��� ^�d�$�T䂩X-�b96�g-n:�@X���12�Klp�_� )�������R��,�"q�</��p��N=ܞ���9���x^*<�������>n�*|R��Q�˪���|�>��7����Qyn��e���`��O�x�@ ���g�#�w�ctd�i�Z��s�@�� ݱ�tl���!�h�P��}�P�!�7�V�xJ����#�Q�CjXJ5!8�	�UlX�$�i�"ǂs���pU�e@h��<�Z��0���\q��G}��^p�ͷ��1�}˷���Y�f�r���hNi}�#�����!�7�q��p�o��,��2��|
���8�Ls��G�%��1EeaJC�è��o�%�5�c�oc2G� ^�+`H&,mcB�e���n�p!ص����I`^7�"�5iҤD��u��ul�/s�%�D����v�"�0 %Z�L���L+�Iy
-q�Ó=�S���c��) ��8��ۄ���W�l+������V &�{Ka�5H��R���T���%�Ǥ�ER#��`�}�����}�V�SH�c�[��R�d��}em�ZT~S5>��
5��ңGos����d�|7o�\�wyy����"���m��+��`�j���9����k�
��#���Y����ˑ�m����u;F�b-9kM�sػ��Z?�� ��R���,t�ER���(mQ`n�u=���SS2���u�6*��W�3�2��W�s�'v�����D��{�9����o�k���Q�����y�J��\�y��F ������,���O�<�ȣ�����A�IX�/P�����w}�B/oi3�c��o�}�l�L�tԯ��� g9q���qIֹg	'ў)L��}���Û&P�w�#`������~�Vm��+Uv8q[�u�RB�_H��ʊWl]�9+��\��a1�e�S�]Ь�ͷ�o���f�V	c]v���ňL��\�����>ߵ�t�^$�L)o���1֦�{���Ŕ�;�ѹ�������.Vl��i��䫣��0��RKY`m�`��6"���a>ݏ,�z$�ƛmSgϞ�r�1d�����-/���)%�	����Æ��XJl��7ց�7o�yIj,����5��N֬@�-�z%��ך��}��\�C+fM��u�8ø~�C��S-g��� �k�Bԋ��V�>�I�(.͹%��3^=$��$�y�MҳE��U�C�רp_��<+FB��U����!A��A��Q�Q:J�!�
��5c IKχ�mL_d����{��yl������Y�����n��{�m8֐!�|J[�s<����g�)ZR�e��Z�R�<�4��H���@_0oA� �d��l��Z�"Ml�/��~X�2��k��?�Eźe�
���٢�j� 0 Ȓ�gH�b�P��v�6o�'���2k��<�bxm��w��C�{ذa�F#@�x�U��b��(���Ii	��IE��Č50���0���Lp�UN+��[����9.fL�
=r/3����$��	��R�Z�;Y������7V����L��-<�Ee��\Ф����l����0��К������@`��tk��x5��pC�T삅ދ����us!&�m({a�ڄ���4vY���/\��nD�����nM���˾�)	���f'������B��<��k^|ʗր��{Ǘ뵟�#��`��!('���Jv}m�=T��;��;D�`?����~~j}���F����g�)*��c�>�La<Y�
�d�؈By�|������g�����8?��()C^'�7�o�E~*<ƴ�:dM��A.M�����:�gп��w4�R>|�{�+U��"(�]c�&K-�k_*��[Z�����j���t�z����:͘>c�ɓ�l��X�|�s̱�0�;���+�I*�Ih9��&!����Y���P����i�*{��m]vɼä�Y7g8�?Г��?�n:�*E�luVY�8#WA����y �]����! �9�Z��>�,�Ը�^�
�'��i59GiS���)\�kR�oZ�$�eeZ�J���o1�B1V��˜�������h�.f)s��
�B%�QR����K˩�%dѥ�[����y�Mg���'�����1%C;�{�7f�?*)�_�y�	�*���O΀*�1fN��A��刑ϛ7���O��,�@�#��u\��]
��ɕ^�n)��-�@�Y��uDe��*��{̹r��ʱ��n��<�%<4Z�����z�|�W�K��a�rLz�i�s��<T̞-=ÜK"ˍ9�g�yƥ;��;�^{��qZlc8h��m��q&�˱�Э7�B�/����T5N�����m�vQ��.ᢷ�z�;h���S���I'����E tq| K�V,+I��@P`�t�{�[1�[���a\\����qm,A��PزB�+���?�&�Q�뼲ȵh�l�*kt��;�;����]>lU�-r]{�5����}/��8E.ӽ��@rW�V�3�mT)MJ ]xZ<C�FhI11/�n�f���G*
,���`�<�z�"$��V*= ���Q�������c�Ә���'ŻSYd��1#��.�\�E/�B2�7 M��Ѝ�2�d�8��M,�#��������1�kt��B���X.zU5���n��s��`�y.��<����(�I�眶I���X�³�9�祽����1<�y\ ��h
X�ߙ�'P���5�g��'<a�>���4�I��g��j�W� �}m����^�3V9�hި�����m�T���h�>��<���x��sX$�]w���7�����޵����H ܥ�0�����ʗ0&̓x�I����&k;�W�,c���;��6ĵ-I�?��7�+�ű�m�J-�lňC�[��=p-g-�r��Z�@�n�L�Z�IK;������B���yS������r����p��x>=�r�i�����
ᘴ r.&\ T&RJS]��7����=|�뭴.\x�m�:J��x�/�%*��q{��Jot�c��'=b�h2��>�@,+�!=4Q�	e�y.�t���ϷujC�w.\�zvF��dTT:Sr��ґt~���a����䜣�JV}�n��}���P.Tl���S&���Q���55,�I��c�x�B0׼A.�����T�,�gB�dG���ҩ�D�r���1
�|�+l�TWyo�g��W�%T��$k������뗵-ņ�����8%uqTB��i�c�=Y����!�K���Kʆ]'��H9�:�3"�����q*�DeC�+'����/?���w����%��K ���0V�<�H0Z�S@S���&���k����.��y�C�}��O>��]��N �jY��eɻ��҃j�H	B��,a��x���҃��
<�W��	��Xa7�6�n���xR𕢴x�h��dF��`�Z�^.4!g r�%�Ԑ�i���>b��<r���O��q�T��
s��1Ѣ�1�p.LZt�pȊaܝ��⨖�9�a���uؙ��<��!�Л=aL��R�R�*�K�.kyw�$����-+;�,f�'���*H�g^7���p8GC�"�M���;ݥ�g^D��x�,�.y�|z~�K�o����$G��Y�ӧ��>�T�i���d��T׿�Cr�
��Sf����u*��9mo�	�M��Ϛ�~��j<�M�FYI���U�V��(��yķ徲�5V)������6"�I~�������BeA�!��95����zF�oݧ���U��h���8A	��Hy�h�ki����t�����O��g�n�<�k}J ����y<2��7�����?�pt�9�>����|,�Nd�����:'�Yd��-	� 63b��~��)$-|c:�S����5���1I-Q��;+���0���k%k[�ݖ��S��P�U:�S<��;��KJ:�X�o[��	j쐥#&2�#Vl �R��e���p�P�A�,m�E���%�\����Ʊ�E���R��p_Ń�^��<���M�	�9�LZˣ&�<V4���b���u�b���ۋ��n<7�i!ӵNE�dY�t� ǲ��u^`���@oS�"	x�mFM] �*���(�)0}�4?��ұsG���DX*_��g�LT�2����ȝ�����Gw;��+�@yw�\н�5s�����	�
:CLU�bcIe�BpN��:༧l?s��\�|�ȖVN?�tY�LT}|>��8��dZ�O9�$i��׸���A���^�W�q;&�w|�{�G�VS<�)T����|NX'?�%d���ىX��S'9��<����ea+^W�%�m��pnJ��5r�V�"x��j	��!����h�JC��x"��j]�'Zq�Ă�М y��>���c�/Sq�"fH����??��{�w��j�^��:K`�&?�<n�}�n�6/�5�9Tv�6V�P��9�����׿?�"��Z���rEY�;o�s��}�B����?C<(��Q-\���-E� K��󂛰`�֜ [�j^W[�Z
@���c�a��gsr�C���E�	�5��	�\*x��].D�r	fLC�KU�R�𔣡�g'���\\X B]�Nl�b����,+2t]B�x��e����ո/��z�"Qomt��/p�E��R ���D�t,�t���:��b�W�Ȇ��US����F�'�֪ ���a%��s!�<�RQT�E�S���2K `0�GLz*�E���q�M ^��&˗-c�c-v#%1W
h+@Y/n��P���M��͌S�x&-.�ۚ^�)��i�w�^��%���`̜�o%� Ζ�L1��Ă3r���?.�����0�*P�5iyψ�s�Z�U^TV�<�3ܟ`.�Q����C�4���TR�v���T�IֵB;
�x��!���u~�c�����,$�+TF�њ���J�h�\�Cc�h�yj�B�5$Uiֳ�O���+Εp=L<�Hk�1e���Q�7�ԛBA����9�r�(%�]`�}��g' y&*-"���E]t2<m���:,�.]:/�ܗa����Kv^c�"ü6O}"�[V�� iF#�}kKzΪU���ü
�,,y��/�췗��o'�ܴ��k��irs҆�';�`����9tm�.:����ԋNZ�Q�Z�oI�6��=B�n�� ���\�eJ�2�`B��/�pe#6ʉ@���K�,]�Q��\�ZP��;�_p%��-�s��R�G�&T:#瘹�� p0��hѤ�CkA�T�~ҒÂ�6���L��*�ѭL0�}�uO�4טi$?��pW�U�H�[�]�/O�<��3p�"������Qܞ�'�r��ef�����H<S��D:g]����9//���K��=�e�c�1��V�<�۷�����s��yYJW�Ԋ����8�J�x��T�A�
u��y�?M�)���uo,�c�ƍ��z�t�^+�O�2OLj^;�Uѝ0�(�V���p��<xR0d�R�4:����WE󖼀RdQ�[��x�x�x_xr�����$�Py�iSσ���k�wZ��[eB@:p&�ۼ��^��A�1Ւ2\�fE�m��߯��y�[�⭾��z��[W�^�[�./��79X+�'O��ٛ�ǟv����nj����Z��(Bwo��������!k�N��a<I���������x��DE�?0���ơ�%�LY2�7�@�\a�OsaS!�hd?j��v���E�������@�.�a�e�� 4IⓌ��K�2�XB׺�\��I����-F��y-jdbnO(٨��1�*�]�I��d��䯁2�¸����<+;î�b嫠Ȱ�ru�ɁB����&�t��9|�o�)	*z#�\2�e��o�E����x�rS*�׳��>�Z�y}Z8=���.:��/?����<2T�T�V$7)�����>�Y3�Yj��g�.q|�5�yʚr�<�R}xyudIx�@�H���F�q;)ߡ�+���#��(��۞�ȥ�1q_�+U�6�1g���
��%�>�&h3̢mD�q*�X�c @ῐ���H}F��qw\�_$�o�v�0�	��~��k���*
�h-	�`!7�v�3�
�R�ۤ>債�g����O���v���w�QGy�}��	�Y6k��oT�H�k/�F#<�z��y��.�g�~����l,(�8���q���E��tG�y�U�tc�����'/"�p�G~����C7�P%Ţ��?4�d~m!+PlkO`�{�y�-*C�q��MZ�h�,�B]���X~�K�*���S�����x|Y�Tk�EQ4f-�i}�r]7��Ozq��	��P\N2�k Q��p�2�
��(+���N�8AOy�N(썰<9&��mx���1q�#���e�8�ʌ�qgܧNx��.Eû���d*�C�6*4a����y)p�X�ǰ>쐟u�B�tz�B���!�sN0ݐcP�vze3��c �<5�+Lɐ��1sq	BK\`*+����O9ȵ- ��턒T�|I��9ON�t�X���(k_s�8xK)
�k�͉��=��^�4�����i0z�ʜ��C�vR�4/�M���Α��ȋ!����yj�V�3��bEZ��)pϑ�/D!����"�����"�1�Ő��\��so��=F�5��@!�m�K �|u�~w+&�ZΙp��Ev���3�>��7�������8�O!Q����jO������-�h-&z�l�h��$����탘ܞ��@����k$��-��ܕ�"�E��D�HZ>?	J~ra�ƅ��	��EU�h���/PI6zI�7ݸ�����)J�d�"�τ�p����)�4zZ�Z��\7� *_+�,9��]��|�]�l8 �E.m5T!(��G�+� J�60 ��r��i�(�ȬP�w/D�\���9Y����t�K��5΢5��sL|��]c�/�"�H[�}�|�ׁ�Va�W��I�<�\Q�nzA�9IxA��y���n5�<^}����4z&��,���_ d�9& 	�-.��f� ]cL>_�Կ�2��X�hyD/)󩠦��I�+����q�ܶ�v�k��e�� =U��O���lx��"������k�㉽>���������6�o���}q��m��g܆(�D9i�I~��
���ɢK��*��ջ����w���l2�����%K����B%_Cc�=�/"�y*��R��_�:Y��<��9����P���4B��O"�{p�&+3��$Ӱ�NN~j�ުԻ%b��
5@@�?�Im��F��t���Nd�����ֈ��\b_ӝ���|���a^�&�˿X�\�x�QQQ� ��Z�f�66g�ܝt[���)��y��%Q|ۻK9��\�����.��I�������M�=CvuT��Ð�ʨ&�;��E)KH
��	�k*��΅�����&�.����$�����x<��L�^��$Y塚��n����%��MORղ�+@�h21 WC��#wr���>p܌���oD�4c��y��Zo�|����9��`�W����P1��B��,�������Di*R�PF��f�ŎqdQA@�3���rk�¼��-���Y�,�˜�"�H�CA����,[�Ԭq6ѡ�g�x{�`����'KV:O�������*�� H�H"GDR]�$v����XC�c��.;�D!#\���`��CF�s�CLv��vm��P�/#@�gv�1أ�zb\m8�~��9���~f���	��p��s/�(r�'d�*1�����x7�]s�r�sGEZ��}���J���Be��K�����=��K��w�n���v�� ��H��Ů������pk|
>o��g�z��W_y�j6ݪ� �   IDAT��\5���Iҭ�� ]ϴv���#����f�"8�ڪ�;�Ӄ��0'�������� �EZ�liQ�������CjcZUֲ��'�P�Pk!��:�1nǅ�7���z��"!��o.Ы��2����f�F�ģ�,nc��	��p(��[�v�pAD -��N^?����q k�4��i`|�Bo�4��� `����XT�V�R���щHfPZ�9�9~�B����K��)]�X�Je��3�;/�_c�c����$rK�"n��d�Ll W9���k�,��B!�:�h#�T��f��1
�Pq��g��yտ��)�s�V�ע��4���ZW_m�o�Fmn%{�`F��3*��S@%���G���z�䑰� R����6�g�� B��@�M�6qf*�ɕG�±5�SLz��f��ʹ��$J����Z0���Y��(a�F�$��K}�n��х���C���s&���D
RB�Dĵ�����A����'I�|�7�|���'��v�<R���G5BD�/L֔�)�2ٴ�~��v�����?��뎿�r%���
)�z&����f������)�e�s1�C�>}��n����xbT�A-��s�)ġ-5	�PZჩ��xÐ��n�v�f��e5�=�	������Fr�KO��y�p�
�
-��H���kT̗֞r�uN�~ηԬ���s*(�z=�yP��rs���d��PNTV��\�^nG ��G�u6F
���^˖�����ѭ�Ŗ��W���`[XXl
-Lz'|��VS2��9K�Y�G��� *[ih*$�qʵ�{aJcT8��I��3�z-;5�ɷC-�r����\��T���η:�����Od@��ר#<>�QnvYjJ�3^ ���!�oR.y]M�fO �� �C������򦂴��������X���p�b'��꾩��s$=f3$7�o�e.o���5�p�3���Ŷ��y���H8m�I�|��J(=�<�(�ۯ�o?�>��d&�kc��%3m+�Ƕ�Eָ�Ƃ���$+��c����?��u'��;;2�x�/q�M&��pJ�!S�[[�w@��'���V@M�	lXu�ȄV��ED@"w_H�
��^��X��&]_T\�I���i%����|�v��ޒA����!�֬�S�
�c�� �sҲciR����"kV�A=p�n5>-&��~f�{w��:����k�r���6-�Byt}+='|��\>\0�:�\46~�ء�`E?Lic����ڹ�L��	f��i������+V�U�_�5��"��~���̽'&��6l�����N'�2{@)`���^�p��8�
�R-G	�-��s<ʝ籨����>Ԋ�{%γ�)W��YW�R�0Nn[	���:�X�o(/�c��2����s{kDX���r˧Z��3P%@(�����2�c�z��W��B�v Jݦ��7�6�]�nCYi��h}�k��밡����������7e:"ˉ�IE��ס�=�|���f�E�0��=���Ϋ���T�����:�I��z��2�y\s��?y�h�Zc��Z-�	}���߾�n4�%��-w�@#|d%��S��A�v�#�Ң`
Bd�˵)�N�� �-�LnU��j�7Ԡ�i{)Z����H��b# �D�҃*�߻U����M6t�"�M��ԅ�	uX�"$@׿�x�"W�����w�3��J�B�R�{�'�vƑi���ش��p,���M��� �� �p���N���)�X4���%�c�Um���R҂�5�{���a�\)d�׆�;Za�PM*X��T��P1�^o	�N@�<���{u�Rn����})��q�lq*
?�,Yjc���nw*��m��8��k���V�P��V,}+T��9�<�W����`�0"I�
��P�oo{)��X,tb�Z��NUd4�Be�=������nV���T�a{�	��2�m�_õ%\��}�����5�&���]PF8��e�BFZ�ß9��Ӯ�k�=_��濬mjĿ� ��F����^��B6R�Fz��&��П}��K�7�Š�J&[��r�����~`i��ׅ&��QI�ZZq\�,��LBH�L]C�\����}��MP�uвd���*X��+W/�b��������";��Ilc���GK"\=Ȋ��5�P1��h	t����1�t�$Ĵ�ض�[��$Q��7�3o99y��)��+eK���D��0N�X�KĶ"�@�	 UY�<�G���S��YK�z�?6?��N��
�K���I.$я��ۊ� �9.����`G��&%��ĺw�唝�k����kQ�jy�8v��J��� �Xlb�@��t����=�YTTlY�cWP9��ܞ
�BZ!�Z|Z�4�C�Q���p]ӱ4�R�<~/o�����54�8~)GkZG�x�"�߇+���Ὰ.�+�זz�(���
 �v�:`��w���ƃm{�n���5C�K��s�'<'|q�h>��Z�tLT{{���<���y�/���uT���&���B�s��;4Z�8�"+�O�5��
�舶=i��M��G�b�.b-�<�g2r=Pb�d�[�k�PKլ"���κ�������s���<|h%�Py079.Դ�PZHJ�2�n�Е��֞r�&��P'`�\��>#���I�+;�Kx�t�p���	��t=�t3�y�.��T��,�U5��]L�}t��F�����&<��X�޹��~�y��ܹsMv$�Q)�B�*�����ǣ���p�b�sp�^�$��G�L�{�`ޙ����b�$V���9S�X�������
�7�o�إP˙�~#�Ee\Yh�xZ�<6�,��'���{B��ջJ��a�rG��d�����{<g���g��/$Sk��9(�d��|�����d�� �����2�J��6�*1���Ǉ�ϔ�Am#�<��1�;ck�)W$[z�w�Փ��+���1�]_(��8�K�Eb=��q�Z�kZ<%_�{�BA݀8�/��tD�!�Y���R��бg�8$�:�����3ϼ�'�x����gMC���H$��/[��!��F��<?��R0�8��ܠ���D��!�������� ���5#�3�F3Ұ |���8����8`V���Q�%E�i���TNh2PM�a�K��DY|��hq��#�'Zf���
 \+N���
�b�dX�Z��o\H��ւ��,.��VpO1��"��2�xY!1-a�XV�����Eθ�ʅ�T�zV:���8M.
�8���c" qL�<gT�C��
�ߣg��2F��miA���r��?g�Y�${Y���]����� �-��g�q\��۳:S������5�h���r�y�M!sg�>-\~��~����ˠX�t0��w�\㬭n�@$�D��J��X�q�5�9�ٕ���X<���!��#~b -�� �(�����*�-]��η����\�<e�6>��!��0��7�-d'�W����6�g��8�C����:�$Bl����aN�E0��ڳz}K�(5����h������dF��&��ga�+՝/�U��4�Ȉr�Se�j�o{�N���*�kr��Z���-�zV9_|�:?�BO��U1C1r��3fZ�H�/9���o�я~t<cklұ��X<�HHs.�����%��s���+̊�c�<_��s-t4��#��h� � �C���9��ZX�Pq�a����n�Z�Z�{׮���-׃ƞ�x聉���ØX�x�@�B���]�E��Т�5I�������D"Ϛփ�x(��^ �*lƾ��jJ��L�	e�]�`�t���5^�9�E@�7-S�����Y�>$Ђ�$zyo�'�_��т���bfJ�H`dœ�]X\d�9#'fUU��oҬ���W�6��u�<n�$��x���P�=�_���ɢ����!��Z�q��F���z�ʡh(�ͅ�@$*Ɠ��ﵔ�3�"Rf�����<����O�S�T(���2�Kڀ ��{�ߨd��yOӽlϥ>�m-뵯��V���T���-O?���)[�^��}X�T�k<Zs4���W� 知ZF{Ή���$��8!�՟*�p�U�k"�Ǹ��Sm��(��.y�V��x����r<
M�[���p�������g_�
�e\p��op��F#xI;	SBc���| =W�F�}����^��r��Y4��$g衵��u0O�iY޲3WT�z�����>�Ʌ�7��2�H"
��&P\��;N8�#L�X>�z����;3"?	�������bfV8*w%��(�a�5*��e!Hf�VD⡆&+\��ŠUJ�T}��r�i�+Sa�D�<�h���
ֻxF�WI���I9�t�<Ğ�uϛ;ǈ��<�*������wx�~�d5��ʕr���A
�<%J���dnx�΂0�Fؕ�f�	9��50����B�C*T	�Ʊdf�1 �(Qq �r_���|�s�^Ѓ���K��%��36�=F<=B� �;<�*~QN��ZR-V=��g�K9N�&T(���DʵƩ{.@�}�rx�6� �V
�m[&>�JUPϻ)��z�w��W�X��F��tP�T逡��m�~+���疟��7�������^�����q��h=��g돿4��������~�a�����o�᳂����%���(�*��5���b�M�O3������\@Ǣ9�ǉ|�>wts�у���gһvQ�>�ފ���â�\j�/.�f�\r�s�!��/Z��^1J>0z����w&���
�B�a\�����\�e!�8ҾE~R�g-8q��-vŗ�Y�B z�E<�[=�p1�ߡ���,�T�c�|	d�g�z�x}�G%C�Zx�z�L�}X���+I����Q޳G/c��yn-B���,�4��c`�x���`Vh�^��܈�x����ck��4����]Ǜׯ�wuu����+�k���ܣ�"�ue�f�����R��^�P���z8.V�ޣ�y/�ܗ����T�'�Mh�j������b��g�LS-�ĳ��xs�����?�_�N�y�L
�m��)0jOQ�=m���?�E�ZEF��{�s�
G���^�$h���Z����n}R.��!�Л�{��`�QV�A��׸�]���/����!fRd4���r�=p�������e��z��x��K`��)Ň~�]�bm��d�6�j^��)�ku0���?�7��SO>e!:Dܗu��j���=�r�%�D�@�gqM~i���n��}.rr�񁣅/&�*��$����s���6�e�W��kh��r�G9�^+�HPѧ?�l�P['#5t�����<u�	��u�CkH9�W*0a�ɐ5+欈�r��5xXH��	�X�\�x.攳7��H1འ�)hK�,���(��x4�����<����Q�<?�_�����m�I`S*Z'X���<-4�e��
4�\�U E� =�W�$�K��t��;�$������mJ�{OK����L��5{��D*է��g<>������$X�����~M���,�p΅���"�j��i�T�׿�0i?�%�j;�$��>!����<��2!�J�� �j5�@I��7��R��:���H	�3f�gO=�?��.�>��#�2�xۍT����̹�����hqA�kN��E�4b,��7�|�Ə!A"a�{=�	M��K��ݗ������©Œ���A}�Y2�e�őYR�|���N ��ʺ*ߙ1	��^�`A"%J��c��0�Z��N���I�'�n_�6D�iE���S�jc�D�u{z��)���*����)˟�@�䙐�O�d�{A�:��&�����`w2�E�±�Zgܗ����=�O���9�tW����DC}v`cݻ��CMSnr��A$��y����*{� .���Ǽw�wx^����ιA�F551�%'��`y��>�E*��єtI�e���F5�⸟ʾ��I�9��,X���2#��:)���\��ʯ<A����Ώ�9�>H��z���=k��
--6������m^����7d�-�����R= �.jV\�_w���y�d�y��1p�\_2�M`�����������c�';�п��ٜ{���N��5���IS�j���k�.���'�h����F��������)�C=��	&|��(O�@�L6舊>����V��#�g��P����X��tV�B��",v͈}e���F!��U��p�҅����4�D,MD��V%�6�ki���?t���S
Ֆ/sk!�1����t�\���=��KaЍHZ�m��[�O���C۴޼.�=��4.����f�|��o���]�w=X�"�����>N�]�ۦbDVv' X��/;޲�Yk�����f��ڴ&tSG�<X<�&�d��h��b�y��,���nOj��G���Er\'�#ҭ[#�e0��&��I@��U��]�a�q�%��Lk��&��A�̺�T\���V�W�Q�6֭���|ҽΘ9��G-P�&<�j����|b����<��1�I���]Q�������|y//-@)Z�d��V��#t��g������wλ	SA\ʾ<�xބ�R�=	�lN�-�6Vs$�� :\�S-m���E��
� n��HƗqZ٭ �r�"�r��Q��g"�7P��w���Ƅ'�i{?�ҫ��:J��|��?�ʫ/����үT����M�;�s��|s��FwHK���~<��Q>O���F��G��������ϟ�Zkz�>�[�������O��f�R�1����_��6��ϴ4�u}�f�]�Brar�ZXx�sr�s�NV��� >`�t�~*�Ab�*{�-)W�%KP1q��Çσ�g|s_.�tՆ1r���قx��9ts*.��8i�������G� �ň�T�O�{��n�;�O�#�ZG|�*z+Y}�	�M�	y����'-I�L�Yt�@@�*�yɢ�|�J�?5�sC�@(�Y�m^-Y��$ǚ�`���˃m92�;w1��
���\V�c|��,s�z���zPL���d�#+�"�A��G�����`.7�x�yo5��c$���!��a��[�y�&�c�Z}Z��{>���������5�R?S�R�z�t/R-��,�Pa`��tMR RC�Q؎+�Z���E��	�?oq�	׫PA�t�h�B�q�^ɤ�M%ܟ��b�dy�ʬ��+�l�.���߃>��Q�6���c��m����K`�yC�Ʃ��2
B�8��z#I2ݣG��k�Z�8��cn���?}���Ϯ����	�M�2%�	�� _㋥��U<��N�����a
�fSm�e(0O��J�%,~ꁖ��q{�.����er͆.�tx��$X�d-zm���-t��	�m���+�9�#[�����U�k��bx#�o�%�T����w��-���Z!A��D0C��ɢ=M�� �2vǃ��i��b��]|�7��>�>
��EN���2�X�#���p� ��t���҂<Y�Pg�g���A��2$�G��@!)4�滳�:�0�B�~�z�
����ὢ�E˜J ����XH�!�8��q���h��x{��g���Y!x���^�@@$�M�0����yB��<(�&|D~���gL���B����z�'���k[��{�B ��kX��O�"P�C���<	I�~�|���A�Xs{(΋v�q��v�q��n����<��g�r_|aG/%��k.�e�kj�j�[\'=g	,�ґ� -@ :�!:2~�6Qt�y�s�;��믽����?81�RN^,r��Y���OWoC�;���b������>�oZ�b��B��!��$Aha��o����Z��@YB�>���{���D
Y)R��\���d>m��Z�x�/,�����u��V|�����x.�h�z�����P&_��e�;��b�>��݊<��y�N`U?r�{��p�*X�L?��Eഘ1��R�B�E��rlZ@5v�T秔�P!�����P�U��1rϚ��� N�]��K���2�+] � R�Wn���&/<�`�X��7��-e.�Wj���t�/�UN�r�></�k�S~�B&�0k�I	�Ly4w�<gh������g�B.���?|fB�8����-0���jc�3& I�3���0<f*pk;�3�� ;]�!)V�o��h�
�V�~U.��P�0�q���]>z��7����>x��ݏ9�x�M^WQ��$0yҴ�:��o4��0�?a��E)�~��"4���wu�����M$t������y�M��~��E?[��?�%���TW�D]��C�4+/Vɲ�. !��̚��n�V��Jd�x�J2ӵ �ҨC�Cc�;և�lBk(�>R�noqH]���\xR:

���b<�*^��'EŻ��+,*0���DY1v̺��|�-lJ@�Z}BFj3�y�.�mB)=����c!���i�3<�һv?"�x�r�ET��q�;~҂%����R10���/�|iGa� ��T-V�a��Up��X��,�&�~E]�6^h�*�
�R� R�`���1W�}P�BL}����{GSdӽN%h��1O���􍌙�����z�+Rj�9����E=��kO�����:>k[P>�w��\XX.����k�W?O���t,~�"x5��|����B
�z��k"��*��\�1QۧO���{���[n��fkx��E\�� 	̘1k\F.-t� �'���L��*0r,�v��_f��wi��6����`����x�֛�zѸq�  o
�Tn҆h�	����Œ�S���������S���d.�/]X�R�w�Z���������1em����c��.X���B?��@���v%�)��N��ڶ�x�Q �O�u-����=."T�jAlAFAh��zrPל$�Mk��]��g���p�r���\Wz���o�`�@V��L���c�9|t�+l ����q�+db�k MUŢe�kT����*�\���"%S���l(�<�#R �Iy�Y�×eս��C
��.�����"�c0~�7��^.����N���Xh)��>��i)�]�R��*D�����=�Vx�=��s���c]O�Z%��*�}��k?K�"zVֶ�P�eE��F����ε�z�#>B�ҧ��g�G���d�/>箻�Ok;e���HӧOùCo�����$<QQ[|�'����P��ssй�:�Nv���~ʤ)����˧>���W.�u��S�R�0�N6K�e:-~�`ltoa2��F�Ⱥ�1n�w���4�����G,t���

k��T���}�-��x8Y��[ ͘���a<����q-��Oڿ�����ߎ��[��x<ʀV2s��^�F$��x1n�K!�i�1������� ������!��^6��|E.|�+?�9�|e�����qXZǱrK����!vo�#�'>�.�eVxc�6;,k�'Z�+p�Q�t�� ���(��Qd�� ̻w�n��}bz]<�|��"�����a
���#M���ʿS-0Y��(��.Bt���Ҳő�Ck��6�<�M+��#�`��Rq��xd�.F�V9�|5����-Q�����@�˳��D$L��'��2d�1d/뤕*�B
���R�t_֤\ʝ'��|�Mnp)7�Fqq��=�^ǐ�S�����~\��a��Ķ.�>��C<H��uݡ�
��l���c/���L��oQ��z(Ƴ��	☓Ǝ;~����=pЀ�G{0N�w,�6�4q�X�8�T�K��樗�0KϢ�[#K�����޽�~nw��:w��ϫ��*�%<?iiE�x����S�V���%R@,��<f�cü�( ���uߠC��~Zɲ�,�-�y����� ]�Q�YH�H+�ށT����$[��@��z���EY0E�'�����]�'��7ךW@V
�"'q�ax"2��8M	�}0Yњ���|xn*U��દ5��f<�@�HM3���rArܡ�Q�^�$g�SZ���{oS�" �)����������r�Q����6�w�2�޴��wW9<�@���c��5�¡�3�@ब��+���L�u�/���㚲˜u�w��g�jփ�F+�x��0� g�� -���Ώ���|�8x3�\�^�R؊��5��nG��T�<��G���£Ҷ���yf�,%�5��������bc2�΀��ţ�d�crPT�o/�=�M�t�8��q��~!E�ׅ�j���hK:}�M7�0jԨ�����8:"�x�X		L�:m��<�\S��Л*޶ΛR��� ��vD�_����n����o�B0�4Z�uu���.����ЊeqcG��d�6�:�d�'�Xo��\l��d0+�9� �,�׃� &�h4�T@׶�U����R���Nng�i鼼�j��GK�,�d����n@�`����2��uXwH�R��ʾ*M/A�%Q�\Ѣ���H(�����D��R-��c�H��bϨ"��m��.g���k˨��ߧ �e�US��P��*� C0"�%��w)Y���h8v���ɝ�{�sܔ:��3Z�T0E���mYVW�aC���9��ҐGd�o���>��7%�ö�W������x�ߑ;�fM��c)K�-�S�^a(�c��OU
�lK�5$�QJ�8S�0�̆
��Ջ��\���6@�	�!��ϑ��P��n��o���
i�	 _�ꫯ�����c	�����'v>���ȱ5D7�j��u]�o>Cɰ+��h:tBGĻ΀�֢�O=�ԕ��wߩx0�i)YIK��|@岵�����򱨳�9c.�!���i!݌r1Z~zkA��,&���P�N��/,X�;=\�SA9����=���ʓ���k"���fއ(��c(voV(���B5�H����$�RP�^��	��]s_�Ϊi$'�+Ii���Q����J��H>�|���[��;>�eII�c��$p�)s�G�7uF���1Ѣ]�~�d��e�A�{$�H(��&8���C�����z��0�!t�S�uy7�T_^�J�r(E��5ʅ���
�R]��C(叞�,�"����R�D���c꾄�W����~/Poo|>��Re"��c�3@Y��q��i�w)&����N�$�K��}{e�_ɉ�-?�D���!K׵���iyã8wȐ!�0sذM>��u���JG��x�X�����>kYI#�v��e ��s"��<Wv�#,4��S�.�?�g�ã�6����5uʔ��_+v0�o�B�Cf.hPT$F�8A����A��`���݂�sZ����1	R���q?��t�T"㷩��Ӟ�.���}�*8�˔է�r�V/�O4KѢb�$"�>p��e3BЪ
�/�
�zmۍ�LŔ�����1�Rd%>ZY����+ras[ɡ=�K�^��*�Z��'A��q�CS�@�p2r?������V.�p劥�r��s�yE�Rv���^�w��&�Y�C
�ѭ+b�]�zt|+�2n^La�.v�<yn���M���kb�9Z��U,u|!H�
��%)��"��tHA����C6��*�:���\�k{�C��ۆ�]��!O��}�#�7��&����'qUU����s�7���u�n�O��)*�}
���5k����X�K�?���*�ۥ������k<^��k�|�owd\��w�}������\�T�C${B{KһѴ`q� �Wm��f<-nw-��b�.u :��t.����B������^���oa�'b��J��p����&�_�"kF�T�s�t_�C����k	�}�"��ބԛLk�euŀ����"s�9.��,I�z�ߖ;Y��L��§ɡ��! �b��)J5RkV����"-Yq_cn��ݓ��<���^c�^gH�� zR(�*��D�D�2�G����������.)��8
b�lSh�l
;�����}܇��9�`�\5xG���+iI�`�Ѕ�qsV�.J�Ksxf��k�����"9�B�w�=��Y�!(��O{�HxZx¹����)h܁��� =yL֘��ܫZ̳*��j<՘�K����� �,f!���W��x��=`@���ۡ��#kd�M,�u�����9��il�p�g+Z������|�Т3�bEXo�����#��0��9��=���S�*Yt����f\��l�s��l	' b��B��.J��wY����� 7G$-v�2:>ٲ����Z�H��x/��G�j�X���J�Y�9�zY�f!a1�ŝ�k����'k�
�{�eR��fűB7]�8\��lnި���@�H��c�i����CЍu���uzH���UO��*��im�X�k�����K.$&���#"�)Fn�Z#�j�$�$�߳}�#��kI	��_W��a��`�/^4����P>ؼ��+:@'���=�������k����+��ҧ"$ֹ� gE���9�]����j@�<z'D44���]�
K\�^��=�F��G��U�ղ,,���g��3fD9���y�O�_�S�9.�cz��1�����Ʈ�+(��<��?��!�>!�h^�ӟ�9��mv���y��G1��7̏K_ڣ��HX ���|�u���]��7�C�}�9J�x@Okg��VmQQq�9��BU����=z�X��� ���X�0ȲA���B�/b	ldx�ͷ�����hYM�%=DhT�$��ŉZ�?� �Y��_��г��rᡏ_x�����|pR��|�2掳�g�Ҋ��GV����ć��rF:��0�&��+!�Ȁ�_n��}!�������ޚ%���%�7�r뿞�P��oR5jH\	-��D>4�1�:z�	�'A�c7�r�/�'7�-��A 1�9~^�Y���,���0���d��g��xoET%��'[��~nI��z�Ar�FN]���fut��!�]NV0������G���/�,8*o�U%���ŋ�����`�/5=��k��w�P��=��ǩ	�2	��ͩ�H�S�߼<c���p�)~��_)�/?�>�S`)�%��[�ܔ(�8w~^��2e�'�D
�����)��q�a.��ʐh9V-�SI�KE���!�3�7�:�O��/Ɇ��Z��q���>p5�C\�)d�9О5����܈�˟�\��q+�
�1��:�H��ٻ�B �
xB�	�L(]��W@��ߟ�E*q����x�7��?^�����8��K_\�i�C��K��Lw����:�wd�2ӧ�� aZ8-�0{�=Z`�B�K���/�/Zh��[.f�NqQ"��ר)}+�	&�,y��k���^���[S�P�B��LP"�Ks۞֫Rμ�l�(�h�f�dZx��x�չ�e��$����E��[Ț�1}���J?[�M.Y����­z�*-*��[�^�H��{.��ib_���V�23�9b�� fZ� Q��9t�-l�B7��m�R�8����<J�j����,��`/�)S`�s����|�vT��ֽ�Y�����Ў��dar~L�:5�N��=�1���V��R� ��ٌu.�����eHSH'Tn��\����mR�R�;]s^ʀ澗MN�W��V��u�m�F-��O���U��|㾯�wUx.V�{lS�j1���Xu�{t�����q��7F������(=g!I�/\�Kωb<ݔ�d]t8_�C��`����_~Eg�3��D������ �� �&Y�f%�٠��@FV��"��i����.Z�l!ȴ��']��&��F�]�ooM����c#K֫������[�+��'�c��cp+k!���3�]��AZ�mA��C�HJ��+Hr�Gd7Z��5�^�C��Z��I��߿��@Į��}�	Zs$�y�.'�!t�x3�N�23F3���4���u̇|v��U?�@.e#U)KIsG�]E����c��?�ʓ){�XD1y�88o��9<w߾���\tq�D=��1�J�-eK�~ҤIв}D
��XsL2�}�v�\T-T�e��� 
��\C#��c�:�jݏ�-��	��Ɏ�5�>��w~���8F3�I5?q��ixk�{���'H�p{�5���F�w�]OBKI�_�6~��%�V	��އ=�>��!2C�Q���>�,+���HN-���֓Ft��jk;aq�S�p<�Y��x]��D��rf�n���2�1fZ�Q%0�CY�<A��r�͒��K4�{%�֭�;�mvltl�ضmwl��`Ŷm۶�ܽ���_�5�w�z�
�&m���Q��D��a�tS驎VCSyˑ��G����}^5�V����4@��d���˃��:��d��>0�68�8&�ht�N
�J� ���?����&���5���R���z��_�G$f�a���ە&#I}�@Z�}�ÙZ��X�!���=������o8U�@��"�`���b��o�2t!E��Xo����*�h����y3~��5-`4���N p�\΀'��񼧄U�81�
��D$TZ����������'ٽN�ֿ��t�rb�T���c��(j1��:��c=7;my����'\�� �1ܬ�g����A7�Z�Z�H�w��h�����?58}{��.����g"��t�*eS�s@�"��CE�!�l��[��>;�1�I�]s"�g�����E�7���H"�w�9P�,�Ĭa���1i(���zےy�}�ʒ���ܣ� ��*d�yt��e�dƹ-�������X�
`�>�g����̽شfN�k����z
Z��ǝ rςDid[�\����x)R�*t��^[�]T~��}��,t%��*�������z�u�0�ݖ����F�Ftgu&�Bh��	��Kw�#�#6���x­��v?Y.{�/�C�|d�C��g
D�
��c3� ���vu0�T�����J���(�iV�z�����K�3l~3�?6}���Vw�.��
�%EM�FNVl�55=VZdԈK�a�����7�Z��*�=r��/^�a�	�/��=�'�%�[�p�.�7���n�{\��n�%�Y�D����1��,�_�u����eyW�Q�n��z����/��`;!��Vg�Γ���0N���B[�>ݔ@%K��s"A��6�`�|1��%�!��V����}� �34b�шE����k�Y������U;�).g-�C�>Ա(2�䣞�m5��6J��Ud�t���{�P��>=��{�F��XJ&�D�[\��3p��y~�;�O��r>�Z�y� ���*��k&T����GS�+���#��HJ�7N9��=�j��Gm��69��p���k޶Gv-��^�~Ǳ��'�� T	(K�h�԰WQ���|��~l^�N&�����M�v���T<;,i��1� �\wװ�)n/Z��o��Q�N�����F��%'��$d�.,��	��?��^:��P�f1C��"]N��cs�H�`(���H��ܘ�T�Q�a ��D��F�kڂ�H�x$�DI��Z2O��T�)5K(�(�+��0��Ι��S�r�U����yu��`���+O�sZ�kᣦ�7cf1�gS��_��`r�k���pyS�=	60�5�{Z6��AR��E��@[�b���ÝD����	�a�q�M੼�*6���x)����zN��	bS7|��D�9⛪:O����������g���l���c�"Y�ņ�U�n�K���-cZ�G�Ȉv��7m8�77�YV8�=vt������{ ��W������+}�x�q��z[[��|ϲi�|�t��߷1�@Yq'�?!�-E�i&�,2��zc�'��9��,�H�x�d��v�
񳨴��h8���(ӎ�T��F��3c�dw�)�RAgj���_���$K�d�t��#�&��F��� ;�]�4�{��ԧ���yݯ�����,��m�������S�^rF5�[,��,%�mX܁n�|��2:j�� ��GǊ�K�#5j���qEfu�1LI�4�RF��V�K��*rr���F���.������rӁc3u(x�!�@�a+o����㦔'(������En���SnN7裇���>�6g���vS�~>�?��tB�mY6�>c	�rJx��
Q~\_�Q��O[n�f��dJ}���:����3���)c��m{:��nz]B��|�ٖ����~Ds�!G��/L�y��:��6��e$_.y�n��h��Mi�zS�j�n�l��Y>��?1���|NLO�K78Ȁ�[)�pK����G:�PTKW�-Uoݸ��z�<��iܢ%!�Z"^�W?��)��7�ъ
���Q���)<b�w�����'������Oj�	t���SX��x��4\P�(��2n`)51g(5m15�I�����d>���{$��7,N��џzA��#�ޫ�=`ʾ2R&�F�7��W/�j�f�e=�[9��Ⱥ�N*��	��
�Q;~�R߁�_p�M��������5WE��B
���YQ��N���91�*����B$��F��_s����|=��Gk�}�9�wؿ�{�<6����/���C�J~�c���hqxߑ8��0���7xW�?:�[s�g#K� � OKe�?��1�����3aR�p�������Mfgͫ޴��ӹڸ>��ר7�k.*Mc��5ή1"�sq��7�'�d��j�۠nnp!$h|k{��v2���7k\1���ߢZ$�\�~����rx}�1AZi�Q:�_�U����W�9�Q�����vfny�^Ƀ������˰�nb2wvQZ��F���L֕v�i��`jUY����Q�Fv<�u�~Ď�1���pv�����
k��K��ٶ/�)�m��_;g�(3+�����;ѓ����[�7�w
��V�k�J5C4��jt�<����pc��l�,���r��"����m&�\O`[���u�M�"���Z;� ���x�����p�����z�'&������GF_��ɐ�4� ��N�F���i�R��Zv���v������JԼ�l��u�o��_&&M��%.�$�uU��
h��q�A��4�,����|�Vp=�Q"D�/Ռ�g���=��7�L zWH�I2��\�I�⪖������J�)�uJ&�FZ?9i#Emt�{��&" 2)J��Eq#���]y��K;���K�F�_���;x��E�p&��#�L?'}|l��;U�}VV�T#z(C�Xv�y��N��O˺�nG�{���`F����aE�u��&�U�58���ݪ>5%���է�8ac^�_�#>��W8�渿��ǆ0
`��/��spfK���?��
��o"�I���B��x��q�w�d��2*��ζ��x|�s�5��?��w�,�K�nD����މc�Ω�be�M����iL`#V�Mh��t��\m �d!> h�z,��>���j�9��:T3MĒl�z�lw��\{�XHQ�4��h��`����D�5q욾�9��t":Q��7QPB�ǈ�3a0a�P&:�Ϡ�(�'�[�C����-4~M)� �D��$�J7 �e�
�]^Ib��Od��: ��O\n�:�}<=�Ҁ��zD��HTk�n�!�F���]�3j��൥$e��w�*�4�D�~���o�(ȏ�;�P�w]�U��@��qa��z��y׼�eTh5����DG�@��!���1t�`�[�ˆ��W�����X�"`vݯ�׉rܗT����ts+$�����:O�}�1J����U�A��睌`GIOܠ�nX��+x���_��׍˺��B[��.�p�e�0�V �l�9��nce�x�v[`�0${��S,�uEqd�L�$�4�Oc[&X5�s��������в9\9)��Nz�
�Jq��xCo'�1Ji�fA�Qw`��K%�m���/- :Ï6�	�=�
�UzݾP'Y�]�P�X��nu_��G��}����}{J�'�	GnQ�G1�o����S��3��[���88ϗ��$S"��ͅ�M���{K_�Ʃ��ӵ�����V�b��~��=ەIt��x�*Kbɰ�Ə��0��*�Acv�m�Lط/*�H��&D�!��՟�gV1�u�;?]��\�oU��	�7�d7;��Y���%�>��`�����+�,���%3�LP�}h�2XJl�E-P%fL���1��3�z�T�?O�����f2
��W���{�L����	�
$-H���nԠ�U~M����u�S�jo-gC��.
!�-ѐ����ӝ#�1h�<�zeW��~��WuH���JZ��ZP%A��Fぷ)";���L.�������M��MP;?e_ҹ5����'"����-FiC��7}�l�J|��WV�O�,�5fd,)B*NV����tuY��8���8j�/�h��̎IT�Q"�K�Ƈ�Zt2�lO	]�^4up����ȜU��\H�r�ON
4��ytc�%���F0j�����@f6h��[ʳx˧��\7]�#=��?n� �(Xu��^��)���}a�џn4�n���e�����q�u�0���"qu}A�ks���;�����}L��"F��^�5��[��1eφ�H� ���Yշ����+�K���`��w��J�0�%:C�w����ë}�/-	-��6R�l�؄���-g>�L<9�0����Fo0�3V���� �(ɪ��Ճ�L�E�0��io�I����"A��0��`lQV*%!��[-*�}���n`����-� ��j������� Ǣa�^�ӝf��
������e�#�Œ�gԖ���Ը��y|�{�ya&���F��s}����飻�i�O2�C�y�����Q֕�P��Z�.�� p�Rz�$�
 ���^� _(R� ��{[Z�#��t�R�Fh�1�Y���[��l�%�&�l��i�+�s�S�i� D�..�yG`�0l�Ie�5M$/]/�SX���4�0-?��2Zy���yϵ0|$��"����#�9z��ǂ�a�ll��l�M��g�������n�ʮJ����^gS'�^(ہ	7�%�?�`����`Z�*vq���|"UW�R)p���� �o�[��cm�s]�yQ|��4 ���e�6��#OJJy0���d�8�l��i��:LV�jyl��[��µC�Ǫ�%��4 �	?�Qq3�"�ιy�qS �M�Fw����˞���^�� ~^��m����(�CPspԎ@��8oC���/����=��t��W,f��NεW�lޛ�xNɋ��\)K��1�T*�3�㭠s�,r	Iq/W�� b*�GxN$WݾՄ�#�[KVe�U�>$_Gy���PO$3�r�[Ι�8�Rq���&����$mu���O7���0]	/�䍎��a�QmS�Ļ��?;m;�J����C��K���,o��G1*H֕K�uqT�s��#$Q73_���Lo
��N�1�c�.Q,
E��=����s��}�r��M���-�E�Cǖ��!�<'f�����=K��z�������D�=~�N�Ǩ�в���㦩� 5`Ň��n�
T=U{�1�6�vT<2�?����Z���:T��{,�h[9�ۙɩ4���āSp�BTh�0<X���
���@K�6��:�$�	tn0����2'��P	63�WxDC �B1�C�Ƅd���SN��η#w��ƧGG^�@'���z���? 8��ÝJ�$n��o�b���xpD��x�|���\9&�4�c��=[pU@���5�u�~܊x��$�ZN ��&q�ԏ���U�]��ޒI1ۧ��� �UÑ��Ğ����Ij�V<we����ǹ��<|�}��)����vM�2�ݥ�:@5�uE/��k�[rm���n�hX�X�3������s����|R*�(�<����ȗWX\��Q��t�l!
�r$�
���
5�1&ŖWGp��B�󞮏����G�HOf�?�i�l%w�0�3^�-U�~�KBs@7*+��7�̫� oL�X��p��j�H�,:Q5�����a�s��?�Gq���mD��zf�I�Z�����k���z 'ٌ��;��lG���w���(1�ZKJm�"�@.��qx��㞟����W7�|��[�W
���>qs���FSm'X�Z}��ڏ���/���c����}
��?�C��~!\�Vy}f����0*up�l�h�C��u�b��e�����j��gDy�����ꄭ<����<��T
��=����u���}����
+֪PA+�U�yfiVOT	��������N��<�*�2�zO�Q����a����RHhZ<���C�UR	>���'�]a�(-�'�,����+���%���'1aƆ��X�ܸJy6�Z}��ι�I� ?]����	c��]���iC�۽�y�v��%����)��U"��5��+3��S�*@9� �|���)�0�_��<��z����Ȧu��X��\�/�TFB��<���?��=��s»���`Ǭ3ge-�cG���#
|L��=.��n�pP偳Z2����r:=#���)�b��%���-�kVt�V�V����nꓕ�?u}�~��k�	1D0���y��Q��:xH S5?3I��� �6�!�L��lYt��Ri��#{�ҁU��?��mJ�X�'v�=��yVI+ǀ!P��8�Kdk�/�����y2���G���#�"l�ckxmP�$d?ŵ��N!|�Ň �u3^-�e2Y�SSk�/�����e<��	���#`3�|�����s9_Zl�S���tK�9�{�:~��z9����&�.�V6iG���σ�s�Q�MH�I'\_���ڄ���p��Źim���#2#o��:��f��g�[��蘮�m	2V�A�� �Ǔ�Iy�؂w���p�(l'�b���j̓0:�/�X�᪌����`F"����U�J�&�?cȳ�XN�������ҙ�5oT����<�?Y�K|ZI�,���^�_�3���t�N���,<M-��/�F �Y�3B��)n�6j'&B���(枉���f\[����Z�w�	h��<��������e��}��������L;��S�	*;�M�-08�u�?w4G��:��;�0u_,���0��j^�D����<�_�;�-����f\9�H�?�^�r,sf������-N��T��'x�$�P* ����k���_Z��K7�Ü{��i�Ge�ؽ��N��W�����lr�Oz1ⷄ#y���Ƃb�ƥ���� ����#Ĩ,���)�-Oi��s�d��TZ��S!��n5=|T�<�9=��}kC[J��Ј�����ޙL�^��b��i�K��pG�\N����F��e/V�?��NH��I�mQ��5�`��=�~��/���l�X�)�Z��d�Pm"lӣ�
�l*l�CZk��f�iD��|.?���)!m�^F:�:oF �z6��kI1�f8���O0 ��)Y�F����Ո���LQ�zu'�Ѿ�.��t�FJ�mV2g�0��Zzp��Js�E����ڨar�p��r+�-�.����J/��q]U}�w�H'�j�@{%s�:A������j+�5���"��+ɗΡ��2O�p�w�f���g㚊����!�x,��x���綃�4��3��;8)��2*��H�:y�X���ғƨ���i��Ȧ5ϊp��[�Mm �%��������Z\��� 0�+j�9g�<��kPְ��H����|��Q�K��l�(��&2�o�O���}�m��˲N,�v�d����k'4�:�X���J��U���9��%G$�������[k r�c�2B}�8�<�d���u�NR�VB�v����1},Q����]^D�cu�����R[�A{|P�5�����5-%n�L���/�35Zƀ���Ϯ��a�	�"s&^�mu��P�V�z0��V!J^��?�nϷ�3�������n*��Ęh��T�3n����~����AH��'�KI��JHq|�N���9��%�]��-~�M�\+��|h^�=��*C�����M�g�\��f矮aٮޟ��-{!��/|�$��/f�RqKTh]�C.X�%�:��Z�K��&�]B���+Aж� �o��E&YU_4��>�li����ѹ��'��0�0'�ϭh��ƹS��Y��]�ؙ� ��~��zz]�� �Y�Ŋ�%�
��X�0�z �O�c��m5��/{U�n�{׷�|.�X	���k����Jy2"Wފ�;����ߵ�Z~����������L�@S�<�$���Q�J�&�=��9u*	��W��K���|]R�{��劙n48Үg�g�1�jm���p�uu�N���̔|��:']���'�n�oZ #/���C���M��� �:�� i�pۊ=�:i�ҵ�:_��/���0!�>�3g���]����bf�6� �R��2.��sH�򜑬̉F�!�E>��n��J��x�yt}&B��!�Q��RQϿ�	6�x���Ϸ��76  N��2���zM��*�z��CQ��LJs�|�i���1��h�d��z߷����+W`�]�4Pʮ��n�;`�C������~��y�`m�i>9��c����z��.���T�����8��Ia��"|U��?��\��,&!hm�z��"z8���0���O�:�4�sk	bl!���:�s�Z�لMJR ��]��P��l<�<��j���g��+��r��\��??Ò�Qj���1c�6���1��oVO�-=´��y�N �x���vl����\�wEf���~���L;��yxG�[�#v�ŃM��C#����H�J_(�NJ3���=~�G���^(Z��s�Ն>tHi����N�d�i������di�Ugc��3�#SRZ���v�e��Zwz�|x]���=��w7���.C��3.U�5�ȑ�~���LҷL�3��W3���,�yp
��Y���T��j�'��x-�8*>�mj2}��k6�b�`}��+��"��t�C��X�h8b3�V�8x�)=�(g}�՗v_5�!	�����
�{��%��a�Th�	��O"�<Bh�[��.��Ϸ�J��;��Y�n<RƄ�����}�)�nK�c�g���bc1����Nݸ�ܒ.�S�֩�ʉ�a}�K�U9���C�7)��w�����>�Ik�{l��xv��m�v�L�-���Ú� Ky���&Ox����Sh5(��Q_��징�r˧·V�h�z�<M'L�P��﫹I�Z!��Ʋ�d&[,T@5�mu��S0n�eRi���3G��I�h�>�i�I�q|/��B�HBv��E�w��J�C��̡��V�(�Jq;$�Ϯ̜C�>Z�'�ެ��T��A�����0��a[K�V.���e	����ܿ�/�S�/�ڕw=���-���m5>�|6MUU�W9�r�X���,x����>O}2�
�jF��p/�S�SOw�2��&C������1�����j� X���K0I'��1�>�Js_��L�_�(Y��[�J;yXR'^8�MO��Ln��L���P:���b�����|m;�	�#?Ŷ,����8�!���?(_�]��O��8���9�_� z�{D>X����JF�o����=�G/��Ǐs4��ʣ̐ �xq\e=e�<É��a2���c���D�/�.�Yt�9��4j�"k���Wtq)�#�ڮ*��E��~������]o���W����MN��n*��Ϯگ�2��#<G�4�\��%���c7�Fв��Ad:**�X���UW�ڦ�%�:o�~���J�R���f�� M����������2f}�QS��t�0�H+sw%D��|��6����*$�W]���ƀV���e���Fad4�a�'�H �,��g;k��X��1'�x���<�Hc��Iux:A�R�Җs��bkԅK�t�]�8s�۵m$�M��#��)5����ө_Ǐ��k��R�V|�8L��;���A�ܝf�O���T׷�I���^S���fi@��Sl"��s�y$T^{8�K�c�����}��fŗ�F�:�����/��v{�/Z��j�&���q�\�󙙱B"��!"](4
m8:�օWI�X���.�HF�_C��c�}��:�6��w�Δp�W�#�a�9�>�#�r�U*�����r��@��M`J
4�[kU�� �7�#�e'v�0�)�<Ջ�Ju}���� gX4	=�^�w�^z�4��+Go�{$� N�Kz��S1��#���@���:�x�3������1-�fȿ�i�M����e�r�hf7CH���lg��}8���;�uҀ�H{ed��	�v��0���AⲤ��i�ۗ�x̧͕�kRm��|����i�l@��`<�삖Q7D��N�B}!#I���Q0k��Rg�ʇF�oM�
��n#?D.n��3�����Ts�B�ʰ�6q���'ǯ"�a)���A:|�T�f�ѓ��KppR��￢��A�Q��9���[愮�J�N��K=�ȏS >䔕ZT��p��(���q���fMUz��\gy��]&�\y��ϧ����O?ER;�j[+OI�r>(�1zÙ�3
�K��Kf��tu2�֬c���҆�UU�d���V\q"����K��],����W��σg`�ಊF#Ȱ�q2��H�g�Pġ�(a
I��֙���:�����h+rC �_�m�e�7�0����Ƨc�N����!S6"D�~Ƿ�!���Ə�4�����q�O��EȈ��G��>�n��ICCFT�A�������HH�Z
����}Tߏ��i�˒����#���@�Cl�}��OɊ��z81�=�K�mL����(�:V��U�>�v��
�茷����1��̞7����s�������Om�㑽�B���&�k���Ja7hS�C>{��,��|T�B��L�]2�L���x���kXz�#ssh��B|��V�/Y^u/�(x��=��
V`��t���3̧wG����E���kb���Uy���V���#��E7 }4Yt"p��E��X(���ҩ- ڰ?���ߙ�G��W��V��)Ô��'�1�[gᗎ��j��*�I׭r��ݠ���β�������n[�~�y�jZ_�i����8��{�K����V���(��=�B��WFzD/�esx�q �=D��{.Y{����eᯧ��}��Jg�̛��!�G��|W� ��f9�M��\&��l�=][������-�f�c��y�� ;b#���,ɰ���q��e�)����z;���Cc�#sYBa���NeF���3~!p*�JTftn&�*���e~����DKN�0���/b{����d$5o���>m�A���P�]0���� 8/�s������c��GZ]�029��ӊ��ΎI��..�����;oP{��!�rҲ��� x��H�S�H�4��x��D�@�˅_�[Ö���T���-,pű�	F���F�DA	q�z����@r��޵Q{Ì����QP��X��O�`akvة�^�/#ID�Ȉ�D��F��l��ݬ��al����1�h�Z~�G���/\��`�7#R��W'���I��<7MŨ[��=����������دr�b�_7�h�׳KK�d3��.i�^��L%������F�d��Q�{��p�b=U��k��o���@����_�AQo(���!N��ұ��\��v&�� �h����q���A(�
�ܵSvqI�2��/m<��%o��;�+��f��,�>��~;��tޓ�<_�xؑ�Ab���b}��=�=��A�\��2�f�u���^��� B�4X�6����YRni�~zep���᜞��RqS�'3K����Nw�K�AP&0EH �\�'a�ۇҠ��	�չ1n��/
d��"�#0:tNp,����3KeȖuMr�	�׫ q˯��)����)�jR6�u�%����j"w��?}Ey�+����m/13eu;��5���f7o[j��m�����S�O���2���	�S���i�� TS��i
�Sj:�n����/f�_6���}����5�`/��<�Jk���e��e���ީ�t6N����7k1k��al*!U����v��_)/{��|��S�+����vYW����O��G�2X���%f�����W��-j�섶/?4�;V*��HɌ�pT�&�R"����**�(3to\Օ���[��J ������\�c��,=J@^�y�|j҉���Q�UM��r������>2+/X���:%�Yߤ�+�m����ڏ�`�m%�ݑԆ)��1.{�l���p��Z�h1o�,�����U�7�FS�\�*�a8����ŕ��>��k:�6�GA�	�/aښI�+��G��e7���xK�{#p��^���|t}V]a� k<!� �d�~V��j�lk��c,C�8־�#G�H�Ng=�<�T�|�����̤������>���.yvʯ"�#M��&�hv���d�A2N(w�2v���C�;��Z��`-�x2rq���RN��gy#�e���?�m)|ְT��_�!��5Y�����a�̥�"e9��T���l����i��=�2@�?�}Z�c�M�E̢Z*��L��J!�,{�ibNS[��wѢ~��̺<��B\}gqS�nw�~+����𶕹��F����0A�xn�Ǣ�m���z�	{�����
LV��/0і�0%;R�b��/�R�7ɗ܆~� 0��E��mY�~x������r��B��	ަ(���B�h$b�P$-�%_�����Rna�8�����W,_�'c V�/����ΞyR׎�Q��ɼ��{�(Md��pZ&~ �]�����5NC2�~��t��8f'�**���B_���;o�9u�ܱb��m���6��3�q������n��/wQעu>h[<����C	�F'O7U�,~�^��\K���
��}�!��:2��X�+7D��bZ�;m��� U�\�}6�@<�s��r����"c����^F�.�ө���86��޷j��n�1:{��Yi���s)@��^��"]�I�!)A
�0��� ���y��Gf�:|�=�^آE��M:�iti�]b��C!�fcW����u*�ӄ�t5��a�T:�&���D�)��c�����)���~�E�Ž��X���V�;ER~B`Z��9�����0��e��JP��
yL���Y�� I�a�Y+93�yK�&T�**YV5��2DU��i���9�
&�#f"�V"%Q�z5�+ ����n���@�_zC����tj����b�Y�%��`n[�t�ₚ2�q̅2�!�����0�w���d��0Tr�н}[MI��rڣ��b+��b��^L�ޓl���8Y3U/�#&G,��橄\>>��:��������:��Q���o�P�����!�5�p�����(OD����G�nc�-ו�4�--����W��#�r�wvҺy0�S�'�N�2%�\��͇0ϑdL��s�9|�=1�<���M���,�/��G���>STt؄�H)�8��L�\'�Ɖ�"�������̘qy��5�9���I�� �ճ�@м7_/$c+����;1a�dbO��]��Ùz{4�j�EDD���`�ꃲQL!�~V޼a�$`y��c`
��:f�Y�2��Ճ;�y���N~~t��x@'(	"�χ��j,n������S<���8�\:���a~�s?�k�1���M��n��yu���˻�x��z�
��7>R�H<]�'hEQ����<�����n$���2�~L���h#�q��MC%�5� [[��Xj��zw�Z�`�W�+�\{�#v3�Y�~��3f]�9�G��J���i�	#}���ɓ�j)�w��d�^�
'��و��[���e��i�j�i�z�g�~:ߏ����(HVa++�0��F��<���Jڱ[b���p�.�pm���̥� �'��G�8yz��k���[�]T�N�3�n��\�$�[zR��Чn���Ђ��}KCY��w�w+��%�U	�FE���I����o��c�i �?�V/A�T�m�/I��ΑI9t:�F1�	�]�e-�z��u����n;k�N���ML��룩���	��b����lm�_=�݉������suR5�`+�=�=��%�:�-�bY��>��j0�������~<�f�Mp:2��D
�1<p+��I�Q��N���|i�(��+������ �ڇ�Hտ�&Н}�/#��/����4u��7F�Y' ն<���:~�.��v.9��E�^�S�:�x QH]�J/#8u���k��Â��#8%켛65�A��Į�۪,t"A0`U�� r�Rj
���$i���o��\��r���s� :=�bod��P�I9��AT�ƞC�8���zޜ3x�JG+X��5�V^^q����OA���r$�h�̯6Z:���ݶ�^����b��#C�0�2�n_���>��P�"���B@�ex����׹�ح�'4����#� ^MZ??��W�0z4����1B��̘�J��5�m�n���b�O���7;�>��v��h�[0����%A	n~�p��o6�� #���� ��0c"o�񺎷�Y�rl�k�9>2k#��j�����L5Ǝ��T�Gݸ7nt���y�l�nb�;���9��~�b�~����*H��-H�gRT�h&O�q
���F����B���:�&�n�!B�7��Oc��|w̞��E]r�i|)�#��Kiw�Z�l!^��T9����!�Y*��e�����g�@S�q˧a�7+Ca��[/������������=�,mf� ��ߡ����>L�o�~o ���"6*�E(N+�����&��@� cem�a?b���+s_[Z6d�v<�v�?���}d�g��	�9���I!�� )W�S� �i�����&Y`�O�{X@>�ڗ�����!#|���J��6ȽL����P(E�/X��-��1�?����NpS�>�#2��G~'%�α��'��8:�IuW��Q�2(�.*0���,������5m�8�
��[��;>�o�m�{[~U�y'z迮K
N��w�~�2P.eiֲ�v�ªa$�%+�zB[�{� j��YY4jH������Q�����+k{F��_"hnM�D���,��ﳲ�"�*v@�1���q���:��Sj�� �(ˍ@�����:�b��+|���ۢM����w[�_�\ov <�J��������gu`[Hv
߃�x�X�'c�my*�����R�(��d/���X�=���1�3���HS�7LX�=�="*+4�J`��@2�F�$�Rg��pr�+����YUڵ:9�tqӓ��?�\��x�?��V����c2��!FO�3-����T����a��x������j�5���?����օ.�)'g�?���>���e 4�У�a��9v:��X�e搛#2q�I��G2�I݉cy�͸��R����_5y����ټq��NЦ�4����n�p^����e
M<gq.������lAqlF�0�I�^���N�,q�V�b�аI�Y �D70�2��:�	iĆN���I�a���:���'ZM��f�����x�L���m��o���SW������"ءI���i)b��������]��X�J&�2+���,��ȉ�>�&e�aɇ*}�?��=� �fX�����.�����e�kd`~1�0��f\����h�������m������A�+�����3W�E�@G��V _�Q[.�ȒL��mf�P<�Ks�-Z�Ga:1���Q�Z51�-;�M��<�O��j��ɟt�<1)�z��������\ϳ����j��&�Eз���wV�������|G�1h
h�G);!f�bc�`���M:@�?���h뺪���Z��ܣ�!łn���m�$r��hD�a����Fz�K�"!A�R��	��}F�,	s$H�
�:�����[z_
���<���e��������9=
��n���{6QR�+�<���V���|��})�;+63�eORHѪFW@
�1�}B�h�6����ծ�V�"���*�op4(>�+���2{����\����	M��#�o���yڧ
	Zg��z��U&oG�W�:�D�,�SnM��Ad��k>�P�/�w�}��ّ11_Oʆ��߃s\�-	�����^�w{�����qX$m�8=����A˶�I�������mf'��Re���z]�N8V&�_��F���t2���QO� m"�̳'��4q�����:oT����l$k��|0b�di>:]RLO�gS�T@G�_9�� �y!N�}���t�aM>ޗF@@D:��"��*=	��F#�R"% %
R�c���Ĩ���hF�������ܳgϽ��s�s�[���Θe�<*��~Ǔw=ʧ��n
'��g�&���X�]픖�G��!�S��ԕ���:c��z�M_�5�h�(��8�q�$�����{#m�����C�@�ܷ:�t��;��tp�q�[��	�.�1�� ea;�m�#���Nc�I�>*�{Y��F�MA3��Yo*^���������Iq��Z�+�h:}]7�7�p��q]��r�)]��'��օZ.	�����{�d��|���8���0[M�hf=ؖ&*��'����1iMp-%��H8]\i�RA��ٝ>��m�k�U:#Ƃ�-�����v`�Ӎ��1�^]��Sa}�R�4�y���~�rdl6����TTn6����&�r�f����%���Km	�wL���|G���/����[�4|�K��h���	�⋗Y\��i�Z��^���A�O�,���L���)2�D�Gu�=b���q��3���2gQ>�4#�K
W�i��d僚�٤���3�JN;��ٮ���ڝ;��ѵ�fLPp�k`O�=���'�ל�U���2��v�i��{)���;D~k����;Rs���Z�6��h;m�8O��v%/#�Lݳ��j�?��=��ԽF}���0�+QD�C�Q��b3�UCB��(?��Y#-���Xy�����Pz�"fE�����Q�jk�@�L�!�m0��n"�'��/ݸ����|���6[њ��ʮ�@��G��� ��Dw��{󆂜�㧃z�������L1z/�^����<��,ǜ������!W9�=w���8��a�������%����b<a�k�K�~�]3(�󔆹!]��ɴ�������� �y�9�G۟���0��n�v�U����Ʋ[�!��4	.+������8�����0t��D�F�9��a�qO˴�&8�W|T5�ݱ5��ѻ�*�w������n�{���Ƣ��vzp~_��>I�[�~{<�A����L"�|(�׿/O�q0�d.b�w�{z
����fF��r�Ƃ���\]�W��;4�J��|=Ǩp�~��檭�?�I���4ٕ����6zm��C���G|:�bx!XQ�M�J����^��+��f���xULQ���ǀ�h�+w�G��$?�/�ܸ�K-��rwX������QB�L�0��"I�U�J�!=V��؉���%~��-n�p�tW�O����F�ff\Y�`;ȍ��)�u����)��w�8��f�gkURH�|�Pf<6�v�Qv䉼
����MĊҭ����_��}��6ȭ�����ș[%�Uʀ0J��L�x���u����6Q=��@P��	�K?|VёiM�+���s<l�%�$s����{v����J{�+g��[2E/A�9��q]+W@�K����X�ˬ���yCD,��5e�D�����e�ڢ���"y-R>3�g^G�%U{���1��1�ըU��f��ģAo�']l���/`;d^W�O% ����<q��|��� ��O��6���]�	�f�V����w
:��3+���?��p]�}�&��v���o�̷�\\�Y }WL��
���]ޛ`!��t�,�5��~ј�s���
��ϗb��l=>O�s/�b��;t��|��!��F�Eմ�?e�^�">NuL���e\<Hz��j���T��	��VQ�c�L��W��s�]iw�{-�!��SZ�kW�����4�V{s�a�+/�AV�꣩N�igl�Xy%�AF�8�|"�C'JPE�qǀ�=Ε�/fB8s����O"�}��4'���6����u��^�
}SӬ�g�V�~�p������p�;���^Tn�{p>L�6[�ؑ��,_3R�G3���<�[ ^�W1�A�8�6>/�񽓕2Z2S�0�y���s�BU�?�J��L��r�+���=u�Y\����k�y����R�r��.S��`��]v�̿X$�W[[�3�N���w�N������#�!WO�/�g2#��ֲ��=�Q�t��͸�aط���!-�n�w�K�ӣ!=?}����#8�.ڤY�S��0�1�y|r��j�)�L���mY)p�k�-5��M{����J����b7}}��lSj'��b����Y�����&/����ё�F�刓�<�̪��wr8��_ڝpG�.�v�v'�����N�+��y���?!gr��8��?ڮ��-yDT�dj$E�n%�N�0�~�:]�|�����V���T6�N�_�8n�(�I$��f��[�M$��n-��ʉ|}��U0��IvN�f����U�@9��}g�Q^�����l���OX@��s0�G7�bGI�A����V�̏|2r������n7:��G���������_��<�ߧ��eo>���127�j.�ܤ�Q ��ټ[�p�~�>^O�vc�dԔ�Ѕ��lU���V��ޣ��M�Q��3
I?�g�ojD<y�f�oμ��ID�M#f�G��/��wp�VY�m?�zɌ�����|�w��D�/l�ݸ5�H�9��/�;��a�V�H�nDJN����'e�
~��:n�3M���9���Y�q�l�Uo����&A������L��r�ɜJ�d�՗Z��,��=�3�xW2JRW�'	�Q�ч:���9p/����{���e�]R���s��'��XT�,y{t����[�F����R*0�֣��e�:2h�_8����S�p!��/4��{�T�uPXj�����T����̌��:��D*&VY����(%����p�^7�
c-�4+�,sE߰� �>g �n/=�<B�	!� 6�YS��=��W�dD|��/�� 4QJnWc�7<�t��@�������{�r�+��o��o�C�1۲�ܠ��Yx_P�9�ȸ�xu늂yk�UI�-��@���m(�i�#u���Й��s�adeӟAK���	�a@�Y9M��b��Sd@�(f��RF E�9@>P�5N�}�^��j���Ii�W�F�I�"-)�w̿G�֚��<y(v��Kn3�����\BeF����#��.�ؙ���9��|@��>Up�٩���;����`zrdb���ߔ����nИ����jr�����C���2g���L���r�%ϸTǕ%n���]�/�۷�dQ�Gc�n�\��� �����fR�#�<�!�|=�{u������p�+Gx�v�1s�`gS�@k��圲�/�~�bs � �O<����>9����� ����0��z��Ώ-��a��.iy�a����C��n/�~��5���@�k책˨�
=mGm���}Q���-�)��+�Cjك��?fQ�"�v����ac�p�%�Ƌ�mswG��)�7�c5�"�yQ=x�Դ�iD��OT�S�4��gɚ_B���6��ј����G�rE��j*0N����1u�����D͹#}�����;-f�Ϸ�ٕ'� ;�g{�}/�Ƌ�Gr��g����`%�+PX���M��u�.o�ѓm Kh���q|G�V�r�xg�����j��D.<<՗��v�(�Z���O!�8OR���v6!���sqG�'H����Y|������\�gyXi���ь�z�P���H�jz�Q�h'f#�=ˡ-�f��m5�ʪ'J�S�U�x���\d_&��fA�s��x}�.��*5Hj��ۜ0��Q�Tc�{W�;���o/����W>�� ��}�ة��(n�k�C��}��i9Y;`r���e�c��*�QQ��EWf�(��eș�ØmU���n�S�ө�N�U��gL�ߵ|��v��Ԗ��^g�uSrg-X�`��Ĺx�����\�X���9�bkQ�� 3�}@�76�Ճr��R�S���b�?�i����Nӹ%A+G)���f�gc�3����P5C���yt挂(�����Z9�g�m���s�ꇐ1.���5/�q�n_����	!(E'x�����ą������O�{�Z���LU�Ql�I>2��/@��� ��|ل�*�$�B�H}�L3��7*��5�dϭ���%8�]mݬK"��fC�Q[���T5>��� @���R�K�XҮP�k�۪�Vb���#ޗ/�X����N9�����p�٣��������~�%)�^Gh��|�+S!*+�e��9�PU�p�=|%Ǥ;�\��Q�F#m�b�oR��'(���h]��:��dw�	���?>���Ǐ|#���l�=�\�4����K�w��<݅�'{��\���"ev�wE���g&�t��h��\���&���O� IxB{[��sT�9r�����Q�p��h�)n�L�l�6�Iޤ����{T��`���`>��zj�	%b~j+R�+J�{�j�Nד������j�g?������D>ā��bZ�=�Y����H�_ y�c�P�w��t�$
(�&���8Ja1�̯�'"�-�A�����6��,�%X�(��B��'��O�d���M�+�#$ˤ��ͬ���nQ�}K~��4���kA8��\� �(���6�X��A�p��8��G-����ΉIW���EG�G�x�_4�1�D'��}�=*we�U5���P�A�"�7�c����y��0��E�6�@�gmL�� <=6�����c�'j�s2ս�tyLC"��3�7l��ْ<}�(���γ$�c�J�Oա��r�� 7�?�e������xY�>���B?��R	97¼�� տ�R8��J�t���ٟR�A�c}3�g���۫컥�����S	���'��WK�~�/	�9s
O�� U�'��Y�f{҅%���_P�=4��i�����0J*��s�cs ��#x|蛔s��(p���QlY�zx�_����a�I��ؘ�&&�?��Rr��˥}-� tKv@>��Y�cXf�2�o3�(�,��`�v�V��'TT��n܃2^f���\�d�^��=�/�����I��p$}X�^/0� v]���wq�c��s.%�-�T(h�wt~�
t=%���b���k��yt'���1�����y/#=��Yڂ7�d�Pg7�"����"�ei��M�M��-�J�z{�;��?��">0����<2'g\���O4~�"j�M  �.r�;�)�sJ ����Ҭ|/�l�pf�ة;�͏��~f���4���y�G=]�]�Ħ�;X]��c6f��I	��(�q&Z<���FTP:n�p�L�ϧ�^���\��.;��x+l��Ի�)X{|3�#���r��X��?^�� .hW�zʰljb#M�jZ�����z��;Ǵ�.��s(�-WK��z'ȱnW�B�?��RS$�M��,I�U�殟X�.2wN�~{]BW1���y���0�D4�C�#*����o��)$�+��T�U�o�M�5�� �Z^������ �������fgw�fy,BEXIy�H����4+I����t�c�|DH��j�G�+D�L�s#JAg��G�q��9�%F��X�o�y�Z,���GOI��g^�K�e�xK�*VT�3+{�U��j�7��4�z� ,d����36MԲi yp�i��R�~�LM��Y��3 ,�d{F���s��}�;�L[`V��Z��˞��%��솀�����Ka�Q����1gr������[�!��a��ɣ��w��*4��/r�5��ήe��4��S��Ƙ�7/3�� 
���_���z7̦��L��^
��Q�,��5�V�����7�ko̠sEhF1zU��/M5�8$Ė>I��,D�j<nz�Oy��@�*��B	2
�z`cg�ں��F!|Yj�.�h��{c9��o``R|��J�e@zlg���FU62`,p�6��o��Kr�*<y��A��gI�Mk��D��j��0'�<�g)�eW��W�e�HbR: �r!!{�,��l��7-(_�v]�G�z��O����|��|����_���x�7H�t����X/6a<���=��0�eJ3�{_x���l��Xycƪ��x�B��a�Z��u��xe�A}+W>��'���Hu�
�a����UQ�	KK�&�����
o���C�PoZ}��K}_k7�m��z?꘿�:�i�K�g2j$���8���f�֡<��D��T������tݔ2i?2]73�L�):�]�t��_)��4�#+�J?�6_���}?������ő��ȹ|Ñ��.��;����+��$=�$�N��\�w��蛵z�ee�~2>7&=x�e����<n���2���n�'��20v��n��hC�������_c���Ma�w�a1!�����c�]���v"
qa�y�-5)���e����]�n�h�х�{|��=�h9Oq(���:�'��������^��E�y�9��Es�cՖD<��Y=�{�Z�R�"�(	 Ѵ�S�(�xD�-Sc�$=|�����h·$�*.u!=6�B��>�e�0x�w��Ks���~[��&�@�����m"ω�U��?����\⩏8����5E���ct�����,N_�����ޞc�A���9�N��4���p�~�	p�#z������YC^+���pt����l��|�Ĕ+�>ÓM�X��\��y�O���GD˃w�qw$n�zG؈٧�y?w`�A?��韒q� U9���;�y���f)��LU �,Tã�|�A�<4Y,�e�v�͎�O3FND,�#����_-��1�q���S"�ĩD�5�����Jl�0�F�$n��3KP��\ݮ�bv/A޼|���:�����# w�;���%Y��T�e�Qg�4��qoV��{�=(�V�p���@�n;="���s��:j<���A)����׾,Y!�j��@X��%aC {���	�|�A� ��E�VDM>n�Β��®��0^vJr��R!��	��`����2!�ޯ��S��ډ�Oa�	�r��hP ��=��'��L]Ͼ���N.B�IpX�V+h9�]FC�g|��8�-���(�¤vmR	pu^n��C86-KXϢn?��/lh~?4�f��r��(��&AW�g�L������ޔ\�_��\W�����߶��5���C����Q�V3����Ý���]�0	�~�!��F%�h_Vvh#n֟����ٌk�){�p����G�E����6���f����[�sC޲�A�L��Ȳ�}^3���n��t���6��@����:�S�����I�B�� ���i�5�7�w�L����.Xo�L$�à�Iy�
;�g_�$��W��{?�ٹ����f'��
xr��l���.�[S����&�eze���<Bg^�噘%�Ss�t9{�%�c�.��6Zn�ᣭ?���ͪ5��</�o��c��G����%_)|FSTi��EO�g���a4|�ܿ��A����7f!v�bn�[�_X6�i5,��l2��<���L���Dy���t>��^ȧ�}�$?C�F)[�)e�c�S?E�|l�d�E��̓=�\�6v,��T�U~M8;�ń�e���~6����YK�ճ�ʼ�li�@�T��Y.&��xϧ"��tN;B��������~M�x1�(^�t뺺����֟}���� �!�`��\�x<��9���t�z���J �c��<��1�������/?�=#��Lj��@\�o
g��(�
��|[=�a3�m�g=�-�<��?�N�![�5�A�7Y�Ԟ⻔�q��l�cU"��!�S����ߍ�5_�ѤV'�?��LZh=����Y���V�9�]�����tVqnW�����sJ�pk��Z��mݤ��ng�s�Ң4z'��MFu��Ziw�^j�\�`D��B�vLV���*��������G#��%A�Ơ��������9����� ��/������1��2�ނUu����U���UĦ+�� l��?�`!��$e���j]���}9��ip�T���l�2m��ng�C4]-�<������e�Ж�j4�O�cdW�!o���pr���/�i0��ʹ�t�Ə���lCXH8:,Q�'��`�����	��;��κ%<�'5q B���L�">�Ҏ��J��Щ������6*!ʙ؋��(q��!�z5i�1�.@�H����{�7�0$4L�;=��L����s�|�b�z�m���ƦK��{��K㲖ݡfU;5��:x}-���y`Q������A�
�dJ˛��s*;a�{go�=�"d�	����]�4��ry0�[)s<��ͱ���-�IOy#�y��H/R
�07���m���m(|
Bic��_�y�N�@϶�[0� �6ݔx�Å�J_
�x���Q�u5�s���|��� �햔�F;0j�r,!��5���7i�Yf�g �y}W��CX'��;;2as��D2_�i��Zn3��|ft�����"F�1d��tpb'؝�2�iϨ�Vu�~ �}���H�ƊLs��P�_1�F�Ř˵�n,q4�b����������������=��J�6XwK�&�� +��\!lI�#X,F���P��7=�S�s���3b����j鎮N�7y� �nI�f/U��J �IE�9Uh0{�0r�_�`�mY$��y1��-�Ew�����Wi��fy�ݚN�v�x���Y�����6s'����J.�N��vE���{�̣ޜ����)�C�j}��K^w���A��*��2�[Sիf����P[���D����Ί��-���i�6��U#��>Y�k,�㹝m�@W$S�cuiMٜѾ��Д���g6���Ev�|i��Jɱ	�<�"�Q$�H)�E����󮏞	$�N��A_�]y���E58#��ز0m�XdH3�r��Ɯy�v�X�Ō���"�gy�d�����i�웯���̶i'� �ۢS�p�ݬ7����d��=��
s<rD~���{=�L<Q�.�ӥ�4	����n�;��	��?��6#YgJ�u��]Ce�HA+z���-ܪ�_>Y1]|�=��g���O�h��2���d�gE�+J��4!����Y��g|���2�y���H_����wq�SD�c��1���� Q�N���~�ʭsn���UCu/'�"�Ӽ�h�h�G+{�^��3"
��]Qx��eyC�M;cDEXm�۳BviΚ�l^�])Gs�V��|��(�|#���9βf��d�HxJz�B1:TW�X��K��)����Go]�����X��J;�]�سU�K��GF��A+��n��԰���^�{$���y
ퟡ�*�rqL���{]$
7�0N����e�jч�N�t��j�2���������{&\9��Rf�W*��%�\����	�$wm���A��tЅ�lۤ�e�[R�`��E��2�����~��R� F� ��J	��i�^Ղ�!Oڼ�-j��0=%�}O3/D���U����3���~�u<r�[�/���L��
9r�
�l"O���qn���:�C�i�� ��֫o��p�C7\3+V<T�-����n�{��Q��o�vb��]�������+K���G-�.�&�@�n;�(��[���jp�I]=Ɠ�q�b����:#���mt�=��@ܭ9�������T&�F�����8�I��N#!r������	~��u��שׁ���Ġ�6f��m�<��Z��|��$J���a�S
Qz��bQ���s���(��|!���PuK��o��"�y��K?�W�s��1̈4���,���ɂA���w=K�}����%����fr)�D��p-}j�s�Z�IמL��+�C�L�� ,m/���J"zUǌ<Y����n�i����D]�����ޡ�ֈr�y�Ƃ���a�� J+8��Ѳ��ȱ�����J*�	��F;-y��S�kEa~Rz-�8��Q����
�-��;�cgHq'048_��"Bo�ұFͮ:��ƒ�TiT;S������ ��%$.��>��6a��x�T��A~���P��`�nm�๘��'/G�S�gUW�J]��X�{��Y@��?� �����ט��
��\��J��]^�{��4��	X�"���8_P>�9Bن�ِƥ�L\n���_+`&�^稳���o��	�+΀���~~~`E��l_ŏˢ�fw����c�j�d���^9o�ӄޮ9�ǯ��J\��ms�?b���P&�[
)ӻ�����j9k�l�I�p���?)�2�Ω�6�&k[�]ڣVL���MT�#�#����X�ѾlY[j�ƅ��K:����t��S"��a|��vM?���v�Og_f���Ħ�%��R]�\��9X�`Q��C��z2#_��Q{�ْq�'��}�E.��.4�]F�9:'7R����^Il����uC8Z�P���-)��4��K"a]za��M%a�IW�(�~�_���i��O'�3���llN!�}v�;�
�)��[�-��]x���$��%z���tr#�`�t}/�:�M��]�I-Ľ�om �������LA�4Ne�܏��2Ъ���ҿ�[���{��03]�f�Bi}�+�)]O�3u��v���$���v��̋c�B��;=�ݽ���Og=��r�tE.TF�Ϸ��5ғ��cX���M�u��?[�shB�s���vױ:����@Wp�La�+�\��5���&糙Xެ��������	A��0�=������|6��;�C��5|˶vx��@=���c�?M�]�n���z��@�?�3�^R9�$~#Zޅ��ZM�"�g����B���#�����Tq���X�$.�n�L�-�\��=�j\���v&�,-�T��4�$%{����f'䜣�ݱ�u���~��/d���xl��w���~I1v��n'�e<�;���R��]����qN��b�px �V	Ǿ���J2G�m���#4��T-�{�p��Ew[b=;�b����B�ԝpM��bd�o��t��l�P�+�\�|<i�?���CE ��A��GۀI�ˁ�8Kv4?v��AU�S%�i�P�[��1bL���!N�=b�nj�)��;�8jdo���Ch̶�Z����g^(E�y7�9��s�r$�R_�+�Ƣ7JBj�N�z��~���^'^@�s[Zͧ��֩c:aK�qq�pE���������"�)y���6.�͡��t7���?�Cg5'?�^W�0������199�W/ �/�;�&���KUsrDY��� hDFߓz�ց��~�����ۤg���.����8Yv�pX���n�WC��?`�%��p�:4�W�;�w�m)�U9.FE�j�(�M�g�Q��{F��	�W5���n�O|��W�z����-��^s��bb#a���&�	��C�!�X�cމj�ћ�)�	>��1������ق���|V�y�\E4`�%@�1�8�M�����U���H��B(��/n�� ����~��ˇ̔�-����,�Y̽9d%�;�p�jku\�X,b�OE�w.(.�:㻅}�Mi>O�P�$k�Y1L���@�r�(Q��N��R��=ya[��Y����X�t���A�ݿ�v̫��\�s�Ȓ u�@���:c��M�n�*d��Z~����H`���BV��6�V�L/�i�oq����Ɣ+8o�$�VWM�V�;c}e�
���$�[s'g�_t�oN|*��W%r?�ؒ�
�����6��Bn/�������4'�v�teiew�<��B�]˕�(5����s�S���!�5�z�=��HZp{4}t�"���'l��g{D��Y��Q�3v���u> ��gc��H �`o���Q�r��+��5w
�ֵ�����Id�n�S�̗��������09�����:���d(T܏�V��{TF6ѵ}��)���Q����k���f��9��wq�84@q9��<i�;�����\oO��J@W,�Hv���1�2!�x��KoӏR8h4�sϬn�i;(L���tR#�{CG��{�� m��U2�%M��}i.�=�c���=|�ʓ�sw�/\/I!��"�mpP'6�f�{�u�Ф��/?���wa�-C��ez�~Ť�^0����WÏ�/WD�^�C�1����������~�/42*e�'Y�ی����.>�1�#��p�P�o�<'��?�шc���k
�{�O�����?P� �������ݭ�o��k���qOc�2��&��j�7df�����v}b�M��,#�d�xV%M!�444>2B���e�?��g�A��j��w���N�IQ�G��_u'�D��X����5���?���G�N5�OU�raߗ�;�z�R�Y�T�
-�a^�+1J��0����n�'����`{y~��J��!?�.��O y�:��L>�.ԟ�g�kݣ�"�Y%�p�R�X&
��m~ĥu/|vl��υ�k�Bg�k�޹䅔�,N��^f���!D�v���|��a,��o!OSU^<����T�S��uVw��i�X*yx4�MBP��*;�僽�T��^@�\�dW���˸sv+�M6�flb��г��W���z�c�g�C |�� ~�f��H�(�*�4tO<V1��&"�!���? �Ͽp�N�_I�s2K�6�|�&'8�w���L�B���|����mS�3�M9zN\n8�)`[�;�zm�CZ�+6�`����^y�{�r�w����v�V�Y�zo��CnO(c3�&��t�Zx��G����A�KH�DU!�qH��M��]��?F�4^[!oJ��8���>��Y���&��nٷ�sJ�R3��N<>e�n<#L;�#Ԛ�_V����X��)�ܢn	3;"}�yiE�[L�����!Bp�(H�����EY�)^��_
���֑�q���pJ��ԄSup72Ƀ��K�?�#>D㖤�����Q>��|����,͡F�Г��L�����c0����+�z⣭��@����kV���&��7��)F@�q�;ߺ ��/jT�u�N�4uӞ[G��/��i�ꆛ�v~��R棰�6ϝ}+�����.G�����pe~�u��~[��J��!�L�~a�|ܳѺr�6���j����D__?1���Q�G~���Q�JK��t�0�<��z�Ȭ�uV���/;b~]���G?rCl�����7B�Y�kE����!���ЅW�������å�v��C������f):,֗Rڣ�7@��~�йR~���Zq���I��\k;����ͷ��1Hq����K����m8��m��T0Aa��'��rctn���
��nx"Gh�ￗ��
m��?���䑯�l�c�i�E���l�0˫�j����b7��Qߕ�]�/}�b��ޝ�l���7�<|x��κYO�e��'ܱ�7����x.$��=~&3&�����f�9��qv�?.�Z�n�e	��u�����寮����S4�!��J����<	/@9H��ݢ��m�EU��z?|,�t�e��@�P�|��p	��xם�-��m~B��u�{���euXH�/�=�p� ����)����ߤ�(1L	�'�� �����r��A�.���;kKc'=ca6o�����T�J�iف�:��y��tI3%D�- [��IPYetѦ�q�ĸ������ϪV��e��	.V�'B�.��3;��K�F�#N�]�MKT���X�7���UY�?�Ss�N�`��$0R!|6��D~l�^}��}���r�\�'��3 �ƃ��V�|C��bfk�4c�F���L6�kV|�p#���vL��P�3��N�gǕ�s=L���������G��=�8�v�����0�ɂ������b��߽su�'�ֿ}�@v�\�=\Ɉ��Jy5Z>ׁ<�,M^]�k��U� ��6{���������[\��`�F��׽��̳���/C��L�}VY��w��d���������q��r�ײ�1ۍ8n|.)�'�PG��O;Fê�� �x��_u�9?m��ɖ�8� _��4ސ�9�m�cN5�%J��V�Q?�f�+>�?����F����-��E)�K
y�w_�IM(�_�A� ��/|��?�m���=T��FH����{	�A	RH��9˴��se��݄����m��)���ҠO@�gd�ma��V�
q��A9��zZ=�s r��D *N���
9j�Y����B�>���o������j�`�s�{7D�����r[�l[��#�>�`�<+u3��Fu6���>$@}Yhh&��-U�R�|������S0�4��4��u��Q����y#�
P��=0
7�p>3����2�nP�^&�iH�A�߻�-kpO*"�߿�y�K�/Bj>�o	V�;�-�8�#�r�:k�X<rjD8��v �Lj���HMya;�M�̖��a<Y�`{����nE_B�߹`y�=ޯ`��]G��i�Ym����[]ٖ�ʚл�c�����>n�Ԋ��Hd��	���`�$'P��y����Z)j�Y����t���>��}4�Γ������-,���&���\��r��i�$�[�/#�lKR��n�΂�����?܂�/� ����,�	�r���h�YC>�Y:��w���݌ͳWi���9jX��υ�� c�L��"�3�@�+�[�Q��'��^�:&}�t�t��4ӕ�lԴQ�
݉@C?��~���e���֫r�0����r�,�`Խ���:�\�7����W?�8���mL�_;`�b��/ϲ�������u�"r�G�'��u��ck�u���:#Ѯ��A� ;�_��d%�������Q�q�6c0�[����q�2-�Ē�m�̫��0�����W�( ��G'T���ֿ�|��Dh��� ����KAs��m;���;��!�US]��I�쬗��o�Wg@Ma|��Ѵk�΄����	��;ƈ����xt��oC�;`�����ګ?��/�r(56��m��P�4yE��k��=����{�k����V�����%̌��Q�sgzʔ�>�tn�I�o�4�(����(���ڼ�*5���E��H���Zyk��x�|Y�s�B}�+���Z�w�{��ȳu��>�.I�b,q)N�����s�*o΋�l&�
�[�=Ҏ����hj�-dw'�����O9�[�78�L:jV9�Z�L��d��܀b�%��H8��̸f�|���Fl5��8N��P��ͽ�k'�¡7TW|����kcY+lW2�I$+�����>�Fe*��+D�31Fqhg���m� y�S��"���J��������/��M5�"�v���՗�k����j����%�_$乼��Q�i���IY�J�o����1�*n����ߧ�w�u9��:�3:�{�-R��hS�V4�X��P�#����J�;��g��F�0�M)C��LвqX����bn~$�d��&�*�]?�:�wટ��f�~W��5�]��\畠��<��<OH��\V�3ⶪ�=Ų!��ɕm#W��9�8o��?���5c����^9Ay^�Y1��߅�W�y+|>�z��878��[���?`;����[P��\�q3�x�\�����qr�����}���z�uyZ��^繊G�)f:7�-?M.%��zT���̝����R�<$l��Q��ۅI?�p����J��F/�������L��\�bg8�G}ů ޣniX�
�%{���Xv�0%U";b�~�F��8S�	���"���n��Y�io���s�ٗ�bl���U\<jM��@x��~��z��["�9֭i��ü@'ҫ!�?��k�
�[W#s�������n�/;��-���ʭs3�����=l���9�~���q�~9hV =QVG��򢄋X�ǋ,�T����k7瑛9�h��\���\�yP��y��G3:��FŒ�Ml¿{��$R�R����kK��Pt�[�������q����-i��w����B���I{�RB'Ԉ �%��m���w>���,kT��2��4H&_�2Tz�V�ߧ��٣�mȅ��5���x42}��b�(�"�M����^n8�o7VCx̧��q7u239�nM{M�`g�Â����JfV�^
,�goa1<Px��3�2���PM�j���y�v}���/,�דɉ������OeZ����m� ��7W�����o4���(;�z�6ن� 6#.�X��@� |ܯ����o��xt<�vq/��!r:��X8cq̮?��ul������W�t}�Cߥ{}�P����mo����%]Ay��ֈ��h�8pg~�A����+��n4��'In1�u���,��TB��_ߡ:�ֻ=�y��+f|���oK5�gt2���W�Ta���r@����A�5��t�ʙ
���߁+R`���Z&p��г;��S�vg��Q}���W�k��_����z4��F��Vg��7k�L7t���3r�!ۇ��b�1_͝�f�5�п��7��X�: ������aULb]��p��s��D�&�Y�S0ͧN�����y���u����7l�H��{��?���{�:\'��uFk�[���n=��Ͷ���)����Z�-����{o`�y]��aff�F4bf�2�1�(��4i��6������%iNC��8�e��#������[��&j����;��й������k��kՔ�Wo��c"B���	�Zf�u^����8e3� ݷS�����4���1KOM�/��_���z�f�Sv�w36���y��0�8��*Pfɢ#�����)���h������o����gu2L�_���Q��~��&��DN�>(h2� �K�,����H�.�E<��A�o���t"��SO����M)��n*�v��yY�
��(ϚYB/��:[�Ch+)ʧ?�LX�eA��z�ͨ�!:�hz<B1��;2�7͈�7{�r�i��&��P�57�`@�n�M]�j�F;|����������3m�ʼ���G1lɴ=̾wt��36�u3&:5�X�uv׻ߺ{�Y�<��G�5��}y�q���Db"��C�P���8\�J�s����N3]���m������0s��0_GФW�.@�R��'N�D�5G�����Oϝ[��K�s�݉���+��x"�X�G�����2)Q)���&@}��7��u5�Q(֦G�Mh=��\��G>Bj)�g�"����@-e�ʖ������K/���2\��`;ds u͗K�%��D���,:-9��<�j��dC�uK*5V{o��=uƲrl�.����C��K�@|��ev�u[-'.Q��ڸ�ʘ��?�!���z��Q��΢=l��u[ڭ�� 4�2� \_@�c���J���TgW��9�9 ���)CG�F6��#C,�����+��#%%��[�X/�Sx@����y��3������F���ZC��P��O��ck�:�Q����ag�@N��|���δ���1k��{�{�e���س�u��T1�=a��� ­�tx��d[W�u��XwG��w�ؼ%� �~�݋�^���CxF�����!�����jC=�ɍX����6ˢ'��S��knB����qK��t�bK����y븯��A�˿�k�f��BUҰ���g�&�ZY|j���!���3��tF�C���tc�3]Z�x��\�Q�����y�	z�T��^����������޵��6��l>>os��?���O]D�(����xWf��� �(�����-Zhd�b���F��e ո��	��dע�̸��K���ޮ6 ���u ��q+[�֍�	�y��z�C�����ʘ)ԣ`�wQ�W����t��ed���ɜ{��MI��.F��d��Mo�w�!?��ʴO�#�i ��,�^hx�E�.O����|�kVP4�&pqS�����?�!3�!\%�Mk��{�	�ìs�c���@(��鲺@\��Knoy���R͋��ݎ�ʍq�1�"��VD�+ŽQ����x�#Pu�r�W��w
̥W.��I�L�v)�	��R����.#����W^|ޮ�j��߽��X��KƝ�+�g�	��=���c�leROGHE��	��|�9'#`6dVcP���`�m��.?s���(_��{��}�TZZZ�\**u���b�N��x$Y��U˗Zvf���۪K���Y���)�a�M�\`����#����dJ�f?����O~�ۼq�#�C�����]��[9��s-��O�9,v���9z���1�K`�
�$�<Y�r��oܴf���c�����?�������M?��? <W	�$s�K/\�����"�I��v;mk)��d&w�tk���T����G���z΢Ŷb�KIK�¼;qp^���v��!Ғnم����)�Gٶ'�`|����R\|� mD������������vt� �QX�Ƣ�V�,��8Lw�啐������m�'�"��g[jB��j�O�<�����1��gϞ��!���>�ܚ�y����r۸a��A�Sf���kG�u��������/ ��ｴD��Tru�)ΧQ?z�߹b��ކ�|ٟ��e�����#�0L�SO>�}�ڥ�Se��~w��a�!���/:0���2�ٳf�HV��a2Ȕ/�oA�ث+��/�f��)/���"�m庫�b]b3��{a������n� �TYxv�Ŧd ©�c�6F���3��O_\�!Ueε��´���q�~;v���%��j{G��9�ŷQ��Q\h�����l�d��c�P�x%��H@��^���O�?��?[*��'�*Ĕ�_��F)�w�7ْ������	ޏ��+\���}:3�X�<޻a�B�뇜'�[����d bf������kV�i�.ܻ�~�>e>>�#}=�a=�/�[��3��3���S'�C(���5N	�J�]�]����f�k����o����߳9߂!��gfX�v��g�@��\yz�=��]l�ɒ �f�_y�K�Ō���ÃA�H��Qq��3OX����^�r%�`��dw���N�>	��~G0ӵ�7�f�ZvV�E���A
��b��Sl���Pz�O���#��4��t�c�##Ӿ�l���w��CO���s/�l/>�,"9Q6���������쇓��Q2�NI�p?A���Hpd�C<�a*
A�/�����_�#�o}��Jq�3���>>^ښ[R�я~L�x��[C�@K�L��*[����j.������r���í�������C;U~ʒ ���x�hmB�l��(=�^��`��ut�2x^!/��If��Y��w��}B<@����?�|l.o�+mw��J�.�s�F�5!>��62�QF�N�x_��Y�-[�ܒ�=xx��K�?����Q�{q	р~�]IO�Lu-�z�K�B-������6g�r{��Se8�f��0�	�Bp��)����gTm*�&IS�|?s��h�����xZ� �����J��-F�]�`������/�O��uE>C�����[��"���[J�W4�>*����?�m۶96���Yو�`o�mi��%�F����l���Μ<j?��Om	��)��"�i/\�؊���8/ˆ����Η-����2��,��[^|�)e�����<�q�i��02��G�phjj��m(�EX,��	�[L��Ѳ��f��d����.��s��<]��9����@�o���V~⨽�� �I2pHpє��P�k�}��h٩18�-wv�-,LF)�D�`J���|#,�tdm���Wv�=��^�z)�#��s	ƌa����Ą��nڴ�j��?+��_��_���������l:x��N�8�Q��2r͘��T�R}s�k��}���I2���<۲q:*#X�VC����3Ӣɚ�����~f�����W��l���6>�[�V�`�n��-Z��"R�iY�@�B��=��қo�Ax����}�JA(����F������l<�!��̙r7��r�
+�Qj����l<�*Ϝl ���f��os-p��z�y���ȓ�X,z����{�=d�,�V���N��m/���N�}��b{�79��ۿAi�љ?��{bJ�8ǌq���̥�����~k�����?�?����G�G����y��M����"�iFZ�����5���o���D,x�~w�]���<�N�.[dU����8�D(��6�VQ���/���� �xz����75�Zv���m�`�j�F�<Iۆ�kyy�+�ϛ7�{���22"�ƀz���`&M�XHl�敺���cǎ[Y����K��	˜{jnpķ�$��� �	b�gIX�>��v��5FUa��$B7��	���Nn�L��߹�U����v���Wn���{�".c(έ�w��wQ���9���}g~~�'�Ι�������������L��\����7m�m�Ğp	#K7F����w�(@Wv�N:�V�f��Ͳ$�T������ʵ�lƌ��j+�9�,>�F{Zm���Y*���c�-#�؍�e0�����ȯNA�� 4W�`�K>�y2����-�|e!@�=
�Rͧ��' �*��f��O��J�h3Ќ_�d�]s�5	i�Q�A��S�-19��$g��W�%�c��
���;x`�]�a���:�)Dc&�G$f�Wf�?�ɏ�ܲYv��[�������H+�Q��n4��$:���(�d����O�W̙3���?��s�W�#�#�" �<y��/���}��h�,���z�;r�ɨNR��,I�ȡ��Q�Ύ6[�0��5� �2 Nd�)��H�l%��x��K�0Hɣ�=d���y��eRƎ����+�w!�
����Z,������/��،�M���B@�%Ԫ�OYbb�k([Wo<�4����S�+<�q\�q^�i���͛�`�+c�<�R{��eɴ���GĦ�G[���������NO�\�y���0A�<��Z�o㈾��J_�k���jˀ(�Dg�W�d���&��)�[a��6��3������-]tUA~����h�.oC<��A����x� ����ϟ�8}���Ť�%Ϥ�	@����_�=un���e�!���Z���C6����ɧmN�"���l�B�5��D;yx��Ua�(*�N��<#���u��Df�_p3�HƎ��3N��2����}ϕ	;C�PV�xM,e�=�v��4ܛ�x�8S��M>2�i�p�\+�Yh�����eQmW\{�-]��
�CW�^�Wo?<2�֬�d�2�a��}6Ie@��V�c##� �����N�.����d�^d����g��Æ�mظ���ڿ�i��!eN��X�}�r�[+W��*33���?9�7+�߬������i�y����L�`m*�޳��^���v�l1�����,��aH��&�ن5K���	z��h�gς�Vh7_e%��fӫn�=۷CtK��>h!�س�'>.�r}����D�琦Q�H���%$ �o7�o8���\*p�Tb�AI�䩣�˵H]��#G�Jg�{Y��_roKԷ[Lbs�ef�|��2]�9�� �����[��n���t{������ٕ��)�w��:Mu��M����@L"�
��{zz������>������vez�+�{��ziS��5k>���t��v�F���.�G�/�G�G��E���f��c������k@"�I�����e�mh�O��&��3a�0�W�]��8Yq}�% �����"(	PG�������:�����FO�FFG��ž��;��|�sSkB����Z[�Q��w<�fw���bB>��������:0>>���󖸸�WQq��y2^�}�w��������TS��ۖ��Yn�L�m-M�B�k�-b�l��=>6e���#�w����ئ�k���dr��f�|�H�Qf�����j�z�ַ����f�o3��=�_��e��7`Į��}ϟ^}��_�ċ#�/����Gಏ @��#�|g�����аX���S���c��B��VV����V�����ʰ�C�x�|{���-�~wf�6dUU��3�
l����� w��vc}z��N|�m-�7�[.e#�q56ֱh8�2�\YF)w����N_^��Q���T۳g�����1��3Wy�Ё���+�����_��/�ؑ�Z��,N������\�O4xS>����ڝ�8@�NF0"�!g���A�=)-���c��G#��X�}���0������������T	��u[��
��~�#4쓪��/@���e������"zX�R}.��������OL2Fzn�\`.�uٞp�ؕwt����X��Ԕd[�b��D�^`�7�w`��rfZ<�/� 5���"(�Ϟ�؆Ƃ,6*�BǇ�ڛ0I�'+o�EKV:9W��N���n����~�_���>��.��N�,G���N�8�LN�q`���MV\�k��Z��*��DS}���w?�҆�� ��%���Tׁ�]s���m
=�	�_��/�L9�Ȫ���~�����T�:�z�k���L_���¨z�T/.Z�Zǎ�tNi��v�kOlC�~��?��|`����.����xﾇ~1>5�>�Y:���z�3ա��B�F*�@����Ef^�x��iʮ�re����`%-΢��2e�d�OQZN%{-(�cpЭd�Bˢo�C\�2GQKI�u�-!h�'�f���N����/��@����c���# �j�[^��D_�˫-,$9�I����I�|��ѵ6$d�-�~����XIq��]�<q��;̢�S�_Od�,��� f�8.1�i��;��I��W�/?r�6�߀�|�������Q����\�uq���E��\�QDc^��M���a��̗��s�c�Q��/��_��_�����/��>�>Ȩ�J^A"�ɾ��Yoɐ��^Y���Y�����fW�\���V����g�+���yҮ�d��h�m3�Z��BU
h�ن�j�h�w� ���Գ�w���
�fki�4�U�H�6I��Mٹ���2?}��M�Rg��lwYo�s9;��0#im�L�O��,&��$��{v[oG��()��y�hD1:&�3U������!8�u1{��M�MBr����@��2`˷RB�ƿ��E�LZ��bk��_=%Ϟ�5?����"Ʌ�����v��;v�u��>t�=w�{��>[��=z@����'�K />���8~�O�n���ӻV����9mJ�R.F_����]SȠ��֥�v�+��|�vՖ+�{��+��)x�wbڋ��$�����b��CGvD���P	C���r�1&B�$=i��[�[��@\�m*g��.�?�-55�Y�Je.���ֲx�p��3�����bQP`����dz��L��MX�9�=n�C�s�#�:���14��&X>d���.;�{O�[��G��;��=�;[n���i����+�P�?�Q̄c�뾮@FV�=�d�JKK������%𱹬o���/���o�G�@uU��g+*>��Ф�.�7�Ў?�V��Ȑ:��(i�UWm�to�d�%Ŕ���Yo��7�n�?�0 m)yH����f3JP��O���&{�Q�g�V2�IK�bl,9	��4ۿ{'��VW_���0�p�v-.��.�U�W�����a�h��ـ2$9<�ϔ����\Ӗ2;��J��bnU��G(D�1�M�=:^�r��y,b�k��4�b�s�"�5A�豣����@c>
s���O!�z��� ��Ļ�}ũS6�t������V��-[���C;{�l����?�����w�^�7g�M#����x�"p����?���l]hHH�c�J�p`>Z���HF�N�Q�#G��v�=w�a%��mG����P�dC�<���C�����,��.DWR!�EE�1�>���;^|
-�U����&��|l����u�e��Kw]Ү���E/e䒐=}��]e�f�2~���̊W���>UN����b��\�Jl�����ƹ���x�֦����۔�k�2�}��4��B$���);q�mX�yۧQ��r��Z	T
a˷6�Y.��q��5�؀4���̙k>���썷�z�.[���7������[n2��.�g+�=��s_'㼂Q�pY��W���2I�d�������cp6S�������z ��}����h���_f�(��'</;�*�0?q�%fdZ�F�0e�ʝ��k�ˬ���4�����?������pF;}�!����n�R�2u����M���dֻ�1�T��ғm��0���xu�E�$᎖�✶�2|v����6u��~~|4������dE�-(�Y�V�����	�g�łb
���Ǐ!`3�2��͑�%��&;��~CQ���/~!0���'������>�?��N|�~�<K'>m��z���G���
�B`���][S�H[��	�k KY�.D�5���([��J WC�)���PvfV{�f�-�n��]��z;�ء�6���@9=���0�P�k�.OMϵ��*�flm�X��ή^�\O����7�
�|�����d�]V�.{!L���S֌�y%Y�"�1m���#,�L���O��Q��{1|�m�������W�~vN�mZ�m
�G��0d��`!�x�2�&�{HH(F,,-3�`��#D3�bcdh�r

a���`=:�� ��Y3w��=��(��}��_����'����������֖�����Ӻ��wd9��5J��q'�� ��Po�|��b�����|�m6gV�ػB\�%Cx��.5���y�u�C<���%ӕ1TҤ׋�XGW��A SO<.��4�/��
|��τ�>���\����566I5 [U��c̩ϙ;���x�ǫ��"��H�����W[TR��ݳ�Z��dYɜ����a��Ak��b�EM�8t�����Z[am݃�n�&{��g�u��WU�^=ĭ���Syȇ_p������k��k����w�}�'b��T�ۥ_r�Ԟ����$X�<��OL�O(y稄-Y��Ԯ���oC��ev"�X@=�xY�8��@������&eV\:ۮ���-)��,"�Q�>p�ui�f� ���Y����+d���&Ƽ�X��EqG�u%t���z��"����ɢ�l��Yd�����)��%���e�b�r��a���l ���L�5�An���,�R�R��饋�w�6�Bb�ΝT�'`���j��Z��	l`Eċ��q�-�Tiб�����f�i(�Q�w��D������>���"��[\�/��A�o��x���^��:7�u�l&�<�5��l� -���ҙX��a�z@��9��M�P�>m�>;a�b."wܢe��ag��Z��+�P6��VS�3\����6�TfϞ���"(GsR@;���a�Z`h��U8^zF2��ю��������ft׮]v�}w�P�ę-�z��u�z�%��,i��Pޏ�Mr�r�Q�J�ZD�Mm�.����W󵝹�.�eU���Z��Hx�T�˟�c��E`��h��J�#�ϓP�C���=�xw��k�����?��_�O�_���%����?�̓O��6�[#]���5�-�x*#�@ ���q��0�.�o�z罌��V���wu8�w����P:���\b��!�t��<FǦ�����u=�z4�i*[bJ
jq)�#��n����3�)E52de�Ҁ�(�"�)c?~�$V���|�2�1�]�<@�6�q5���"߰�
[�r�͝;��A(�of�Y���	b� �]��s�s���uT(��T�>i؜9�H:�dށR���ĕ�ć蟫�>L�]�w�40�ch'��a����)�������y���?>>oY^��҇�=}����t�K��f�r����8Wy[Y�4���Rm��e�s�̶�~�s g>>�Kmjn%�
r�l�g(�W[rZ&Z�#X�ΰ��R$Ws,&��۞��n��;�B1eI��.���{��]g9��!�Qu-"�	ԕi+�mmme�{�	�h.� ��/��k.�E��#�Q��/Y���V:{��K�(�X�SM���5�V�bF@��������s&��RrW/��-xT9���`��G��h��-@$�*g6-LF�F������lw*�~�t#�Iq���w�#pAE`�Ν?t��_Sf���.0��]y���I�r2��'$X��OB>�,�xY/����r��k�I�$>�i����ÄovR��)�h�:��{������#�"C/�3G�����(e�VlR���3�d��aJ�2�0GXˣ����i�X�׆]�J��q��w������e'0`�EK~���v��>��sM�6!/1%͍�)c��
�(�fx�;�;~蠫<��,��n'K�ŏ2ܬ�E���݌͍:^����i�crg�5��켰���AL�0��L$���訃�׬�򖫯���a��D���VP�@�ڻR�>��;^��F��Y*W櫾t/%�3�����&,?/��{�ݔ���ԉ#6�,����1 j���w�� �����z��;�cܭ��4�Vo�b���K�M�m����\O�	��%�֑R�@�r�J��0��9�����a$m޼����"���:�vXhvۭ�1w��غ�j�U���`�iAz��d펴F�]:���k���U��ʳO�(cm����~���\W��U,�r=��By�����ғ?J;b�}8��D����0¼y8�q����>v��$^>�%���Y�;�x�#��S�}졟<���ԩ��^\\lEEE�:4��M�JCã����")g�`�r��t��ǰس���H�";��b�˞��������9���^��˰�d]��f�˞y짌�EX����(��,$p^t����ݕ�%������:�,{*s,��1��t��g�?�+ �۷�(��c���*�=o����g���e����$�W^�h����u7�̱Z��?<<�u�٫�_B�&�9��ADG���S�\ey���uka0��}� �߂!����͟?�{o��'|[#�Y�ok���}.��:v�����t�$�ب�~��A���E_���,���2�Hc����r2R-/#����a�=�����N�<�`;����#�'�Zs�)�����H�v[*B-����BU�E2ߍ�X}S�S�sNk�z��S'�A�+��v��^1�Ճ>u�8���ljw�t����^}��`�����я~l��O#!fų�l�M�ɣO�91���`��p���O�[x�UU���0��P�k�)u}��L��/p���E%�i �>�M_u�����,�����B'����q��\��.g�.���?>>oh���"����>�o�ߣ�, �LkOo�&�s�v��Jȣ��]��
�sPz;cMșΞ9�2Rɦz���ed�[���Q@��%%��0�N��ZyI�ȱ�yK(��N{x���r	Ҩ�j����N7�݊^{,���'�M�r��O˸��qt�E<�����������M��:��}�X'�O���7ٜ�K��������SC:f �u'���*�K����W����Vn������\�H_�4Cf<wG��^�=U.�a�˜F�����6L+c�8._��ἂ�G�\}�w�Ї�vQD��E��E�\x��'?TSQ�Q�v�2[e��O�޴��23�01�5����rr4ٮ����]w�E&\j�����%G1+�
.!ah�3�+17)Ĉ�l<5�Rz���'��ִ�g p���9����{C�p,"��{i+�˼�]CW{+�rփhMuM��}KbV�ًΟ?�������L�O��ǹ��6@�<z�sv�L���3,,4ڂ�RwTr =��t��\5"�r�1*��}�yb��i���=�أ��?�df��B�"�u���0��Q��gC8��U�Ha�N�gf}���<��_��֋���͈�Q����#p����N�8�� �l���Ff%{��E��%�.��kd+�q�%���/K���EȦ�����{���}�Y	�o�֯�^`�9)V{愝H����Ȇc-�Τ̭�G���S� ���W"���}���^ǭ�l K��9/99ٹ�I�N�.�r��2���\۸iF/��I�mϿD�>�8+�9�f�JHL�~�+WN�_߻|�2&͏oq��V3gO&]y��E������6�j���c��"D� -.��ׂ@U������u��L	İ3>���g���o�?v��ϋ������G�G�uG���������pvl0���r	���Ѻ�z��yoW��_��iV������|�f�ȇ��8��8@8-5ݮ��N|A!�٣���DZ��aǵ��l]*j��ƧF�����-]����ϡd������V�e�,9RZ�7cd��sr�\+ <"��U�jma�z�J{�ݷXtR��V�������۪u[ kdca�Kb5��^ni���'U%v��)-jȜ'�Fl�K�YY�|0��;պ��67�6��]*�^O�-��/KU��ջ�r���,^$����+Yץ˗�XP\���6���~�� }<)���|޾���E=���|���o��%RYww��\�lWY�����t0ni��ń���(}�R��G>B{x�v�؆+��c���3$l�^x�v�u7�Ɗ��c�%���^{��슫����f�B�-{?=�޾۶�Y@}��D�.>!59f�cb�~7�{��1�{��g�(F�%�Y#_��Uֻ>��=�І��7Za��ث��'`���Χ�u���ǭ�r����$�s	�hS�^w��_}�%[�|�=��6�ܧmS���W/�9��Z����pU4"�s?SE����|�M��rS|bR���	�g��"�K������#p�E���ۿ	@�C)8J��[�@H�1�K��I���]Z�#�¨Z؄;���#h�'��߮���c������=f�͵�L����k	��Ⱥ�I�������Hי��D/<ɢ�� ۾�y u
�3��@�?m��([R�w�����z$f�{��*]Y�l��`���cx��S�s,-��-���J]x8�14�o�d��`��J�=��:�C�v�9w��:;�]I~&z ���Z+Z���7�R�"��;��E�s=y#��mWl���/�0o����M�?�����榦��g+?�gϞ{�]��+ *//wB1*K>U /���K�Xټv��q�D,�����L������vŕ�;i���Qzֹ�Ek��~�j�Nۢ嫭��%�x���vF*��-����ϵ�Ɩ�9��L����gu�����,��"#��m �H��Mɽ@CN�B�<'�RW]�z֯��î��vd[��5+?�z�*��DL�a�����H0^�� � �0]��@��qcy�-Mr]��!���> ��V-�ci�^ /6�2�	�\��%��~�|Պ�=����_���^�=���������}���w��]����@�@I����v7G-@�����Ν5�����m�	��D����D���\:�� �Oo���F�RR�!���u ���u�ؚ��鑷�cO�}}��XZ����z[�f�d��MG���a�*�;���P��/#�����a�'��w +��qh����ۖ-W�a;����ۨ%pm�DG&Q^u�sXD�#�M�; �B�l�p�f%U[UQnUX�N0J6�*{�ǩJDrMC��G陧�i��Z�:��y*�W@���J�Е�O���q�]^�q�W/�ϝ���9���?����#�#p.0�������Z��W1��Qj�K�`�s� ���]@���� 0:%��N;z訓u�����.�_6߮��j2�4�\Ra�?���;2��A d:��E�)-59�v�-'�k^W����dBA�1n��W�mi=�xO72��:���Dt���rd3U��O�r{N^&e��V�`�˄_���M�[XT�-^�
�����r��"w���LO������=VP��gA�a��M�>a#�CΚuB-C��h���+ช�F�T�p�}�G�S<e���ɼE��9k�w<���������|��������>���yJBb)���%����J���k	�"�ur]-��AB����<##����6�h�]s��VI.�q��0��ط��V����1�1w)�.��)�������A���s�`�r2�&�o���vPb7��8n�1q.�Wv+�2���� �=M�b]?�����jmŊ�6o�KbAq��$g���ჶt�����ы��#pP�ޘ�;�9PN��E�D��_>@9>#3�ѻr���Cd��q �ء�6�t���%nf{"ew�ɩ2������a����cg%2��3�s.|�w?������w�l#�K���7�#��"Py�b��={>�*�H\	�&��k�Z}� �+�lGn�������Pb���M��bX�x�G0t��HdY9����ȚG-�>ttd��6kC��״��,��>8��Me�NJ�՘�0��;`�.r���a������^G<�����
�.a���L�^��(���]�Lx(�����!3۱����O��yWX�[n&ۏt���70>� ���G���ĘZpP8�6Uv��^u֩�쑇&��r�2s	�h�L�p�!tM"�)�@Y���m�������/�۸�����_���{]���~9?}�>�CZ[Z�y��')��IK�����R&�CZ� DLq����n�!m�R��F7�_g�\}D�;r|��1ge�̥�J���+�g9�3 �a��沆����[������~� �EP.�~_K5@��)ɩ e'���ʀ#��G-ʹ+HϮX���\ ��v�b����/���Z%v���$�� �����-�bA��`/D:z�-Ag}�*N��V�+ڠ�9��v�່�8qS첲�s����]��r���R�K`��ŘkQ9?19��?����R��_r�����\f�o���/�5Y�\���]*����\�ۚ��̥^z`X�vXTZ���K��z�%����x�U �^xA���������Z�e�XWw�zf�3�,����^�ǎ����J9��0���K����|�+��g���w�����,\�nҋ�X�5_�l�%%'86|
��ƺ&{��gm�-�@�-�f���IO֩ĕ�+���)�T+]��:��M,:XĴPh�G�h�$כ˽�6�[\t�����+�W���Bhz]Lv�����x�פg�?y��w~@��>u�v_O|��z����#p	F�l;�~��b���ݝ]��םi���X%v�677:2WGG�+/C�|���\��C��YR���}�8�y��p�m�F+���Q�����`��m�]������l����uw`�Ҁ~9r�(��ΙC���~y�57qnJ�*��]/y�n��ʴ�យ�>4�}�SUU	�׻6�G?�1�&��C8��V�ÞSdKVob�<�e�}���gC�M@�{wls͜KҖ���={pm��k��Oz�2X(�#R��{43�\s�zgk�{��*�k�a}�������а�����X��b.�[o�-y���a|��(�y��ç�9�y�� te���3�i����[��`�����	�i=zıǯ�v��s�]Kmݚ��s����(�cd�q6�����r���̃'YW[��:�ǲ(yw���@.5%�bm��A~%�A;p�0>��,GC�HF�����We����q]�v%�ZJ/�ܙ�x���7<.)Ֆ�Z�B\���,�O��>���x��U��ʄ��$c;�
����B &����m^�<Ǡ��0�>{�S���j�E�>���'z`$-``�yZ���x0����\`���{ �r|���޹��CB70cΈ6�(=��Ү�g��d���q ��`�6of�+&z�e0:���m� �t��i!����+mي5d�1���fG������(�EƧ0���Z�ׇP�67� S}��1H�� �2A�TSe1�WUUS^��0{�s��NfO�;	�2z�ʀ7n܈��+.)&K�1J�M�wz�U�j��)�7�:�	�k;�������F��A������x��L˵�S�HC�F������(�����2¦���"驷��_�4!\�T�\_>4��-W���Uk~�v>�;��~q??�>oH�}��?�����y���zi�����xf"-��L��55�P.������93!z5�"6`E9(���X�.{�TJ�[���ٟ�'%;��n2� /��<Hi"�ő��I��t=b1-]���s��0��(��>H�u`��?Y|�&����� �Y*u��U������
��;|䘝�����j�6]a��3Y�;�Ue˪<Lo���7'}v w�}�:��Ȯ��~�V��h/m��m�ki�Un�1���r�@��++�l{]]�����7�f���0'@��w���;R�ӟ����~C�?�eO��l��q��|����*�n�

W��R�z�/��2d�KJHr2�*O�^���3'O �!����k�}v��Q[�|��*;� �w�l� v@�����^� %�P�S]��i2���Kf�c̬��?�b�-T�b�ю��k�,
"���a g��g*�gM��F���Gvv::�e�E���^y��z�VK`nVY��f��ȏ7@/�r"�	�����v�ɤUߗ��(�o"��x�%3���c��{ �:_���7����\�T�}R�x���e����D-�Q�_:k���-\��,����E��4ǎ}��=P� tG̒�Db�h�LP'V���0=���'!�a��f�i�a�F���}br2����:
hd�ԫ��Q9����y�3f����6J�-诇E�3�VD���Tߺ �UQ�o�o���Q��F(ch�ԛoiid4�cki����6�^������S�\�_��|�J{�>b!ؒ67�ώ�izf�n��Y h���~dcwR��3���t;z�}�&Z�#������?�`M����.59X�X��kK"#離1$@G�ՙ����WPP�����33h���G��G���_�|.�`{��?���~�rp�2J��J�A�^]h���>�f�gϞ�q�|2�	z�mּ"���d�1v�����~�6L&��[l3�,�Դt�B=���Q@4&�~q���%$e2&����-?E�?x��79����#H�C�b7�
WVߠ���6$d#"� �B��Rɢ�b�����z5�z�j�*--e1a5gO;����"�MH'I�{�1�#��Ykmj)$�8�Oķf�|\B1#CNf����ϻѳ!U �	�UVW՚PL�#�����ݹ�q���w�wﺏ����������sA_�/�_Џ�_����q���R&N�b�����+���	�6��x�)} ��:��n�՜�����������?��?>��W]����bp��+�� �}��PT� �1��Hkw�qF'��[A&N`c�#Xx���p��[�ܕ���%��/�.2�d��5gOB|˲��lk�q-2&�ܠEs�����Y@H�u�sҔwJt���'%Z}n����$o�h���DY���Hr���Gĳ�{�V�\i3l����]�2 ��Iz�a�	��i���}�T��*&c,.����P�;z`����?C��L[1� &���Yޮ~��+�+�q���V~Kp`�4�u  s^IDAT�Ž	���Ě��?T:{ށ����񭍀/�����g��Oط{��/���_ �فq&�q���	�0���t����G����x���B$}��i��V����KV���+�'O���ԓO;<<4!Pƻ���w��:�F�4ť���t�N*)�7b�ky�VX�c7�x#��(�ŗ��E�-w�d��a6k��A�p����6�m-��tQ�O&��vr�q�Qᚭ�z73��	E �g����q�!,(�h&������螗�__�|1�sٶ}���qm�{�/]j��ǜ�|�sͼf�������ȹ�1n_��1�������F����Z�9S�T�F�̠:���W�|l73�����N���P��&;K^V�Q��5469�ve�z�;';�o��OfΚ}��3�x3"��͈�?���k����^�̫����	��=���@OWe�I�ָn��0��P�����6���v�l�E����l��{��cϿ�K��0߽{����-��W�p�m�RJnG��
��K�Ƞ'=�Y�9~����0�F���GR�^�f��[��p�b��&0=�g����^�9o ��j�s<��mw��:T��)���_��ъ�W�a�����G��������	��H� �]��:K?ew�~��Z�����l=�3u,H�����r�ৰ;톅�@i����L���ô?������~�s�	H�vsf��9
����F�b�b@/��_߀|8��	���� �)��� [�x��+V|�l���^�����#�[G��o:�F��.���<���N���ӽ[}x��HS��|��� ��|�ۆ�+lΜ2�L���(�����ھ�d��#�c��42��?��#��)���f��ߑ�T^N�Y�����**�QT�q��~7	�\�ʖ�\f��`k�:7#�k�j�9�v^a	��Ռ��[<�iL镋�.R]q�F��!-���;��9Qz�b^]Ҩ0�]�����K�\�����gT-/�R}R�$'.ӊ7�i@=1���ۿ���M,L��0T�m>c�|�x�v�q+���e����'11ѵ��8Ո}/�` xbz*Nk�������f��_2c��<u���M8��ɻ�&~�������	��������G����j~�O����k��'Ž�X�=}^w����������h�9 �@�@`���@cZv5P��n�5e+�-���\���xMN[d ������dWOG�5}��+�|�ǂ'��cb��7�͚���*b1�ۛ a�
6c�,�G���Z8���
k#�|��w����'���p(+�̬T�r!��-:&P��g�H�&�7�HKt�! C)����@/���U�P����r2r��[���'|ˣ�f��lA�e�������CI>..��8�6n^C�|�+���} u7f��X8�"X��x��,,��X�9 ���"�5����>�⡇ED/d�Q�:sR\�[dDq_�Ȼ��V�R\��i����������-���:��15-�F�F{֬]�w�_�?��O�{�������ե>�����-�hK 3W �l35��$V�5+c��Rsb|��2�l�u��Rvd��ԝu��8��(/�bmْ���lꩈ�8���<)+3>6E�?���_��!a��kI�z�`����eU0�s���uQA�ER���gm��g�'Fm��E�t�l �������E��+��JJj���d��ǎYfv َ�M�@�K��X���sB+�1W|�x,#q"�e�����wҫ�1y�=g��<s�k�BV6�Y�v ���VBf�]�	e��B�\�@ܽ������Y�lߑ#�Ճ8�(�7���sh�'L���_�{��؈�1��磅���X�
)@������.[������|�*���z���������k���Gා v��~�� ⹡dx����������8���3�}>+��8Ǯ��*k��+55͕����\ƨQ/e��Eh�z�v��e;w챪J�őX���L�"���̛ױ@��y�Z�z�-�?�*�OX
�뙀<c���ǂ!^2c�-\�����<j+�#�<̋g����Ȇ;*�1�VO���yHtǉ�~�S��[ ��l��[�5���\��;��~Zz3婎Ů*šC�a����̟X*v��X(�bV|fq�%g�b�r�e^s���^KH��^�p��۔a7V����O�����68neK��3O<a/ԕ�EB��QU[��j����X���d�}�49�9ͼ�Ңq6U&)�oذ�_n���?��?-��>�]|����Ϳ�G�5G`��]w���~�Rs��'�|ɒ#(;\)�W�2J��i�N@��I�t��56�]�Ď������ �(Ǌ@EM�,e�cӳԓ�d�h��_��r23���Yp�5��櫣!���yE��{ u���[W��f���{�}/2��%�f�f���M:6�A�g�6lFݭ�,6�
 qg�:^k��ﴂ�9\
l��ҙ�4�Ҏ8ٯ�X���(�y�%1�1Lo��e�,�:\|�<'�:kV��Uu�1��~���߷ x$�j�}�h�bW���	�<���Fqv�i����,�f9��&�s/���Q����u�;���	I�9%<1�!�UU�@��Jz�!����{-@�!�c ~C�`��Ϙ1��_�?���op@��|Ώ Jlk~衯Rލ%��M�mʩ��L
8�}�8�(�uɑʲӑ�& \@�o5s�z�BKJ���/4.�ym�;(��-�1e�a����|�)ǰ��U1���o�'�|���d?y�%�bHB�>�|'�Ry��EOp�,Ho#�<o7^w%�Q���]\0�z�Q�} �;vh�-([j�,�B07I�T�t*cK�&�y�!@�5�� 8��#���[�{)��vQ�~r��>����!�쌵��3�����yI����V��f�+���e�l��U�P[Nܢ,�97�Z@�(N� ������`�c��5�v������㙝�
��tٻ*��H�n�փc�>t|��W�w�ˇ �S��%��
x�������#�vE���y��"d�3�̑	s�fd�#ί[ �ްJ�#��w��P2�Q&F����Η,[b�sˬ����T�:k[�;�n(ۻ8 }z�pZ�j_GȖ3졟>��0��,��
�6�<�TO���4�e�z����k���.Kf&���.�Oƽ{�6[�x�5�5�^w�7��SuЈYVf�v�f���8�o���=���SG6^:��f�̲�8��"�j-�p/����Z�̊f[s�+�����Xk[��L-��#0��g~�~{v�/?Sn� ��8�M�K�N3���ek6�x��QN�*������[�뛖��r^2Nl�T��B��@����5%-u��}�ë.����:��~A?q{r��v�c��4,f��@��d��!��݋X�J�}�� _��8v��g{v��{v�7��_���S�^Q�%�5<��(��wD,�e:3����:}'�e�0g�����v�uW�4��b0�S�h�J�F�yV�l�3k6U�H+�g_s渍 ޱ�!�E��[:%�8�w�I�v���d�*�S�n�0�E���q*jb��ٳe�Qkl�12���#�Ĳ�a�@\#jA�z�/=�l�e�7�"�������k>g!1Y3}�R4��`o����h����qQ�볐�g�Lp�����\���Q�0QT:���ؙT�8��A��z����O/~�*��q�6F,�Q-AZ(p����ݷ�~��_�S��F<)��x��..�|�߿^K�D@1!��qHh��L<�)�VV(���>��������j̈́D�?���:����w�(j(�*�?w����~����a��B]fII��Ru�����o�}V�_b�)v�UWSV�B$�τh���zP@A�������-��?7�@���^Iɴ�7Gen��s'������1�5N��8M;}디8/=��>2�lG��>h^y��`�\�cU;9���z�����۬�a��ɤ�Wlr��,l�-�]P][��.^��_������5{�uصd�C}(�і���<�`�U"W�]��]��z.�T�8���'9\��C�QP�ŗ�ά_�z�/^��G�G�_�e��_f���[�̬�݁�Yg�f4,)9�n��fG:KMKF*�s�Y nRb�3 If͌K�,|jľ��_a,p�Xb(b�����wP�S֮�7p��@ &��͞gW_��f�23��[|t��zy�r�M�#�p�Ν��i�ŧ�A �G�3.�G:����R��]��5U����J4�������Q����Ow��'+(�C��Ϸd�]JK�-''ݵ����[~^�m�x�mX��
�:��>	裾m��E�%�9�������NJNt�n�G�^�<z0�?�/3�I��lq�2�0J���h~\�����V���*)�Q֮�iQ0]yqpdxræM�������������t�	�x�#����4�L��Kx�7�-��ag�j������g3�Z�x}c��3JaY� ����	7��o�;�t�S^Sg�|U��ec���<2���5��>��X}.Z��g:��I�q��k��{a���PO �0N�K�\�B#�{�Hׁ};1,��N�A��(XȊ����Ǐ��@��̼��G���Տ����Ȁ[�L�N`Gz�r�M/b�״k���{�p����/R�N�ܒyh�/��sf!�:��!�Z�K)SF0F�x {�E���ébt;n�z��2�hi  g���<�Q:U��wS�hon�X��*��/���tUL4=�S4B5b�S�}�&	斕}o���O��x��8���7��f C?�rZW�b�(�}�?~h_�Ʒ���/��^p����#ۮ��D��4�p4k�ώ2ڌ9X��u���(�TÐ<���8M �U�7�_΁�+�S�� 7��ZzV��v�;-9-ǲ W�xge�#�J�݂�K �X��)�8T�4:vKQhtV�C���q���-u�P)ǹ�Q��s�j}��5Z& �b�mF�$-Ü*?�uQ1H΀�6f˖/`��!�UT��Q�;s������B؋��iY�X	�	E�͋������OۙÇ���n�)kF�Fb0�Ξ�`�>��:�n�¡A---��<U�] N�.&���&0����{�T�����C�����'���#��D���ߚ8��\����	�hk_���5��������PȠ\�:02?>1�#�/�Db�(�E�Пn�&Q6�`�J��n�����/Xb��ٱ��-�Rx~~.��`c��WW���5i���� ����8����9a�����]�X�����Ҁ>����4�w�.+��s��^�y��ž�ABu�u���Q��456�VH�N?[��h�K����^	̐y��10��5�~��1G�S�A�8�ROF"���y'�x��P�?z�(܁>ˢrp�=�u�����X[
Jp!� s�X�Na����rkc|���ުʱp� Muy��~u�q~���f'N�;[�v�j�(���i���s�C�|��:59�6J��=�����⢟$&��f��K�#�o�������K��#�ҋ/}dϞ���&�ÈTD 8������	� p�9���2K8f�m�͞Uh����m���i��(T4:�v�M�Z������8eYi�d�R������o�:4�Q���7���uZ~��;�~��9�4.!P���s����鞌F{:����s ��9� �>@=�)�56�0�^��i"+��x�]u ��~�O�\c_r'�5�G���� 8v���V�UKW��>�I���ށ�	��V@>�����0�0סc�Q���?%/s��]�«<<2������0�S �5���>4�56���#��m�y�	z�b��,-uw�k���J�K=?7?��?��n��?���|�\��||~�=�<�{��/�N/�"r�����g��6�!�Qe��y(e㡮6�W:ˮ�z�7���h��o���fٜ�E�pPC�mﮝ�����@�
F,%�9�(t�s�'����[$5���H�w����~v^�l�܏�̛7vw�+�geeS@���2�O�����[eT+�"�c �E:�-
����l+�u��dXRSSs�`��d�*�Y�l��Z[�n5���pO��zjf�� �W���E ��蜈s"��@N;C����0����	���u�nښ����O�vb=�Qb��B�+��K��Ő�\S���J#��L�efg���w��������x�"�3��+���e:�:R}���0Z� Pe��Yo@�E��j^�D_C��k�jd����f��>ā�����̤w5�u�O���q�2��Zw���w>h��m&�lE�-� ��P�G~�V��W����(�|�8�to}z�*��;&�����+�UV���E_=�t�!�[a1%~2[9��0;߈�� �������W��P��}��t%wI�
 e7��y07z�=�E��1��FI��U����t���nJ���eDӋ�|<��`ٸ�iN�*ZM��r�=,d���m��sY=�̳Ki~d����)��vW�oE��߸��2����^0%x-@Tzwz��λ��Lɬ�o�fd���7��">C�(���!-M�9?�Ƀ/
̕��[Tؠ����.Zjn�Q&9���7o�՛ָlS��NZG�	@(>!�Jf�:���������i�;w�#?yo�
�=w=�t�ސ�N����%�,V��	P���}z��NNI��K��Mކ	L+���L<
o!SNDF#p'NT�mO�_d��r4��a�H�Jmm�E��˔���Uf�]�XX?���JfX���p�X^~�j����'tU� �wZdO�v��{ײ`���X�4`3ž�\սi�$��f��������`�KO_#ib�k>��*�3�c+7l�+�¿:�I<��&���^�8�g߻�����1���a�J�)��)	�H�]�4�$���h��y/@4�g���*��N�<e��p��=ŷ;4��o�Xa��v��w����nE3��i��b�>�c;|`���nm���͆��IU]��c>*p~�BAҥ�t �s���,Y��5�1k�M}i�ZQyM]V��)ɫ�ב�'�TF+ܞ�֦�q�©M�.r[x�`���[��A�;�T-xN@�Bo��VX��.�R�"��}	�9�)�6{�j[�j#��9/�:�$�����v�uc,rBXh�Pf�fl�g��{���&�E F��>��e�� #K��=���:�d�n�x ^���@� d9f䣘i�<����
��
;q͍7������o����/�_ԏ�_����斌��|�;�mm�ʞT�����g�x��^@��t�@;ī<�r�f�R��������DϽ'�H��9�)��T�f���"��'�6� ��+����-���hsJrlъyV�JZ?�9i���|u"�.���p:�4�]Ǟ^���-:������L�,�(=�8f��([�S_}i����v�l��ɺ�;�k*��m̃�⿞��c7�x�#�ձ�8ӽ����R{�����G��n��\҂Y\L2&�������3 8)ף�^���o�i?<�أG/	�q�or?�=�~y�w�_�O�P�SZ#׫{Vy]���3�`�,:{�5��V���>݈����Eo�r�=0�om���o��$��TJ��$� W?ׁ1�gf�����~��$�>�/�k7��:ڿSd�b��Ht�U����1%�"E2��T����W߲�Z�m=�^�R�"����6�G��n�Ŕ��/�������2yYp��c
s.������l���f�$��-�-�e�}��R:ǅ�ch1��PZO��^YQ�G1"v�L�s9�!��ޫ��d�Q�-jU�%V:����vd�NJ�i̛�69=�Xz�Q����sm!�h�A�@����L��1���m�>gR�����!I�I���T������_q�`L ��9�3_qF+��\�jJ������`��|.�����������x��g?En8W �MV*��2斖fg�WGG;�gƻD �%�1��Q捌�3�m�7���m�^9�W��W����4��EmډM�j�ăPEKJ�d�9�Q��auM�ۑ�Zs�>��rUE
5�^{�#���$%#ݍ��[�h�� �§�~����L��C�}�5׸��ꁊ��������p=l]���1�7�����,de{��v^��IVT���Z�+,�4���'~� �������z�n>U��ޑ�{'8���V7n�a����{T*?�(���Ւ�}����>�h[@�U�8ݟ~�z��_��닖-���q��x�#�3�7=��k0�h��h�hL@�HL�C�9PvY5e[���{�@�Y��NN~ϐS���)g_e�?mt�F��/��=yN��Z2֟��H�}����)J��;x�N��v�d5#`�v���?�����-���1�#�����=�Z�� �;�t�R{�'��)�Q����RRUboл����y�,77q�BG��rY���O� ��C���~x|R���x�*}�Pe�E��gD���l,�x'Oق�k8�K,+T��Ã��g�N�vB;=,��zf�UbWl�to���"��M���e��^�-,���-[��b�����8?����G࿉@JJʉ0���:4cg���
@�:FM���@oZ�t�ݢ(��ѫM�vt��Gыv�ss��Y���N�>��*k�^���%c���=n3f.�f�������}�������C�7��lŹօ�&"��T ����Ano�ٸ���&f����@�0었���u�\]��~���-!1�

�T����:F�*��[��[R�IJ�ݻ��s���[XL�� 몙t��'�����:r�6F�#��hX����Bd�����TB`�+.���3s����~1�Y|�M�.-Bt��*C�B�����5k������7�����_r������74i)���b�5�<�Ƨ �M���j��^8�m��'�%�v���0�& q�e��فC�m`lآE�w�d裔�Ce���4Gm��.�NG�R���9z@�.ax�'�{I�xװq�6
���P�
��'lr���9�|�h�諷�<L�L�*	a\%�����y�No���^!R�S��zՁH]����v��W�'O�f��H-.�G>��.�c��@ܛ�=^A�5�bqu��h�]��f[�%j��I�n�녠��X����������.F��[��*�A�%����_a�4jm��h�G������$?wp�A�g�E��om��GØ�`F�$�����I�������v�}o���G�����!�K�0#3N�~�ewr�"Cws�ʙ�5c�/��42��h}/F���{@�v�/��0AMǓ��4u�<	���]sM.kV������}�_�j�����-^j]C��i;wd�Z��  ���q7�-F�(�s����l��.Ҁ�8���OFqQ�붺rzkk�ˆ��s�:2�9��8V�SO<�A�0���I����\�?W	p/Q��6<0�B��^���d;^}���U�§���U��o�M�~�����e_i�k����]݃�ܴy��\{�}���*5#}z'��\B�%�K�a�[y�#����#�p�s5S-���Ą���ǿ*q��/8*#Uf�w�^[�f����X�e��J��#�iU�_���B��4Ӈ&�����h���=c_��XN��؛���_g7�t=L�*7��vu�� H�la��0]�� �b ��u��o���4�r�άE����O�ܟñ������,�ت� ��F�BhO��m�QF	�-^���>��d���d�R�Z��2IQu@/]��͎?�2p��z��^����"ao�shє��x�[n�����#�\8����,��\����z����Wh��P`PCwT���yjܪ	�Jĉ����Q��<�����K�q�Ў07��20G�[���x�1��TcBR�ˈ��1�ێ۫/���|�v�}��q���k�dx��M�-�PEph~N����1�u��%`�X�����+��,�B1� ���Z�f�n�]w�mV�HY�q�&pk�q���������!�a3�C�\?��C��CY��M_q��b��C`��P��Q@VV��r�sR�T��!�E��
, ��,_�����/�G����74��`�Z�s��`�8?#���e���ڹ10�[�R���D%x)��ٵ����ux2�8qvڧ�%9	��&x���g�ڭ���~�w���e6`���'O�����;v"�ڏ�JV����CI΁�z�R�;'*`�������1*�/���jٙ�v���e	�y��A�:%�dgL��6�TG@�r���U���>�e*@}��	kb$p�J49f����\�-��wy6���4}�8���$2�)@�S��z��r_�v��?���k=��&�-��E_r�(���2.�t������Ӟ��t�0e�!ܿb�)�UL�o11��_m�U�W<��t�����h����{��vٹ���[kϨ���A6����OQ~����m��s���4+,̳]����m�W��Z|�s�!�;c}���@�! �E���g�VU�����*DGg/niI��}��a�����x\#[��� ����J�*ѷ#嚐��f���[胈_uU�͘i�v���s�3��]�@<`ݪ�����b���o���w߆����o�gş�G�팀������s_�=w֣�Q�J�%�*MW�$%c)��DYb/�ð�{�������5X��#VQ~�k��#���k�v��k���A�����b�#l�z��[�Ț�ZL�0g��V
=l�Q���ŵ�xlI��s���=�������e�V�����ZjN�����6H,�p��`���&�1�5�c?�߇�j&�޿��[W���%�-��Bp( �lZ�S��6�qգ�t�w6����~b��z���d���/X��ڻz�'X�h���b��C(��pt�G�i�ƨ��c���`g�Ai�����S0ك����<�������/����70��P�nrrs��m`��EL&��Jll4���`����cV�P�JT*n���˼��Ҥ'���r{���e˰f���6e���.���� Q̂\_;�Ӷ�f��)��2,;�Yt ׋j���%�=~� js5[��h$@Y�lL�v��i�^�>��_�W2��Rx�`ft1�|� ��>��e����m�I��7��vSb��C]D��3���ҿ��v�jwB1��G{1�%��\���l� �x�2W�O;��F9�8a�����v�m��t?���|~}<��O���k�@QQ�*�j� 9L�1���G� _��նG���G1���绱�>�a�z�]�����%WY%��m��,�`��G�q}������ ����RC��c|b���^�ׯ}�>��/9����4��4��������y�R����������*��1����]� 	�D�b�#�@8���c'�!?g�*`{}`ֈ�8����UUR�cv�Nq ��;�Y�>�>:~@��1����<�%>�1��&2�^w�{����������������X�.>�T<�_R���̛������hw��8��l%���Yqq��t���w�k�6mr�we�R�S����Pj�$�����,43;��A���Fߜ�����:�<�� ��[�g�WI�j�+!.ۢ��mf�j��I��/���ؽ�N"ת6A0�y�������\]����s֪N��-����2:";��]i������y�rz��>D�AJ��!���7�/>��̀	/7��i��j=~��_]|y���Ϯ
��Q?ku��ܱ����a�=/?��ظX��f�#�ǽ�#���D�/�,_��Ϣ���ϷU�.0W.&yhH�3T���Gp%�!O1$���'&F�7a��nQx���@g���_�:�=S� u���P	�4��y���Y_��@� �"q�ϛiC�_u�,E[�?o��Gw�~T�~��v���������C�������xF���	LG��|է����&kX�����(�7ک��)��ƫ� 1�'Xl� X~��ud����]&��=�"S�?8�*\?e�75�.�!�BI,�>b(�K�D8D5�f�F��.Y�����nMLJ������e������G���h'=���+�)�ǐ����B��7�C�������e{��� �u���k�n�������R�9I��#� !n�sOz�h�g��ɞ�#�,��ue�[P��b3��@��c���=�����Jf"�:/ݲ�`��LY^^��S��b,,#=������W 7m�12x��O���݁L]ՁQ��#���'�jpi�������(�yZd��~�T�[T��F	�঴OF~��q��P��e���K^#|�QF����1�U^ל��uk��'��������%%� ��7��;�^g�򎉿{��6����;��J�*GK����D.��nz�À�������;F&QRXK�%��ّ���G�t�,�	���f6}ݦ-6�XW'����t�!��,�(J[=�ɞ:w7G��Vr��
u*�+��s�z���°������߾Ay=Ζ,Y�n:=o@��{R�{i��q�++��(ZZ�n�"#8�;�\��0)#֊@MsK�����t�bj�̌��X܀a2hG�������b�|�&����8 2nic��c!��ϰf��X'�nA�_P��\B<m�5_���u�ME������ʌ���6���LI��G�G�E��������^�s�{<ɣ �$�D5->A�-Sȗ*�MGO<�bk��i����N��n����Vq��E�.opY��߹���\	_�Y�χz��,��sR��9զl\����uk�!�P̓g�ㆆ�LhH�o6]k'��v��Gi���,�\��6;a��:u��rr�|H4b�����'�]]m�;��J�n��|=$�k�k�����ykc��ų��E�(�ty��VV jk�rF�cؠ6�_=�AX���6:��Cx�Kw������:�1c��_y����.��3���|"�3���Y�;}"096��cO4���%�D���&f�a�O1�օz*}^e���Ϣ��''q[�t^RTd)��$%$YɌ<�ю��bB3�S+#M�ʵ9��XuE�)]6�t&��x���O��ϕ��e����SS�^��O /y���LП�����u�ޗ�������̸�2���T�����`�!�iA�F?�E��񚪳0�O��-�p�R�6�6k�'>�h��
��8r�[��L�MV_�c[e]���1)(��r-d���n�Σ'A#j=���`Ѣ=[�����¢o������"���.�G�o�͊��}����O�z�I�������8g�|��1Wj~�w`5��ƸZ[�A@����v4����p�B�E��С��Sx�46�\ds��G���L}4˙��<�6wY�y��{��qо�PE��N�x�sgB�+�5��hL0�qؾ������mgq��8��쳶j�&��݆ �0�Μ���͒s�l���zk�a���fS�DP��'11��!���
Er�*�ǰ`�j�t�0�uu�2�L/0$��J�jH�mr|rrn�ܿ�`�f}��q/�x@�����7=�?����}�,��AN�D��J�7i�t�x0�g��xlj2^����-�����}�m}��3+��t�=��������[��k���N�&׬>2n-S��D����%���֝�q�0���7�f(�p@�]A��jr��L���X���v�uWZg�b;��xuu%"8-���$�^}�:q����|Hm���6ڶ#�����>k��3��ۙc'-x�,O���(#62jѬ���z�[p;��A��F,����&i�9]{ݟ�|
�2y�-�i�N,�e��}��?y��?���E_r������&gΜ�񩧞�\��@�Z�Tr��v�q�3[>�!�2���8��-����W�����f ���Z*-59 ������0۸�JlH�@�"�?n}؜�efZ:
l�W�r�ݍoi�<""�e��!���@�ߋ'p���{�rx7F(��pd�l�w����F�ҕk�y7[r|4I�Ho��C�?""ީ�M�(腉����Kz�cVSYmad���ߍ��M"#`����r��\��r=YxjoC\w|Z��Cxc��D s�H��D�3-�{zX�Ϣ&6!�0W�C�������|k��?������_���_�[��ں���W�EP��kMM5���>��ىc�!~���7�b����(V�t�����}j��~�ӟ��}�V��y��U�6Y ��������V�0rI���%Hf��	>�x��k��}ʎ�s�? �Ǻ�4+G37�uM��z�+#v�3�Jmʹ�M��))�c��ۻ��f:"4G�����~��~�6k�hf����#&-r_rR<=�A;s��3D=lO��rT��9���7^&&���X@t[*q��
u�k�hm�tx�ع@~�{{���Y<�r֧��,Y�����o�c����$"�Y��c�7�FG��L��}�����/6�5f�ð��$D��QQ���(�ǑI�֣�ش�� #]!���n�Դ$[�n��] �3G2j{v�'��t)��I��f���XfF�=������A�]��9�0+?~Ԏ��mO��q��/r�����@� :�8H
rN�%c�5	������\��5��t�>-5��B@��w��&���>�IL�͘Qd���VCzƂu�\$�����@�~��L8�<��Pʗ����b���7�Ȟ�nU��b�ʹtyɀ�kz��ᬻ�\��z�t�"�6{xTĩ�+W|�~��x>�r�e[]5�8	.���-xA4�]���wo����ݡ����晙k~�|�:�N��{m_�C��^�/�^��uu�ϛ�W��wCs.���	A �1�(�ݚ��TR#����:&w��e$�"�skOE����Ă$ �h+XK	ZMSm[I���b6R���K�Mc$�1���DP�'&X,h86�?+ٚ���yź�#���M�����wI��-��̸�K�O�!��n�a�B���~H!�7P#kǷr~�o(Q��k�KI��4��/���\�u=���"��cS�G��q:�� �>�"�:)M�~q�(�Y�Q&�P������%я���N������D.��d��©H�ts�|w��/�Tj�� K�@d�y	y�֎3=
���}��E���M�������R8'��
"h�7�I�Ί��Z22�Gk����|�舚�p���'N=�q�`*������8v3S����t��m��5�5E��t�7��^�R^�b�*���;�C�e����X�	�������Y�H��a�&\v�Q��� _}���Lu��� �����/�5��?����ElO�B֔x�}&�ݵ�B2D8�������P�u�����gd���UD��?�m��`�93\g��9�NP�ɋ�؏���^F*�Uϡ�+������E�O��`��y���D��~�;��1�u���e���I� ��>D�RJS���5��%��ߗ�dl������U��I���)�K��J�W��M��7���[�Ե�5N~�����+�IC�F@{i��Z��=L�b�e,����L�ǁ:�Rn~5A�R��~ϓ�v��iV�����4=5�һ����4d=n�`���u�4�.s't���,��rZ��d��V$M�e��N�3I>
�,�k˩�#E�s�����lJVO����K�dɅ�ٹ�!��U���8��)��γ���%N�g�T��W]^��O^Pn���;x�ۃ^��)^�U���9�	�d�����FU�C����	V��Й���-���#�,:.Z^ՐU<c�Ը[0.#@F�X�F�2��b�v?[5F0��6ev=7���Q�G��<Ac�	�� ƲƺYE*짽�'w�n��Y�:�{� ��=>������i���x�.�=[^]N�����4��p8�֩��U(FF�o�=����T����ú�\i�x���"Q袎�w�����e̓�H綠���K�/rK�	K��@<H�#��(?���՗�x͗i����(��L��X9��cNtR~6�"p͑�LZe��۩<a������4��*��\;�*�/��`����n2�\8�ZSv��Y.����qո�۞t������O�D�d��a�rE�Øb1�_���c�#�t��ܣ�����r+G�l�p�W[B�{&�y�\�c׮֟��s,�
{���ү��m���(� �M�-�'W�K���^k$�URtv�&���Y}yga���N��F�,�Y������s	��t8��q߳��F�c��<��k���"�g��Қ�ש�_���IJ��^���w������M4l��	t���_}���6�X=l���A���J[+��v�:[7��ԓKK1vϓS�|^��m�E����U�Α��W�9fg�k<�h앥O�*��F!�u��=��De� ��W;SD�m_~��*��ϟ�
3~���C�9�����T�$di21]m�P:)S))&�<F� wZiQ����(M�!�7��f�X#՞�m[�N^�gN�,d�Њ�$�L��8�����&y���Q�l���m.��|f��ۇ[��������;����O�&��Xd|�Wŕ�|w`��C��o��ϴ|[��l?&��1�������{��^����$����,|��C��k/]��i�7L�@�&����=���a�R�-&S �W*�U�Ҧ���Gr����?C�;�D#5�-�z>$ӹ;ۈ�yQ(��v�8=fr>[*<e@�U��glLмn�㙑��5)v�͔����q���Q_K��f�Q�L��(�(@d�NE��S>�Q�x��mԸ_�M�0�L}����:[�#���O�<���h?�yg��'!���䯑�%���/a�	@��:�'�����pm�F���Z���ӆ���ߺ1���gk`��I���y�h�=��*G]�d����Mr��k����_FZ�������7{9OqPT�o�
C�4�������ЦJ5U5��{'�e*S8�j|k͔�HD5�R�r��n�K~��d��l�ePE��M���AS(?w~e��_?r
���W�ד7���� �&�ci�P��Yc�GMqOt"G��t���_����14��3�`L�����+�`S���ǈ��}���.�����{�V�W�VVu���#B32��]L��%�i��$��%8�v,sK�װ�e������	�_�4�܃>���߆�����d��#��s/+�����Y
?�{UG��C�^Y �:)��׵ǥ'&����Q��6���^����؍�����\u�󞽒~!����0�9G�"�g�d3�րN�|I:������xRt��p_UM�y8V�����H�&l>���|T3�f��j���!dd�!1٨jH�*q�sz޵��`�O����{���X�'��m�o���S��?�ק��p�*3�e�4��߿��v4�C��-ڻ�OW~�c'U����J<�^���S�րk!�.�/�@i���P@�=��%�eL6���7�7�'���J�G�j0~���ji�X��?J2yO}�튆�/����&7tZ��pWĶxͫ���?7m�"}��N%!}WZ�����.�g����m]��>ʦ�+Db�p�؝��i�n�)�]cq�J���s��6gfZn�m`�,���rE�c�ov��I�u���
�S�,�wRٚX�8	�捠��BK�^]ǂ+��6�Doё�����C���pʭ�&�HCNfd�[۸S�X<{�j~ ��?��4� �Ӭ�c�Ҋ������D6c�"�$ڎ�H=_�Z�|<��=�OOh[�>w13�ʓ z� +�?�[x�n/H����%�^
�Z"�@cZ�=��%���ǹ�s��+�i�.�ɞ����-�S��l�k.o|�=:�K	���������;�E��4n6�>o�g*�
�Fu�|K����:�S�X��:УX~��0����Yp���S$�UK�I��s	�DS8��� �d�z,vmJ���s�ۼ"�02^{pӥ��7�/6�5��<�5q4!j����(P\Њ'�˄��r�B�Ͽ� pT$�Zz|����P��v�1T�kCk y�!�%��"���E�w[Nu烠�ڬ/{�D����}���-5��N%(2jZ�N�������[��k�k�k�6q���L`A�9>w�W�ZO^�z�\��e(i�9(@
��r��S�S9�XY�}`�-��fW�<�?y��
��q�S�>z�:��ƬO�K bܫ�y��}o��e�]���[{�+�����]��}�]���!�ń̓g�Q"990����1���V��\���ڀ�DU=��%������ż*k���o��;�Ĝ˓��鴒r�?�,��	�Yw�0u�޷�^�q�Z<�^��b�_�Cs���NE��Cx���߆54]$�UtONMs7�� $���tm��<��A�Zm��h�"+J[Dn/x�w�c�6� �g���߶��R��������4�ZJ�Q\�@�3����5
W5�_���QH"
�����㧦r��uD��)2�xJP��z�!Jx�v]���Ɇ��:����F�]�iwl#�O=Ī"���~��0��[�yݼ�����9/nԇ�S���/ؙ|��+.��]��M�����V�6O�^���5OĹ����0�ۼj�����Y�x���5�9b<�o����G  ;tM=3]�E��M�Q6�Ҟ����gQҰk:����y�k��3�Ř�6��s�<k��]]�u=��p*�D�UMW��"�Ɩ�h���c�L�R^(�к�R��Oe/�B� �f�.6�����i��/y���T95��BE"�T�o���"�ڈ<!u\\���:`��O3/µ�ߑ/ģi��BMX@9�~y�`	V�f��k١���O�چx��������jsxؾ�.����;�nHmS�o�1w����Mzj��t�0��k�ՠ>(��(��l.W�ꚟ���bJ,"�oY%JXq�Ȁ�d"g`m�;��E|Re��03�t��s#V2�ՌG�jvq��(~-�.��xP�^�9f�X����c�U7�����0.!ZK����A[���ut�(?����U۹M-���K�q���������?��Y4Dк��0����w��qF��'�9��t�v]�c���-���.��1L3��g�(^�!�]b����ʠ?p�i���:�EKlSH�6'��2�sP^���/�B�I&o���	XM�I��f��O(A^-�g���w<r� �ԓ�|l�V����U-Ϛ�N���Cr��G��Y\M~�.��o�E#�H��9�F;D����J�O���Z�����>�م4�ꃁ����� /�쬤��������_D�ߍ��Q���5��#��/�d�B|�����a�F�NiR;�g�����F���8��T,KAL稠V��X�02V̇&m�6��ط@K�M�s{ܼ�q][��R�[��l��MO���Scz�I,�uX֥a3a90yVVj������ �#�Z�Wawio��'!�I����z�;.�h�f�SnK(��a�=��R�p`�;�m�0�Jڮ��3s%�e�};��Nm�Y�.�ܲo�_�o��3ę̭r����ih@���sD�+[Щ1���	ct�}�M����691�x&�#�Q�� �N6y)�S�X����,áuH��)5%F��b.���	̢q�p�%܂.��4׀b���O2�[�ٙ�?�2r1���i�5�35�SX�q������k�n^b[��x��Ӷ���)7*��f� �E�;G>V�?8V���ez�/ܝ�������o7�9rn�T����H�1��L������+��gm:$����ywme/q������]��)�E��SH���L)zk�P�n��*����E���&dD�Z�Ό󘳘<�݅s-PK'͓^�2��4�e�b��4[vT�c���7�N�A}Nt*��,�U�?"�FrjK�7�aa������Vy��,���N��%�-�9��ϓ���"/��H�I m�N���lT�s��S�_̃B7��U¯+���=��ˑd%�{8&���;��-�"	�cca�mW��.!<8T�B�Y��~%]���*��w��o���]�`�Cr�_=J:�1&����p �6���y*�oNq���NbpK���i-� dsN�\���9��1���w̍�:�c	�	^-�>�'���7TZ�2�;]��%����)�����I-!�9:��چm���k�Dv_��` �`�t\d�Cf�p(\>,*�G�qՍ�b�5�-
�}���uR�s�l����8��Fs	�n��^ٲ1։�y˛�[W`�+���'c9�v��v��]<�� U�D��zǓr�7�קn�X��
��U>�	�tּ�+���7'��H��]�$��[�xCQ�'x/S�4�W���L�M������s�s�ȋ�1�&�%���uD�����~���ݯ��i��!��� b�5���Q9v	OCV> ֢��	0���#������v�O�Bϫ[9o�i~2?}�xu��`���0�5�"�,Pǟ�ѷ`�7��kl妋k6_?>"�NI�;
>��s/ L䗑���/�Ժ_4av%k�D��N��ͱ61_��Y��� O��BrD�.�,S]b���_�o�2�KU�%�yМ��W��Jx[����k�$�����r���8cO��T��;d��4���|�U_�6ax"�ט�Rw�8$,&ܕf����'�fE�R8)Z��_�x"������2�:Ry����_%G?��%��9yE�|����Lc�拃o�3j��;W�6EbD�w�ͺ����p1v$���y���y�IB�����5��e���;dhe�Z[+-�V*R*�;��>)�?"��s���d���ƅ̶�d�ͩ4kXu��ݡ�ɜ��q�Md�3�3mĎ@\*oX5�!������r]ơ�����Kc�pj�Q2�AO�'�݀w��V�W����m�-����e���1V�Mw���8�ѥW�I;�q}�P����プh�4M�:4I��S7�V���TX���t(�>��,���*�iG?�"�6ހ����|�bz���J&HO�ŧg�����y�ՂK���f��8]���G���e��V=��*��ܯ��?�!���"e*��sqqq����ӗ��B�1��h��{9�3�2�V]�{k��� \��@1���iP����������y�j�%6ņ��1=�����Q��|y`'}�o]���=�5L�/��*��Wqa���?���C+�m��s�"8�;ݢ;��x������H���?�R��0w��vm�y4<����g����D��Ҭ�f�~����=f�x���DL�yT����;�\),R�Æ[,����ԼY�M��=,�RR��o�)��%���sk*zh9������5���q�lӆ��~fU�8�0���\��z�Ǐ1�;n�[����h��5\����ʁ{��ZZ�����U��������bcE6�\@},�.)�[�L4�	M7 ��U��UvT�����p�##~�p�����L���\0������L{�8�� �DR*]�p�z���a�I}��R�^�TG�|z�+���Y�l�S��u�*$ ��J��ŗ���0a4�~���䓬1(G�;���K���fW�Aު�3c����_��M��G5�(����8-UB�!뜉��a�F+�mx�85u��A��u��u=��O2uK+GQ(S-�4r���)�j?����E��OO��1Ϟ��p�q�Z5���b|��	�jϔ�`��,!{���z�H�/�]V-�^�KN�:�?5������=La�ͻz���d*�4�pM��|���ćA'�3��'�U�AAX��'�bŎ$�p�KK�U��5�5���e�pS���a�ƍH�L��#��IGRϏEa��""v��H�\'��2�o���?6_�$#D��1�/I��E?�~��+��}���rF�W�O?z�s�O���O�'\Ev�`b�#_�1����[R3�	��"���:Z�����f^Wq�O�ϯ�!����iC�������}�aa2���XkhTl1���1�N��y�_� \������θ��p��0Zo�a�&���1��в7�R�9U������2ߧ2b�E0V�'"8[�y$x��-A�Ͷ��99��]h�6��">LCj|-�X�����6��\&r�SBZEMD�U-]�ے�ۣ&>�g�O�3�꣓�mG��b���.��0W�ى�Oz���lM�O�I�ۦ��\������3B��I��	 ��:�ʔ�~�1�\���[��9���U_i���E
��xAG�J��+a�������.��Ѯ
�����i7;�.�����%�%%��7V���`�-�4ΆY��G�%��yX�47MsBx(�v@#�`�
[O��ڜv1��� �����Jz�+����Rce%?^׆���������Z� �"�}�������.��㶁����4vc�#����N�c!h!`�5��ky,�4��2��sБh�A�:��Z�:�M*��6ϠXn�t����pC�v=����q��pX�>�s��m���3li� D#�������s6���A�xnx���!��JjlL�j�ɏl�Ķ���(������'e|OgC�Go �_:��t��>7����kI�:oܓ������o�J����.?��;���ʾvVJ�]#�d�����!뻲L,_�Yw��eM��?"<3O��
�$��=s/^tj����Ǐ�՚Օ |���/A��?^U'�Gٲ� �^�����9�N�S����?~.��:���5i �u`��&I�� �j�$�d�~;r�f��t�z�rsY���|���+�ZA���w1^v��|��W�>�Oi�IdJ��+�(���ݖǀ��ۥ5�}V��7�cy�!scf�}O4v��Կ ��zWÔw*Bp&u�+�6�̶WK`�;)F ����ۗ�J�5�8���W��2=���E����ә�E���$/pk ������2�׻%���\��#�Gey��(�7�W��G�t��HR���>e>/,��*�?��赌N�f�N���̊W��oO���cA̸s�(��L��|�^������P,��=��e�~�	;�9>����ҝ�>ڝ(]қv���s��Y�_����5V�c_���#D7`�	oS��r�D����bC��:�B�k���ע��C����fz%�?=�6��C�W-	А�ZxD�/u���oQ�*Og�yW�Wi�ś!T����|b$1A�\�RXG�m�����[F�w����J/�w�3�́е6��/��J̀$��yA�����d w��eu�E��h�͓'6`�b�~���&�mUpv!K��~�گ����蔈v����w�e����𐜬-�7z�7�������.�Ū���NL,%*ܔlz`��>=��l��$N甼Br����0)��;w�#d�T��������z$t�N����l�]���bu{���!��Y<3�_tJO������Ӓ�����X�	[Ab���EF���-��$��4�+���
4���Dֆ�6�M�� J���Uxq�1Z��B�g�%���|��C%E�δ�&\9,`���(����|��5�;3��E+PTz� P�wD���ڌa��~�7k;�����������:�x�OL
���y��ʑK��d��'���ֿA����Ǜ�bl�Uܢ���؍��k��3��!'���c��YA.κ��+���)�ܡ���rꬶ��kކ�5saT3g��p[���s[(V:HL�[GO�l�[[��a�s��*��9��d�O�z��+%�*������hwh=��2����<i��`2���ˉ�y�DU}��"�	k� ��w�Ӓ �s9�5�s��`�`3A�IKA�v��^�s�s��˸Ul~�_ҧ�Ue|9�?�v�9C�~�^�v��b=�/�7/g�/�O�ڳo�Bea!�+�_��m��Uz�Ft6�IK�q>P��M�{����k�  i'1��-����8���C��sW:vXC�J�!�)u�C��1�z��o�\{�	�QQ��l�����?▔��U�kAX�N�5��&\�����zBaӣ�)�6uਸ਼3�S�9DU��2�Y��x���w�B���nK&�@��8)��ek9�[��R�ڭ-F[�l	hf�'��F�e��D�\/��V]�x���/hT��g�	)���dQSZx0�V�l����r���<���uzW�B�P��q]<��ք=��ҹX��k�!@��i*��6�I�Vv�W�*�Ƈ�w�8���Gޘ�}��DZ-�pQ�Ҡ�{�`��f��+��
���U�v�|ϱ�3_y-E�&��ˬ�9�z��&@�nޟG�P=MBB���R�$�-'i�#�HTV�0�ʉ?��i�;d6�Dʨ���Pl��Dyj�|�,��߇�|#2�O ��gCfPNU�T���c�T���B�"�Zf.�O�ź���r����n7�6�'y�i1w���S�#���kқ
�T��%� V�%��txn�먒upv��Y�$�G��\7���y|2�w2:����!4
3�6?g��<+��cy�ҟ,�j]������8���t�9��~6q�A9]߀	&��ϻ��S�[���|��8k�`��6�g��`L?�Y�E���"�=�����kv} %�"��K\0����?L���T-��CF~B-���91���ӈ<�pFx)n����{��ý�� 8-�~��':S�� ���z���}� !���
�Wp����O�vIm�]h<��ت<u�Ǵ7�����,�{���C��Oϥ!؆p8�{��i�٨a
�ի{<������Y'9��	��@떁�&��mW%����C	��ڻ�LA�1����Uh�ZK�����zbdd$]K W8>�����#�{�����`��,{�˶�2���N@����K�fr.�:�p�F6��'��j�l�vc�%.�a��֑�����yp��G��j�S����u6̲��Zk�B��~�6��סS-�Ǥ� ���F�� �a�����q��.���l�Լ��Ѿ���&��y%���|�����|< �YNQI4����ca����O�!�-x��CgxՄU��D�[�ʬ�"��H�ے�i�/S���	M"�����`A�|ї����#�e�6�gߔ[�����Դ���(��C��������^�'�ͤ{�t=9;��V�S�f�8+��Xn�0���F�X������.��
���j2ބf�\������F�K��k�^BY�er�9�~7�+Q)�;�4���ݩ݀(������C��G�T�����Q���d\���4I2,A/�/�1ĺ�p�U��q�';dV����Tع�7��| rg%>!f�˱/�EP�[�V�uD����=����,h|�S���)���K����y+'��@�H��G�W*uR�5�*{yƳ�k�jߌ �t���F�nC�
�݄Fi~_�����[��_�X^&����-��Zl����˥+z�B��sp�=��������d��^}�|CÝ
y�Fr;�)���f��\�`���OfF�$�ك��naa�i?i�Nȩ��>=�6���a�9�ͯ|9:qMX��݇>��o�Y��߳�4��.�5�������`�y�}�M��(D�̗����f՛E���������;��״[�ᛸ&Nx�fPᮦ��ϧ�,��zn?c���Z�
�ԾQ�x]�Xk2�;��tT+���:�
��F<��|:iе�t��6��M���������ҷl���dh���`�q����6'��a���� ��i}��+�d�O`Yn�'��"/o��[v���]P�W��LF�a�rٵ[��'�9��Jg~f�O�@^�_�������h�ƿ�+=���i88p��
ʩf,ͭ�h{'�וĳ�j�Ө���m�-��8e"��'#���}*nNJ�
�8����.����q�`L���.�,{��#�6;2C�R�o����)����	s�
z��7�e�VNj�9}�#�C��/P�|&c<F'��������b��=���d<Je|�$��Z��T�'h��X3t��?;{����O��E�����;�s�Yc\��F�(c�9�����v:�w��c(b�oR�O@���0�ppsa ��	�G����(hB
��§.�"h�Y�Ϭܨ��-�,�����z��e�/�9���Z}'�.AUU�����.���@/݅�7��|���!!�H H����4H�/s�K��a%L�A�r:�A���u��.}HF���HՀ�&�E0F�����x_��]wP��)�G�=��L7�+�l�j�v
���������|M�M�_y��Y)iA�t�y����r��_��g�x(�Ľ����]�$�����.VB��r(�X�5:�lR�����ϛ�G���Nz`���i���!�8r���aj�g�ßg�% ���F�K��	,㞿�=�U�;�gSrSW�]��
Xێe���0��N6�>h�=�Ϋ���|���X,���9�aĖ����&����?�h,>�35���@���K��gΤu�{�]j۷E�}w��s���f���zq�~tA)[�����:�TG���u�ns
������i��$��a��+6���)���H��v��ʊ)�~�l|�H2�jZ'��a(~�I�S�ĝ��n�#��¼�ŉ�e{�����y#M�L�}�f=�o������5�7J�T⬐\!a��6y�iVuhxT.��="�b杖��h��~PyB}�}��)�(|7��_���6�fn�q�$N��x���R�g��wt�%���,���Ŕ�C(i������.n���H)�wwAI��^ښu�E��.5�_���8�"g�J�tO/�J/�/�b�*���/W���W��Qq�4��ѫ�O�#W�=�Ս�����yy�3Q�t#(�rmUU�����o��B�4O���|� >���Ɩ�������2��hotRq�X��Y��J7f�U=�kچg��gh��Z��Gr����(�U����w�G$@w�oɆ�\&��2��M͸'�~����je+&��4�rF*.ة�p�A�4�Ț*-��Hw��q��}��)�S֝R�І�a�'���n,���O���!��Z�=����~b7��S�dٰ���K/F�����I/;�����\_L��e�qh����,	���f*Jʫ�����G��-Pv%���v����2�~�,X?���
 �-"9ͫ*����d�4n\�W8�x�|�2$B~�ڎ����eZ��lԃ�+�|��?Uf�*4�\�^�n��ߚg���@��+4����N���ӗ!W��GD���bn8~�o��h�H�* o�-�d0F��1QUQ&70i�Hs��{V`���� <��Ȩ�ٳ|�u6[�5���&Ϛ�M�ω��×'w7j����!w��ȴd�bb2�N)n&.�����9��m�?��G|^\&�����
����O��~)t��pZ��w�s���W+�J�$�pZS�`�^"]R�R`��T�(�咒#obo�VP#­S?d�w����"9�����c�-�)�J���6���BW ��Eԛ�w;7ޔ�/c�BML{~� [ �v*toxX�Z�U�֊ a~�~�x<z$�}�R09>"*�)nJ�T-]���^�3=�K��E)�q&�h��vAݷ)�nwڗP�iT��%q��.�D�<r�/�2Q}��P�//KÇ%	)�Y�f��`D��G9s�e�x�?��XS�%ϺÎ`�(Y�?2	�q�	���=pTgٛ_���b-E=Xi��(���fDL��8w'wI�孎�i�����v�b��O(��v_��8KV2���x����ޑ7ޜ����ZϿ�oC�kӫ���k܇;\�ؗ���6'G3��H��2vg,��~?_�X��lq���"�H6�ADd�i�s:.�P)ˍ�W�^�V����%뚿-���L�I^|H]���w�����f���	����𜢢���('�q����ݫkWN{���S�tc�~�vT`��Ō�I��[�������[Nu���B�z����4�ѝ�&��������i�&���Z����"��i���	�w�-�x�T�\��(���M'=?��d	�Mz�ܛ�v��0��c�}lگ��Z+��U�ݳ�Hċ�?���/:5�	�ݐq�Z��-������H�����3,O��T�����?PK   �cW�ADE O /   images/be117233-6f51-4efb-b1df-934e4f712848.png�USLۅ;�[p���.��A����;��:��n����28�ϻ����_Uwժ>]u_�Vu�/59TT  �� �U ����FF��dby' @����VS���Rsw��s� |s�2��4�C�N1`Q
�Qz\`J"ga�H�Q���
̥-�`V�c��c�c�	$�cA2�T�M?!�Q��B��_g���
�L?N�<nz\m�xP �Ui�+�?=J�`�'W�}�ء$��0�@6��? _��w��BG�N�7��>��bb$3�� �҂ߓ�f$������� j]8]{�dc�m��2hPh6y��RDy���!�'�E�v�D�y�ܸ�<�c�dM@�a�q�f3qq�`��a�Kb������t	���fU�;�c�u��ķR��S�7s��;�=G����T�H+��0��� �r�����K��m��� �c:�y/D������y�Е�\7�kx~�uX_A3 �o�����;j@LR�O`�'b�Ꭲ!��<ы�﫥M�2Rn�3��1=6�!m&8:\t�j�>۞R\���54a�+.��{c7�k��4�����7��7��Tf04r͘9c`�,�=-�ap#�\z���q.�)Lz��t凜k�?P��v�����aBo��1]�q����T6��iW2#�oZ��(S���|PV	�:`Z����ĩ(�39����y2�i���N^���ph0�%���M�t1b$�V�A�j�p�����L���+�ʮ����X��f�qRؑ����T?5E�&1"���S#K�I��#�E/K��k�\��������."lE�~9��'���Ą��7`L���r��p���
b�G��b";����v5��$ b"��k3�D���VS_T�D�"ӊ��l-Vk�}�K[V�e��""�M�\�<�2�M;�;��y��$���*4m�J'@'čUa�3�j��͌����`%���67j[td�&�&�f �`n��L�uTΥ��#�9�sw�i�h�non7hޔE��n}=8�1��%�AA���SC��b�"���*�*gK�Iu�+����F��LEC�*~l�O�8;��?��f�cW�:Π���Ğ� �[e��-
d��g�b ��0���1��(��E7��uH�I=W|�h��gFI�f�b�c�R�/��Ưm�¡9���#^(��S� [MH��5����p��F��֘�^���Q̸�Vnկ*`�d��W�8I�����S_KPKlK�p�����i����KCvUv�~���V��{w��?���ĤDr�[q3g�g�^����/lP,�n�H:�x>qn�w�^;~�e)=۩%��V%H��,��#�1O´o���m���vu�Q�W9I��f����$v�-��K�/b�����.��z=����s��kLA<��V(��%�^*��������^�B��zt�}�5)�@����7Nk�r"�K�Ss�OM�%k��QL+�3-����Ó�5#�	B˹V�ֽoe�{���߭�?�<Axz�-�ٿ�N�5D���b,M��+U�U+�f��F�[���#鷭S���6<7�@X�����۫�w��W�jdo��B-���-�x��nEBS���E���ڰ�������ݦ�#��iT�Z#�����:w�����5�ы��K�K�K�-�w]n��60:i�"1z3�4k�cC��j��������Ja�Ӭ��Z�T"�(�)�"x�����7/�*�{pZ���[�;�=.6!m��{ti��ks�*� ����������rj�������lQ9�r!�Hwi�hqL�	�W/vo��ͪ��?2�}���Ȑ��R��vPߚ�ꥲV���{�G�d6��(�Ǭ:�����z:����38���d������ӡձ.�g�^���tˌ~�D�BA�����N�꼟0d&��O}�m���y"N�B�Ja&E� V�oij9�/�"�9�b���"�]����ȼ�<)�51
1�p�>�[@�3��$���y����l>V��ek�5�&�yO#k��/�9�,��W7��}%����&��-����!�3�O����n�������4�jt��������NP����P��"�$��+�n�M)��\O�Cu���/�ͫ��7m���-�o���s@� u��ê��eg��Z�b_�G�ze�q�������͖��]�� c&��m�M��z�J�5疠��4�4���*�+���r��Z��.�*�*�j�+���5܆�ʑ��@o��m�עG��ɗ�:�jP�$�&�9�����˹"b��Sv��>�*Eh���Z��~�>�@���_����k��!g�eP�.(+U�b��MoO�K�°��e��f���x)�R���v��-��\]�n�=�|5� �r0X|��:�!r�!h�8�o�����E���[��-3�����Ay%��4uچ�7��,`�ܲ�ٳ��W�d�78vy����8^����,����c�¹���Fl"c�Q�Q���������}�vH��ozz{V���A��W�r�&/h���iX'�bm!���!��X?�E�L��������G�+нս����垥��y]��d�+���`���~���. �,a�@P��G+��M΂���S~��jA̵� U`+ C5�s^� ����Iu�m:�Ƕ<��QqS��� �p����ݤ3Γ�cb�p-��ܟ��|�z'>�t�)ߤ���n?���H@� �p�^��G  ��������;J�өW^��B[[�{u/��$�d<�C*���|�7&�Q��\K�_)�nܹC
���D�IG�tY���t���𫡶(�'�j�`�6����+?, ��g--�N�eO��T߿��Vp�C-+�02�Z�$�����'�O���?x�����Z���A䷗�t��U�~ᄖH_<ae�;�8�^Y���1�kW�m\�$�S������fV^I����ƺq2��xcM[�s*Ug�gN��Ԯ��~�9r�ӪL_��^���dou���Xo�u`�+�[�a��#��(��wIU�1@�Mk�e�={�,�GM�x�u�1�-��Kk�z@�������I��S��V��l�mv��*.�z�;���:m����V=r�ß��Q�V�{�q���%4�cޡk����R��i��ٵ�jM@*�驀�j���̈́Lew�f��[�6��C��b��撙40쇞r���t�Z'c�E­��Zp�ZM���Uqa��vz��_�E}/X��&�����kf�0�Y�#�
�n�+��[[�Z,��uO��i��3[�z��	�cg��#�gO���m��MfX�|#�p����u]�-�%q�P|F���*��nj���e=��I�ټ{ϼ����)2�� *c<�h�q*Q�K<j�9	wx^���#x�ZQ_�����S�v~# ~}Hq'ÅC���x\��AOAt���=te�N�>G
Q���8������؞ͪH9A)~̬��L[i��� )��[�ٱ�d]s��̈��si;�n޺�E.dz��}���?b[O��Ç�����{��B�'��sp���US�B�E�t ᠳ@�-�h�ō�w0��9Z���x��E��J��������qY�����&3g��S�Ėt�VQ%�۰k��'��V���q'ky��v�jc��C�A[
��[cs�;�Q �����i�����[P쩦���G�&��s��:oП�=�﹆yU� �7�����3EU�����<e��j�Vu�u�:0w��mT����ȱ�U@�"�9���G��k�B'!;����\���X�QI��v&7u�޽a��ݑ�k\��>�?�$�� 
�
�G��۰�7
������T"{9:E˂3��&��!/g4%o����X�}���e��>D��Ę]{#v�]��[,���z����&C)͟�d��Ǌ����8�:�(� ��X��=�z���D�4GҧG�[t�jI_{�a�n�=o,B@�Ȋ����m���OW�%�8y4=� �c�����qF��x�A%z��7F��5�>��Y�:�f�@#�K.�ؙpK�7#9r\�1R^����'c��O��Xb��8dr�|��~+�+��.�8ح�6c�:z�|,ZWs<h�/RU_��L5�n���?�􆤡��/�d��76즧/���T,^�/�a|����r�aN|&�zcg�V��W^"�,M�11�[sF{Fn|�)&WD�RN�^��<{�s���,A���5�þ>+z=L�v�کt���&j�Z�j���~�G!@�<_;3;�\���.2i{��;�)tyQ0��w8p��9��/{���k3��5�v�V\4�	�t�d	_��G'���s����`��Pϗl��)7&M�к���s���}M�)�yAa;6wY�_�hԌ��פ���QkR#�X�Z&���(N�@��W:�j�U�����MxY���j[��B����,�jZ�?�@F�+�G��ڭ�=������P�����}�9���b��rWڜQ�^��0���Mu+5	�� ��,��jb��s!W�q!O� R��щ=��u3�69W�)�6wi�������Lb�dP[ǲ�X)Kf Ȋᣠ�C�y�͏�7�)��S���qM�[�&���*���7����3�P�]�]<����;�.%�%uqQ�.�����n� ���������)��x$��C�m���!�7`�%�u��� �Xz�%�����` ��w���f��eq�vZNs!����x����Ƌ����_��M����xl˱s��l�bÔ�����y���3豷�����Y�i���X���N�5_ֱ�T���M�7��-Ѩ�Z�Y��vvy�@{]�aV'��o_����t�BB���k��t��C�GU��a� !�k�L��b-HC�}�'������tiI@�$`�Ρ�Q;�v�"��ű�Teh0Y�	�vv7��o���Q�k%���ۑ(�E�j�7ljLUn|v+�y��F�q�ޭ�rD�,7�ݩ�#���:"�~�[��L�L�8�0�T��*ڂ�XXu���_?��X��� �3�k3;�=���;��Q[<"�������ɣW3a��{҉OB
`5�ߨ9r��?�����G�wA�K6�C�2|5��u�|D(��/� �~���"oQ�m���%���yv_��KhJC��������Ъ�_�Zo��bϓ���&vU�2Z'�������������㶳��+q?���j���co�����Y���'�X� ��.V�<�Gykݗ��:�g�=%܆}������0<'�:�Q�F�j��{�����7Nڮə��B_�H����wK��bWi��:�*���'1�_a��4�J�)F�K�̂��iҢ�NbI&��ՕB�Y��k.���u�8�1XR���z.���ɤ�,�6o����P�ֱ���^�U�5{e�ݔ��U�'R����$Bd��}��%p�r�����wpn���3��^,
1tD	�)tT���Szn�''��;�'�̬�ӊ�o�pfH��݉M�D�K�3�Fug٧�f�V����O���.�����EQ��9�1y�Qq�E�����r�z�p���'�ͳ����j���+Dr����F[u!�>]�,Ɲ��*W]�]�!%�م�x�E-���Ǌ��Y"�$�~��o��^.v�6�tY�Q��"qs����o&\�E����~�m��Ϯ���/'4y����C���>�}%�ΨF;7���|��8䆷y�w���w�Ed�űF4���5��d� �2 �4��Q� ��ـ��k�4zV\[�Y�L�B�Eܠ�%��F�v�.[x	�$�C��c�O�[L�y��p���9��3_����o�����3�J�Y�����쾳iq6�v�4����\H�CM�M�Sv�D=T��Nn
��FG��%�,��3���/5f����X�!��AqW�NY":"�8��,���|��C����U�!BZ$5�L�#��2���S�G��Yy��6m���&�Wg�)��菝�
��$b���#��l���xF~{��"�f�L�[=Vl�MO�(ba�- �M@�o<ݬDM���	E����l����5���%5+�5b}�!� ��t,�&��]ә9.����U&�8q�@UT�LߌB2,/}'�;�j�K\}Fwf�&�Gf����\�x��g�ҕq7�(9eJ��y.�7+tB��X��7����6�Ƿ�]���Φ���8�8_����bO�\bI����.�La�x�'0sI^1k��W����u��;B�hd�s\�,7�Ԗ��硇 �k�.V��Q�+x�8�1�{Ĝ����$I�L�A�����m��÷�XV��U���#�|�(\�<2��6�s^f���n�ӸЇm]<,<����Ǌ���]C��B^{�1М�b��i�_y`
�}�94.qp�J��B�MN]�$������*nO<�=k��I�.��ul h��Ί��&5�5jI�b�|\ΎIdN��&��3���B+�R���IF�&(�D�q�DWEv�����T6�1kC�{r��2et�ј��V�v�"�/�����>�Y�(�u*���q�N��6Á���1�*��!;cJ�m�n �v�)�g�/����pRأaR�v�
y3� G�K�DQ�	���C�JD�����I�s<`��*k�B�{���,��L9=�.)F�\G�X��F��9}���f��{��j݇OL(��\]���Ñ���ZYM�z^�� ��I��馱�x�ѝ����]�OO��n����%�`F�E2�t������Ƭ��H�_ӑ�+ �����L���P�v�]�}�0Y'�+e�����s�y9u���6�xYx����vӒ3X!l�.v��S/O�5�4+��G�%����	�����I�\���y���7s&���|C#�j\��#<r�υ���ܗ�S[n�,�)���|~(���C�{c�O��F�I�&L\��t΋��"��<��U�yap.����5����=��`\�䤁b�XAn��5e�/�a\�0��ⱊO^�B���H�*U~���A�(x�!)m��PU�q���<�$A��iM7��D*�B�9t�����I���Jn��ư���n���/�g�+��(�_�7�D�m��	�1����^�ӛWB�<>pJ���0mHp�M�eі�KS�Sˎ�H����d 89�p�
�{����Q:�5i��
�a��}t���H�ͥ)�Jn7�/���ߏ�C�o
^N,���y+��؟�IS����;�25����h���4��ޟU,�>���k\!��J�!d�,�8�1���j}DG'O����T�����?H�k[1����E3SWt�hH���#�l�6�q�/���l�%ԾW�P�;�V�L #N/����&��|B�D,�-�r��\����	�����D��0��$G*@���N0�x>M$���Q}��mVkX�z�C�\G���4%0I�p@¸z<����� ,�����~���E��?�1�kK��;!q�y9a䆃�)�c4n��S��J{1���k:�w��E,zפP��)D7̀|/�b?�����;��{GJ�Oڿ�u�WrH�-���鸰��[>'�a���܎�i�3S#�9$H�ˆ�my� �{�n,_�!���kb=cg��=�?�D���)s'_R�}�9�dj
�\�x���k���8�)��1���1�`VV9w���ͯ�ػ7�7m�
,Ղʍ�o���X�}��!*�ނ3Q*iD3	�����E�I�@�eG���)��D�H������ �e��aD��X� dB�]�)ʗ��UY[�����7��|�%)��^��?E�xtuu��nŨ�3��DS"�E�ŉ�A��2����E$Zn�(7�7;js�xw�U��re��s����Kn38����;�k!�+ɽ�N����MLŚ׹)o!�������R�D_��#>�I"0�؞��6.��Ê<��+���^������q�?�ks�a�9�33��4~�am��q���s� ���U���E�/��?��e�ǿႭ)��)���	���c�u�������kۥ�	S�`%��n�~�RP�
���@gki��\��U:�Ra��rqW�ᾥR��@��?(=u��/(֑�|�-hZ̳�<��8ðR�N���N	��%S��4������-�#4�N�I9D�?Lh���G� ���ӈ�8���P�8�8:Gg�ݳ�y��;���r��<s�=�n�~����D!���eaq��w��R���#(���k���f���]h�[�'����~�G�~g�.�yq��ɿ&'5}�u�����o`	��������@��r���>{2T�T��Ã�ӏ�L�:���a�"uI�G�	�p�����(���L���C@�m������
�+���FlOOãwՎ�A ,�%��q�9l�$s�C���V�_[�\�m�G���Y��=<Йi�k�搀������\zya��ݼ#<��^��30�Νߞ8$�{<�@�#�W�7'a�7�~Л��[Ucߐ�u�������P�垅��Zb���e����sX��x�^74�����!�a^
5�:��N�#��P%�w����Vm�,K\oM�~�B��
n���!WZ�\�(6�^-�ZRG�&�c��}M��_2c�E�J2�A ��}��$N�j�"�h�p��y:e>|�=2��(Qы �trG{��{.�gᭈC+<�$���	W�R�M9��$��KǞ_�(�Vol)���_>�7+m|��P���%<:�y�̖e\�f�v�69���c_���`��(�6Y�~y������kב���/'�(�l��(@E�f���	Y��K�-k%��N6R��y�X��~� �"�i*��<�����,o���fr���I���������"u-a+#'��!P�sc��6d2�M��ܗ��>8���_V�����͍^�=?$u<��s�v�t�����0z2�L<�������b>��E�׀�3�i�T��̒�JلR������܅r:>G#R]�%��N��W�5���T��М�Lg�#��o��Tq���v��@k���o>���
ʸ��T_$��!�~<9�;j����F������1R���m���s��%:��mm��0����V�[�P���F��}�I��<4�#������L�|�D�=->���`�D�L��k�5�F�f{����ÉEP����,���K0n�ét��i����g�E_�ӿ�"���%�o������OQ,^8]4� ���k�z�3������5��5�����C�����ɄH�Af�oƏ��<����HV$xI%܏���M�n{����ށKR&B�A'H��bCA*H_="�+V��i�m�����k�'�b�~��9��ih���{w�=������;��e�r�O?�������sH�y^s`r�z\����5[Aj'ԏO[�?-{Cx�|�Fbk$r�&�隷@t�����L���faw4��K#���:�c�NZ��#�ҷ�����nW-�w#�o���
%�]��W������n�^7�7�7C�SζM�v�<�z��p�hEe�����Z)� ��Aŷ(T��I�݁����p��Y�ADD�_N�D`,(���06c�=�H! �	> S�Z.7?�c�0�
�|=z ��ͽs��BV�6u�%�?�#��/����u'C�0St���d���¡J��
{Dm���<��'K�!�Y���HU6����a�4#��l��Dr�]���Kl/f5_��WS��ƹ�L����x4jO=�샲ԪM�rv�9�#Qij4է~�;���u@m%�
_�My6
w��)V	oe���2��(Ae�o�M�'3Y��`~��8L�)�����D��������Ǡ���Yq�Q��
�?18�=+����� e~�CiĖ� &����?�()�-?f�L��14��p��T����������O�����(Tܪ��k��*��Z���>T�m�e5�I�ZU��g��dCs��I0T��v���ZA�#9@@�����*����7.���cS��m��_?M�[E���kC�'ek^�.�i��)]���TE�%�8����&(8|ވ���-��C��P��Z�\�F�K���7�~�]��K~�鐶Hya��ӭs,�V�rO�5�a�s���Y!�� W��Q��[y���(��ax��wTQ�|����Sd�@�����T�����U�s�L�T���VI��>�l�o?s�����R/�/��㲃f�)�|�p�^�!�	[�A���I���NZ9��;�n�N:M��0ܶJRro���^s�=�����f���@[�Sה���kж��bCT�˾���
����UT��U�&��#�>�D҄��y`�"�6��N���p��c���$�\텂�nt�./qE��_���\6sP��>oql���
LmV��9�8�$ֺ�v}7I�o������~��(՛,0a��-PY�w��L;����
��}E/���
��Y�i�LL,3�
������a����S�+��%��\��=���?w�	����`�X]䨔�f8��8r�� ����n����?4<�	������9 �"�v��u�DY���\ZG����{�MX������?��Q��g��(����	`������&:�}
�ϥķ������r�"z��r�\�����}�<i<��4_?�@3���E������;c"ɼ����"o��6pS�� �����QBuu1�D�DZ�z�Ц�*͡�~w��~w��8����$�?����SDU�4\�B��y(�0��E;�껭���<�4���j8.��[�\������]_��$7վa���ݙ�ħ�4�����4�*\����ΌC�+>�IH}�P/�z(��x����<�����z�����g^���]'�!em5�O�s?TMDz_6��]�N�L�f�����L����b���+�i�����xZ9�(�1`�o)��ș������Д�0��6�����&<'(�u)�5�\�?٘�!o�ޛ���2��}��u���؟��0Y�Ww;0�����V����`��Ȯ�:� �%mgB�E��&�(;5 ���?��߶�-�d{ $���N��z��AB����)����W�6��=��˕�l_M���	�ɼ�+ݏ�&S�\LU�"�_	}O�c3�]�j��G�*��\� ᲩW(������aDI�v���3Q#'����x�B���R�~��hi��| l�q)��3EI�;@�~Mbk(#�!�/�Y�C'\�ְ/7��ʩ�Y����W�)m��^���|��I�5����^y(C���呉S�G�h����0]�����Q{׿F6�?L�P�x����!2	��I��2���=��Lt`�w�B�EI(UT���*�=�;����N ;�).��=n&͚�>s$&�#�F	��JBB�����f��GwM������������Lsq����h���'���n}G��ts�Zge6A#?Y'cZ�c�"-רT�ew��Q��Uk��܉f�����;��#d~gb۟�M�S�e�f`��P���	fIǡV�۸X��Sj�l�����#��t�G�n��CÎ����B�;��k�����F�k�V=���g"�*�l�럄��{&�şn���Ys ow5�'t����3&3b��k�[n`�/b�B`�+̰.ѓ���T���
��PQ�bc(7�sFF֐h(e�h>r)��1����L���،�j+�_˸�?�f�0���Y��L_������rw�c)|���q��rC-	��m�!����-F�)kǌa5����q���^�͊J����=y���M�g�%�"��\�UZ|��M.�:OBU����B=wT������1��v��<�uL)��3f����{9�D�5,��A���������NJo��D�}w,���m����o|�%aN��_sf(�kˍ�w�z	j���DL�.O��XF#�v-���RH�RlD	�j�5�Di9�JϽ�֜ۨ9��Z����X�������~CX�;J�'}��;H^I���"�ye��1?���!�#�[���fgܞMĄ��:��i�d���R�t-���1���+A���1��)p�c(8�T�2�[��2�C���ܙ��:�eR{�2�X�bM��=�jň�h��?� �/�C>˱H��Uđ��}�rx(��R�*�}�I�����n���O�D�]�o?X}|�;|#�><r�X���x�f�צj���5�*�|�&?�YY��J���.��?<�4,��S��p�E�~��_���GG^"���EYh"��7�%�����+�i������`ƫ�a^�|ߞh�$E�[���������WE���̚L;R��E�#\J~z��C
K��=Lk���H�JᏴ���Lt�ӧp��z��_n����x>ǀ��?k-E���s�r���� ���'�k�%��~{i�����>�����׾�d4U	�Ҁw����¾��ETɐ<�'�������r��pH/y��^��u?G���yR�u�3${y!}���~ I-
lI'��b�}K�Rk��5����x�3�h��A�\�sg �,:�mA�0mv�N��B�қ�����K���d�2M��U�i�2X���7�4obh���|��R�W����<�x �N	�-�5D�Q��L}�X��-���|�$sr�B``��1ߍQL\?�u'O��k�w��|ނ��0�N�,TLH���X1�{ �{���!��	S��S{�r�ɉO��*1{���]��*O=NI���JS�d�`8�M�<r�&�Q�`������,]����q}�>��P��ȯB�,QQ�xX��T~�,�5$Zh��&�ׇي��=rVRD&�A�ʣ |�,��<qX���FM��o����A��T׀�[0~���O�UI��ur�@�>�X��/��4�ui����\p����xQ�zx#	�7��+c�����o��l�a��l?Y�g�)G���giC_ꃗp���\z�I):�ƥ������5w��c�����\.�@�w���Ή�C�Wj!�iW]nMU��k�)�w��+��q�����C�
�Wg4'�vG M�9�,
���76~��*�N��7�3�ИK��U̱�>��hPAj�3�繑nn��N�i������l�:/��H�%��,q��&[ ���wR����v�FS�Nh$�g�����+ihQ6?A/���� dj�]����h����o^�����K����	�0[��I߀���ǟ~o(�P�]��v�>�b���s^丏/���&Mf-��v���Y }>@�L�'>.�����v�|Τ� V㘚e|�}���:e�@%o!6J��������$�A���=V���z����-�Aj��Q��Pz��s�j�(�vi��ߋlT���$��;F�e{6�H40HP@k+����������<�$�R�%'6�S|\�D��;ؕTjxH��etD�֑�M����>�ѧ�y=�[�ЯAc����y>o��l��/!�����!7�y�Xb�Gp&�O�X��G.k��޿�L����?����v��m���ʪF"�zA�iX��#��؛���w=�a[�z�j�?T�aFa�!��O)Lǝl�9�ԷM,18��1�dvsgJ�b�EK�9�<�̨��j�-^�9ivqg�񤱮�?�N��ܰlZ�nN���C�b]g~2�1v�����Ս��?Ê�m�<�43��(�	y	�Ci�,��&Aj�=����ThW���Һ��0o*�w;��\DOi��0�{fswFD��S�8�Ӂj�"G�K/a�����ݻ�߿�$ۄE��6B�̈́珥�>6$���p��%O=a��~C.�_��N"������m��l� T��頧<tK��lt���:��_��W���UdTI�Z?Q��KfTQnx2f�X��C�5��r�\�/t�.�DM'���	 �g��rGl�թi�f�o~�_wJ���)^�W�|����w�;gɒ�ORE�*!��(��p��l=�7B	�Y2^�C('�k�mG��^��/[	�j�A6&�KR�z̬�M��l:�ΞJ���sH�gm��9�wZ.��s����A
�����>?�������������b;��.b����Ŧ���.Wǀ�&2m��T��e����?VK>�-��˯��B���"b$uXʱ�rt��d�vRQWa�q��NI^���#3�R(�^��6Z�B�����j�uO^�Kw(Ŋ	����H1鏊��\�:�+�C.�3Dͭ�����#T�_�B��S�u�i��*x���:�5�S����R��m�`���3�^�h��[m�0FA�)I��� �58�n;�{1�y�e�[����  l'�Tl����9�5 ������9C�!�����/��!W�D����r��w��ݖ8�Aߠ�y�L/%��WZ�Yl�S�R�m�%�ܦ.�٬U�+�1d"L^���	G�E�-�]�`|T�+�F[���n���}�`@�
?�1esհ聯�� ǣ�U��%�JUKN��>�@�c��HaŮ~���":�p'���ѣ����c��p�eV�h��V�˷�>�x�Pn"�vf�%`���G���ҍ��Z����5c%Qq��<�����pr���k���Z�S�V������{�}�>��r��&�Ҫ���ccя��ڀގ�Η��6E��wo�)�˗'?,FB�;�
*��\7��ۡ�����[����.�i��D��I%󾙃S�8��ަ�C�>k؈Ғ���ѰNH��Ъ�L�ɻ������v:N���=�������?-�I~DV5?ĄJE�ɒ���Q�:��F��Y�+�R!���F	�s˵;�A�N��mR�� �KtSL�Ma�]��#�$MN�*�|�c�7U�1'z�ũ]p�&eI��w0��O`�(��n��p�J$��:h�0���E��������&T�[�]��Ұ� ��|�g>��?���$�Z���̀�S���Z��dpk���X��� |�������tG��=w�[Vj=%�o��<6��)���a�`��Q$�/H��;5��l�+�@�^�XO_W_������Q���≔�g���Pe-�I�+�!cN�8��٤�����i��i����9G�S��/�gȣI�����w ��	�a~�N���XhTU�wo���V��6;9ۈ�h*�R�o���<z�=*߾I��
~�}�yt���+�)?cܑ<�^����ğ�C�4T{/��_H�<v�.$���)��b�הÄ�.��3&�h�[���6����������_�RiS�a!�U�Ҁi)O��6�tطj�9�Uxkk���SoH-��a�d:�Q�;����!)0A��4fa���h
��r��x�O���f�M�t�����S�؞HB��"9ё����-�-��B������:`�kF���D���)���W�����|Be��\���fg�Q� �딁}�	������O��2ny��o��~��c�~bD'ʗ�^����7t6y~�r�'�zA��h����FJjt����5�:�ϵW*"�o�9GqY?9F�5�)�H(���%��T�|Mb6_L�Cr�
-p0����������G�TZ��>�8f�V�����|/忂��W��hb�r}-�YU���4n����1'^Ⱦ�J�$7@�g��nX�a�@]ݝ��{��D*]�Y."gͧs�;�cPҝ���QTl�W�vYaB�w���	�\.7�˚�HZ�A9mmCo�����/�n�^�l}{�X��^}B^6���;�#y�;���.9�Ô������`��/�c��s���o�K҂o u�W�e��_
��`i�C$��� nuB�}�����gc�C=���ZmP��r�8���Y{YVCSaM�7���QX���W�57ɹm�0!��H]��4<�r��og�Y$�?=W��~`_�4^o��tu�\\^ZN��e��T�ȿ?F�9��Zi�? >@��e���ڮ��Ua
��9�1qqb�^�Y�H3}��LK��>�P��h�zJ#o�_'�le5��[{�N�J  ��"�ے���5�Ln��L.)&������W��b��ư����uN<V�s��wX�%^�o:��*9����3|��y�o�r�'��I�n}X+���;���V�h��*�%h.�@@y�g��O����=�Flw���k��B���c�6�p���m[%Q�Ac� ?��Î@WG�q3Pc��uϼ��>C��a����c.��
piLUk�4!�|� �++Ք��Y�ȹ r �%,����c��Y��y��er�C��)�ͩkgE{� O�&n*�)B*�ݻ/c �^�:���B�i�$	�M���1�����b̎����ᵗ�+��W��/��k��c�_x�U.�=�����J��G_�W��vt�3�>�­�^5/|ۼ�}x0]_>�T���*;:��?D<FA5�"C�Ԏ��ۭlw�)��*ϼ"{K��fť�V�'΂җb�X
�㑪�M�MH�>�B�£�g ��i~ed���Z}���vK�1����>^�����h��C���\, <�GB�mM�nh�jKpT��kP�Z��tR���E���YA�6[ oKt?�2~��<hmo�no��0)<K��bD+T-ʩ�@���ołm����g�f�ocV�bY��!o��<<�(.��Sл��e��)��n�+?~�d;��p7�o�C��O��3 �s�o���S w��$�$�s�C�?����1:��K �V���>O7� �=�F��V9�Ѣ�#��l[��ڒ:߾h���L%���w���h�i�T�� ����0u�e�mr�"�{�ڸր$,�����2���Dl���k��75��g7�Qq�a�I�#kcCEiڡ�.������=���&c��q����Y��Rq�=i)1S�̑�*�U(�U�%���Wq
:��փ�x��B�*U�Ҵ�1v���b���n޺֨.>��;�~�w���_u�ů������U9��
/ˏ��s�?������m�ƅ?���{�?)���avxr�ݔ'},Z�,`m�(FCwuM�I�U�v�W����nG����?.�^��qO���ã^v����H@�T+���P1kr�)��A�Ub�,����Җ�l[^�����{V�W���h�
^M2��:���x�ȩ�N�+�z����ٚ���1�����>����/ɳ�;'d���FE���ګ:���B�𒆛S��y���O&�)�d�/��Du0�a�� +�g	̤��9�jy꘱����D�y؛85: (��D'�or���p���|���|��;������?{�}�����0da�s���T�����Ã��x�O_v]'+�O���|���h' �t�t
���6�d�JC]n���3�wI�����9�8���&�o#M�~b<ߓ�"�s:���DŊ�8�U�f-񓘻?g6T'FO�x7��g<��Q�&�����*TF]��b�=ݣ	Y�7G'Ԡ�-���s!)j\݅ �LF����G9iұx�'�
���rQuN^�~y&o]F��U�twTV��,��r�i*ĭS��,{������Ѱ��o^�����{�}���O�xۄ*�xU�@诊��+�?����?�S//���y�O���o��[]��Գ�x�J5��|]�7����ζ�lka���xnWJuURۓgޤ+� u!:q*�8�x��O�C��z����.
�Y�I�QIM�Qwq�z�V/��K�^ג��¹f��C��mv�7�I?[0fQM+T�n@AL��2��{y.J�R��)j,�'4ԣ��T����֝��*o��MG莝�Y�>����׋זǱ�Z
+s\��1� v^##��_S��R|[��=�#�
������7؂`�i���e�Ɔk����M���t�Hm��I�ݮ���Ҏ?���ܡ�s7.���������j�:ϼx�}'��8��(L2'},��Sj�BA�[� �"@��:F��-l_Kw��@4�} ��cH�z��7��:i̍��~�k��M��hA���y���t6fh>6�`�Ҝ����T�˷��goR��t8T��"�#����
���U,i �p��Nz���<���*��ŭ�e�w�f"6T?e&"~�J����C�O]i�!�dGᱮ֐.����lil��O	��;ԭP��ɸw���������~�������|��U�����R ��`
|��i�C�z��Ͻp��ɲ�݋ڕo�ͶRl�zp��|�e�Gݐ4zЍHsY�;�]P���妐 9��]C��䅏?<I��n�FR���X��|�j�A��0F���&5��Žl��v�}~Ǳ6���U!�1@�̅e��D�k�@FdQ��6�APh�)�\UeeN����Q���uG���*�W��wc����"�ظ�Yx��C��7I�VZ����.���{�L��Ѽ�9�fW��|��-�{<�A�P�	��x�߽�d�XY��)���0$t�]�f`2��~�6Ã�)&0?힦q2e��1q�y��W|����~紏���6ȓ���q�;i?9 �/D�.�E��Gi���5^iNx���n{���-F��G=t}BƝK�&��ވ�3�T
��x�c�mJ%�&��䭧� ��<����
#(�& �~M������2	�	1&�n`Usݍ]ؾ>���N�8�^��;2�uv϶}�^�L��H�|�x�)�]@�X
Mѝ���F�kj4x}4wI!�#C@0��dd��6�~��Nʛ����;ˬ�U���hz��Ү,�
��*,۟͎^�lu��ᑭw~�w���x�����#P ���+�3yy�ß����{��v�~Ǫ���o��z�8��
�w�֣u�mQ0B�����	��w�F���E.�d �UP�7��(M���aU�|�0�C��$���YJ}���\	5�R�������Ӎ-��^�R?����0Ql�4��F�+�n��Pٍ����Js[:F�rZ���w��9���9�L/�#��ȹW:q�T@��Gj�i��E���Z����fxuA����y*i�2��������>�Kz�&@�gQ��m���M&⁦n茭!��טb���s��T�V����o;�g^��wc�F�xt6{�^R��3�4~�9�l�4�9Ȃ��{<ݹ�1 /���䝣�8!��A�^k�G	�:�;
Ԉ�5�E:b�8u��jn�m�l���u���<N��-�W��\�S`�x��L�e�O�sia�ѱhm�V�阸��Y�|x�l���3),&�9��BVU:F��v�����!#�g�� �M�ѽ����R�Ϲ?Tb(�|�W�(��H�(��h�8��4w� p�P��n0~��F��?�q����PGk
�GK�z[�qW��%�����H2��mK���\�<�׮�z�}�wW?��_q������Ɣ,~�70��tv�����O|�嫟~��ߚW/��Q����q������I֗��:���o�y��m����h�Y��j��G�u�3ݸa�KPs0���^W����--ʖ�.�SB�l:S�oy�rQm[�޶{y[��s��nr�K��?�R}6�pf��B"��R�j�E]W2��$���ql�H��kq�Ȍ����w,o��.WC-T�����X���'��w�9yhv�$`4f4T���	��DX���5k���P;g��/9��Vy謏�gK�����t@R��9����Cǲ<t��RzV$����oWB�2M8D����W�@=9�	@�=�������Yz��CO:�;�{��.�����-�α��8-����\eZq*q�g߂w�cN���_��pL�XӬ��Ua! ~��5��F`F?t?�s��O�4<U����dh$��`M��c��c0�,��Ps�^
"�O�Q�\y���f���c/������L����ȷ�0�ꆁ�	��C�s����Řnwh�JU�4+�C3�c�e����}|t":��U1>+�5��zC)�/و��������TU�Yh^�(�4A�jb۪n��ܖ�|�_��1�F;�J���k�g����������dミ{�R���<����3���V���=��~����/<yt����'����{���o���#Y߈֎=���`Q�y˂վ-K��ޖ<s�@�r���b���כ�s��\MW�C)h呻��'�4EW(���\�s�P�C�P[Խ���ҥsٖ��,��Ս=�qpxx�<ڱEn�R�B�
�����s益�6���Z�]�\En�0GL�C�ƈ����Uoڜ>�����9(�� ;�A;�@�u ���f��r�vۓ�r��2<a�0�X��{������q,H[�L�F�;�J/9�\}(	�0X*t�?y�9}��|#��g���̨
�@�`�q�����)��DM0�L�u�ϧ��M���� aX�]�a�6��Ǒk�\h67FU���;5��}�%<�����)c�R"[�WcO�"9�������
~�\��@��;<g�_n�B��<N�ǚ~�z�"2!�c`O�����K�6!�� t�<%��,�3�9�C�m����2vlK��~��O�k�AW�<�	��ҪXuN��b��(�9?>�8Nep���������FEl�ұ�aAJM��!�s^:s%
�`P���ծ��*�/7���K�,���*@o�k���nm5���^ױ-���{A4P���o��;z�����?�y����}��������e��S�ٓu�O�|����7�v���U}��o�+W^9Xd�Tء���Z<fZ����ugQS�[�U�eKt�n���e ��d��R>�͞��)�۵�Ue
��8s	��
n�����za/�ʥ�پb�;����y��e~Q'��Hm��2Qz�5k�P���)P�-ME�Rbr�����kF��&0�aː<wyc�Џ��LdYP�	�u P�2�TӒ�''ԦلsӉ��	�̌�y�%��4 ��|wx�vT�3�Dʚ
��-dp,
!�i�r�e�Q��>����=0$O@���~��Ơ!�p�Y�2`��>�9v���q�0ʝ� �Y�1b�8o�c�|��bJ<}�v9�k�������3g�@۶J��x�����*}y��؉y_g��{LR!p�e75��]��O�i�3 N�����]<z �,E�O�ወ)�. O���i�DĘA$F�(
�ө���ȶ��3o�b�dW�|L�L��0N�3�\��p�=�z K�"�q�hQ�i�!
�~
�!N��C�����U՞�pM����D�Ƿ2uP�ʢ�]艔49c&R��V������ZS�ZSP��	��Z4|	%<M��ʤ��௪�=��F�}:��캸��W�?89z��h�����~�O<�{gM�/����w#P ���X��[���G�}��C�����^�S�r��o���TS���Z��gr��5S�E,���2�i��+@or��g�r��B�C�i���%y���jӠ�A�1rZ����u]���(���n����g[b��<������68��b�ȫ��M�� ����:s���lW*�-4���9�4Q@����T�O�M������d��qp�D/���������})#��B㉠
q}LK���]ؤ��kq<��T~���K�09>���{Щ�n�!�R~ a��:F���UHC�u�M=�M��BJ�#��)`9��6�R�,�Q¹G�X��oz��� ל��Kq��(w�9�O�6Ia1��ٹ���u���J�3M$D�T�m������ OB/�%q8#	��@7A���Ȝ��B7b�a��9��u��ո�	�����Ǎ�<��<���.�q��\o�
�7a؅���7m~M�����lcѩn���S2@l�x �-��{�&+O��CΆ�d$G.;�a�gu��k(���eԓ�6/���=0G���ʆ���P��ɭ�+2r���������UѺ ��b��V��9/�"���(��V��ϴ t��5��
PFVF�D�+�(n*s��Ն�u��ƍ��wOg���k����w?v������) �`
���r�C�|�oL��[?w�:�e<����)+{�x��9Pr�k�[򞻺��$zk�b��n�B��`-'�[��o�Z?��|4��0�Z^�����k��D7��|-Z�����h���G.@��D��WN(GIV�������Tۺ�;�����U�J	���Vr��<)�ڔn���
\�qt|���J$���L@l� aZB�X�ɭ�A�gbu:�g���Z@g�G�ʬx��Р�����& pzԩ?C%9�9-_I�s�̨J�(
��]]����"<�?���A�<�����xc��Rj��M<Y�]���;����&u6�B��B	���S֧`4�{�'���;�Dx�8��o��t>��|'�*���襂<���Yyֈ�Gћ;�܆�"��A0�A�ԐEG�����g�M���ki|�5������P	ZހN4c����q�X�:{���,�Bjb��~j�����)��UuO ���q�d��+�b��Âcc����a�p^�ǉ�Ƨ��=HqQ�wD~�1�δ�# �~F,���&��+4��¦AɯŌ�E/�şTti,l_^�XJ����O8y�s���E`�RN�N�XO Ū�9���y1#`�`ɚ���ޑQі,�!����*�f��eЗ}��:ֶ_�m0:9>z������������?������( ��q
|��i�y��O|��;V�{��{��//wn(�������Ɠ����jl������G��;*���M�uq9�NE�߸�S�\���'ZA&����VzR�,\
ˢ���t��v�����/�e�m��c���#�&e="�AXM^<Eiv�����#�oK�R���Ŕ��BB<���'�b���1��)�J��\�R�퐨	�P�Rl�\u^��፯�MU���1P#�����
��X)T���,d��G��v�P�9���m��1�T��b����95�b�8�x]'-�hNi[���r���k�׫E��`n�!����7P�g9��R����s���[S�A���f/ �k�u�6.��	豃 S�黩�Zɳ�EvX$��P����q�T:���D-�ݹ?�O!�����m��:a��g��K�
�r/�:��H���XD�@
%�Ik���3`'WMǅW,������ƻ^�A|�m.@'��Lm��G��w��#NF���C7�?�ΖK��64ϴ�P璵1X�tm}j��O���*�La���k�w�G7��&���1e7�}N��)|68��%v��2ɡX�>X鼨/ͬ�S�W:���ڽ�� ��pݶ��dXЭ��7t�[9��4�eC!��q������{���~�ۿ�����1
�������4�������}��7�<Y}o�£��ɢ��s��걼�e5�����%��$����Ee+����Hׁ�������?��U��dRs�Qʞ��*@'�\Ly)�\�m�t���۹���*�<R�K�;>V�8��� `�`�����bPl��}Q�W�������҂U@|\7帟�ڣEdO�v�=�q1M���7M�x�ɣ�U��f1�[���1*Q���Fe;�t�x2I�5
�$Rӯ��}�� }���(���G��(p�h���G��pP��:E7�'v�L���(��ǹǮB?����,���e��'
h��`)8oK�ll���]Ă�=o,n��'�{`�g�w�����H�a� N���qm������ǎ�c����~v w*��?��k%��-o'^�m�X��1�)z��cj:*����i6B�.NDmcgV�F�v��B����ZF�Z�T}�yI,=����n�Zs���i���O�z:�8מ�P��5
�5� ������'"H3	6�"�$�ĠR���и&�3�9�A��B5Ź��z�l���eRB�Z_�
}M�t�SRv�\������_���2�t��3#z ��u�ѱ.�/!���=�)֮��Q�uuS�MS��T
��تm�S_d��쥓G���Ov*���폟���W��yZ��=�������y��>u��|��[��w�^|����{^�`��`��t(`��L�1n��5䵶uC�JݺMbfT%cQ�W�=�W�:�`�-[Y��- tq=�ݖ�����Fg{2
�^��]�|Q^�,x��DB���ү#��C?�-�nX��V�~K��EQ�b���8��	A�aW2�␋~�Ea����#-�=Q���%Ƴ�G�۵�S��~6���Ǻ�cZ	s���V�#_(�?�Ǉ2��%C�=9-�o<�~�>O׏�)�>P�Ĳ�Hj��5�&�$�����I	AX�p���bO��#e��B�X)�,v�p ����;��!6�<��άw�=��MD�׹��V�3s-̶�r�8��qj$�����m�H)]Q�6�����;�:�Ql>��y���6��}�q�����z��ʸ h��HƂ��y���OX(WL��1�W���ؼ�"��'!���ė2����ZH!��6AI����`\����Q�*V�B0�3�:⸠�U���(Dx��A�3��A� �c�c��qq{V�dC�dq�.�ν�t���w޹�2�2H�U�n�Fz)����4�!խ�h	��-�D�3��q|���b�Ã�l&�<���c$rr]�����'�h�B�NȭS�K�����w��܂y[����{��2�B!95��n��.���G׮���7ݷ����?����ox��Izǜ-����@���m>��kӭ��7|��/W��߫�h�]?��L+�Ḕ�8����)
ճ��%�&AIGÎ��ںYk,dZP��WN�)
�	u̵��b�#Un�֕8�t��`"���m�/�kg�Uk}G��Y���B�y[�)�mŮnކnږn�-Y����%M-OwuLbҴhL��J|��l���rܩ8'#Gh��������/��k��L)Ex�q��VexԱ ��C��æ�N%΍�_ �DP�ݎH	/L�杊e���W�DB�����)�7�	x����� g�%f�g  �p-p�	D2T�0/��B,��2�d�l>�Ӥ��r75<�й`,�S�<߷7�W�'6<��OGw��x$M������&.�6�P�,�@��N����8�M@�����ӌG� ,nǆH�i���`j�\�;�3���v�=�Sx?vdFD�>�6���:hSy��k�"Q�PƯ�"dtQ�|�x�"M3B)!�#��[ 	����
����-1�ME���O�1����a�$g��xp�3�C>�<����TTz�zcp��r�L4���[��:\��W�ؔuR�h-7�&��j�SF����T�-;x��uZ;0�I�����6�6�a0B0x$�+�TaN��XzG-����l���ﲮ��굞e�r;�2�P���+/�NN�^P����[{���o}�����<��=\���M��{4~�S�s�����N���m���Ǖ֣��~]@xK��N(�"`=������$[� ���T�o^Y�(m�����=A|}-p��y��)�i���d�g�����ҕ�m��L����ġb�}���9�F�Т��͹�*p]Y��ݦj�+M��AΒ>ѱ�} �얘�#�Ǣb�r��h�cC����?�'���Âͺ紧԰Ŕ��@��Xhԙb�V;;.K��(�a	�HԞ�i{f!\�i��&**�Za�"� �!��ʹ�,���8�]��<ǘr��t"L�K�ˇjΔ���0BF��X0��BO'�j��r�KU�r����t@��Sl_������o�vN����v�{�w�Y���f\��Xb�8� svu����2
p������c��G�a� � !�Hh����� -�Q36�pÑ� ���g�e�c������q"�qj˘�A)�Ɲ49b��f"43�;����c��px���(���>�kǈ�X�� 1�4]줇Θ��0�򖵾Ğ � R�D��h؃g���i�"1�pܵ Z�������t��{C��R�";^=�U$�Z��N�%x9y� ;~喣 ����<�h[w�+)ve���D�#�A����E��3��^Ge�e�P�y�)O]B�:$]Uk�`.�p�^�'�[���?P^��׿���?�u/�69�?~�#P ��z�ξ�������#׾�?k���������{^(�"~��|�P�+�9%��q�AB3�m������U����<թ�t*��HV�D9�+�f���+G �\Ȩ]�)0G�����.ݳ��ӓ|չ�y�ܸ'��N
�11;Yٖ�	b����m�뒞�-�^���c�c�f?>�dT��[tQS�X��Ky�cj���ft��Q�[�F���z| d~��T�H꾻��Іzq�����,P�w�җ�b�ZX��b���Y���t�r��� ��֨���7���5FAsG�0�����DiX��DW�G1�h��4ȱ=� ��=�8'{�I��2����p�d+9p�w�k)���s!w��Ǎǝ����MB��/�9��n��S/�Nʝ�D�5]��V{~T�܏�(b��X
��κ<�[ jx���a��?_~Ƶ��`_�J�Ʊ��1QSjfY����6��u�S��/�h�c��ŉ4.ħ��![��*�����yi���r��pS��:�! �����s7��ڀ�@�Chv��$qE�'��� :fzȗA���(�J�h����6h��ֶn���=�C��Bۧ�DON��?Q�R��R�W�PG�&�#�/Qq͋zK��׵F;��%֭>7���V:�RZ���윎e]�Dq:�Ţ��]S���Z���N���������7>q�G�o|ӓ�M���������/����������ZW�l}���'���C�\}�`��0�δh�
n/V42��mw]���ՠ���4��Z�>Q�uʁ�Wm%k{Mǂ�u�tC��{��ʕ�������0�n�8VN(]L�i��]-�aS7�%�0�W��#Cb�N�BC�,��H�k�H�N���rӆ��-�����(��9��R�j��Nպ�B	ڢ�^����-�9��N@)L�1�:f�a�"FW�N�a,(䈣��"���u���Q;_���u�U��F �NZ��J:�����a�K�Z���.p>�4��3	�Ң�E��+��LpOu�Y<-{�ᵞv�2�[�+�2�(�C�sS��ޟ��g�J���R�������#`��J���/�����\���GT��юy�D���!������P�����ؖ k�a���c�uǘ�9�=��pT5�eH�Z��4<XS�2����3>�c=D�C.�;-v�ys���'9����y輆�=*�1_"�v�"����u���U򤙑��{V�ilWz�Y�>�cp��`��[�� � �Cv�=����V�脔<00�M �S�a�Ӛ/y�<y��U᭪l��:Q��]�ОUa���'����_��D�����U�f��Pl]^�Z�{M^���J:�������k�Q�^AC�JMa�s��<���c�j�P��D�mr*�_��Ɠ�ы���w?�?��?�o��_��{�^�����E�5�p�~��Gǵ~��G����L}��?Q�>����Q�H�mO���&/Y���H݋�5S(S(�Z��-l�!�M�P�8-CY�Pɒ�M\�"��KTjᢠL�>S�J5�ty��Z�w[��}��r�%XH�m��0 �zWݕv%���[U:��	-*(ع�G2�2@0F^"Ņ��P`����"�u�x7��;Κ�wF6�D,]t%��Y-�ӂ�>�,�ޛ�����N�ф�~����sW*Eby��(��}��H�6��x�ڞ���U w� d��F��ó�� �`�"DnxK� ��|�{��`��� 9�!��E�^e,�6�5ם�_U.v8q�obx�4�Xk��Uɘ8P�#`@����ZA���uڠa�����D�.;�΃B,���P�s.Q�&��\�^i��=�7|��C`��%s|.�.�n)l@��1e�U��GC�-�'�%�`.�Ύ��r���E9oz(b�c<]�'��M�A%�����^wTT}&{�������K��a���䰇�^�����/��ՙ����,m��B=]����ԶÁ���o.�ELJ�Ɔ�{�DJ�I�=`�_��g���X�U��ȇ�''���或��&�a[�U[���9VWq�y��5��yչ��:��]R��E���[ҫ*���Hincy����'��KE�l��-A,}-�q*M��"�0eU����0br��]t�]m�ᒂ9�Z�pq��ޢ��x�����?}��;���_��E\��n��V ��h���}������O>w���W���i����F�/+O��m��.@%���i6ss�H	�(�\>GިZ%R�!@hj|%n��h�P�Y7E���\����ʉj���{먗�|Ku׵-ʮ#l�"V�O[Ȼ��9�I�S��#O�}D�S����tfC�����g� ���j�Ř�]��5��˪�  ќ&+��k�+����bw�&.+*�Qr��y�4 Qz-$4�@d����-�8�W7G(�6B�F��dE�Y�� XX���ql�X�BI�(n"@#�O�9'�,�2�<�]E��7�@G:��	.	����Z�����1  cB���B��&/��	�h<� ? o��h�����y���=���Ը7o�s�w�k�W��J���2��<O�/�Bч�㎟��[�-�i��9F���J:����ܳ1�'-aaW^[IeFS)Pd
��m�$�e�q�(���D��H,��4��㭹BW� p:�ڌ��N�H&q�9�µ�F�;:���>�T*${�W��N{����0(]�&��V�sl���L+A�x�)�<��%)��(c�̓�=�q���}L:�������;����`fS�U�5QS���u��\U�Zb
['P圻��Q��ھ�<��U��!o{�TدGY�q6�m��]�e�V�sOp��n_����WjgP�5�:�&0���'G���n�ӓ���Z-O����[,v��x:�����@�?��O���]o9�c
~#P ��1H�������O͵[�?s��[�y�j=|��D��45�R�����/�,�κiMXת�2��#�W�bF>�\��ƴ��6�	o
��K��D��l�~���u����˗����/�)�}]*�GGف�)R�o���^�MrV�/�W��U��	̛���F���2@�R�J�wB�:�L���I�09���Lm�(���EK�[�.HW#& �i����,�~.0_ȋ��fY7=ծDO��P���ƄNo�-zzE��
a*PQ�A�l�،Vɩ�s��V�9=���y��c�v]�dzL�^��<V��E��h�J/.�[:w��9t��^:#z
�,��Tŋ9��_�q����R�VJ�ʁ� J���@�)VC�Z��5Gw������1pgL�uP��i��쾤�ޒFϽu�-)G͸p.��1��R@J�w7Aa��� פr� PY�hF�9Q�q�X0&�ޏ�؆��޾��@�g�E�GN�+D�"�N���W�2p�=�;��9�Ć����w� ��12�9OF����e�0H��sz\MT2�nQ'�|�r,:+}o!y�P�'y���+~��.+c��è�O5!Ќ��s���G^�Cfފ�d����_�R�qE�?(v��~NuM�Zc�١��dXW���K��Ȯ']�M���^V��}p�Py�j�,����e<�[Jd�ZcV�xY�ZU��P�/jE�,�������%�/����J9��V�K����Ѵ|���sW��?���/��X�w�O��읟:��3���o�/����凿f�j�K
�P�z�+�.�����k��Ԃ�����B�^޺,Zʣ�Tf���&��f�ޛiћ{zs������vv���sv�><T��Z(˫���㈚H5�Rq�-yG�Ďb[]y��SeQ�+?V��'�} c☆.s-J��Ř�ܪxR�(q*�W��[�q⑯I##@�t�K��FÁhI�-0JA	o<�d���,t�7�oh��G"�X,��\�ȑղ4''e��5��+GO����% 6 ��`�UٳOܖ�����FyԠө�]���qN�BX G�u�q�Y��k 1)	����G@Q�xdxخ m%yr�%:�ў�̍���q�#�=q�ܑ��%@�:��7�q xog |:�T�Q��L�y�y�4B(l���h�`)��:�x-�����mz�.0��a��0����V:Ɣ���$��[α�d
� O���q\�z�07��6���,�;�=Q�t,H\z�#�G5�7��E�0B��j��������(/�� ��J>}���I`_BEo��S������A�8J���Ѧ���q�"���Z(c����y	Y�!��1
���]�������z���1�bU����ly��YU�9�*G�����kT���&�A6=�{��.m���_�*�����Pי|V���q#C��0@}g�����cW�*ne/:��E�M���o��{~��C�������B�;���G�ǿz����~�c����Οko]yӬ�}�XQzk���U��R4��@;�ᨄh� sr���D�ub\��u����ͣ�%6�˫]*V�8��n#��������g[��p���'j��v�j�HJ�ۈЈ�u�.^|G}ͷ�-:�ai�8ЎE�z(@���~��$������b�?l�dD�=U<�&(�8^}ԗ+Չ��\R(GEm�h�r*U��WA�+j��8\gO��m	����V�!#[O:y����\h�C�zو괈Q/:ʹ���R$�ދ�ԷZT���'���_��x:=Ȇ�]�����Y�VmwL��v
�A��Y��k���")�	?�;�9X�)rk��D���\��t:�T��P�),N!0�~mn#lL����|h�=J���ݲʂʕ���	.Vf�#
��^zek%B�����-톭&�T(D�����B�!��m�i�Rm�!0A�͸����mA��=x�(�È�X�*Sw��=\�d�qN��%��c�A��{M{�����K�+l�1[>.��=N1&.S�vv�{��z̗\KXqjY+�?!&���U�j{.���NKƢmQS�����PE�>9:k(B7�v@��H-�A��6wUHf[������+!�<��)<��j_N����h�:��*#�V�/��S�8Q�7������Q�ڮv)�5hWY4���wT�JΉ�*LÚE8�5�P�{^ڟ��l�rt���o<�]?���z���~����6y�?����eL���g?��|�l�^�w�/����x��g]k�f/�(+�[�2�B�%�A�M@����ɩ��ď��[�P梽稪�2Q��T�[YuEj�⌗%z��T��UZQ7�P��'�~ `�7R9ͦnbu�����wZ��Ts|Z��@|$�������H`��+�a�Eu�rj�
^�,�R�*�������/s�MJ������]��Őtb�QI�M�)c��yR�b����H�������J����&��G���h��F.ҏ�jL,`�7��Jqr�i&eK
5dDQҖ�;�L��Ҹ�0 x�� E>!�c�^K���c�#�|�n�q�-�f`:Ҟ��
�-���c���A=�j0	�9@񴖹A�-�U�ډ�%���(9L�qgG˒��i�o�6���|4�|�^gC�)q�Hw�P��X0?�$W�X��S����)~V@
���'3�� c`�!q*����p��9%5l|E>�)v�o�;����;E2�2P��8�F��>N����(i���dCh_c�a������Q��� 8����qJ�;pJ�>K��{M��P�<��A�P�C���]�c�D��]���h|��0K��(@U�W�%&a[���7z��7��ze���kr(t��Ӧ
[�t?J�C�9��^�����ӭ[YM�\E׾%��*��4���?ګ�xں�^�V7ǝ�JIo��P� @�:ᵥ�����&�D9?	o�j�5e���t:e�,z���/gO��W�_�����|�g�`/|����bR������������.\y��d\�v:��x��
p���mM~Y��%�YQ�FI����f#���4ͮ������AB7{&�J)]xƻJ���oe<|5�;/jR���
A�"0?Q	�C��g�r�a���M��"t�&*�����MG6(ȑ�����.�d�C\F|a����E@�K���\�?�؊�����}4<��#��T.}I?!����f���0*0��Ԗ�=C��y�z�" �%�j,&�����c�m� E=1g�J�GL�K!	�TբK�my�2Z�h��{�Y�g����Fq*�ѹ�����O/���d��4J�����@���4۲z?�!���X9N	�bZ��ō|�UY �� �aR�Z��Z��R�^�����ov�O�dI${��~�^i~m>rO۔��	y���7t�5b� �C�kf�;<��	8��� mt����r���WC���%�AJA�
�J�jS0�,��s/_s�u�J�i�a���4,��x��|&j�Sm����";�U�,�Ӹq����Oa��چ ��9[�"D�\0���O�(d�� J��xî��掁�Ϧ�,%+��!r�	� �ªm�:	3��H�m��\�W�f�pn�J�J�����qRJ������6ll��=���
�=��Q�G.c��!�jG��UQc':5�DNel�;:�W�n�b��b�9\�G�b���K��`��
#�%��z�po��H?��!|Q6��uu�ڻ�h��'?}�������?���O�����( ����y��C?�/�����������Od~R��E�P����^���
kO��[���ZZ���ҟ�nhKy�P�뺼Ϫb�Z4ʔ;uW1���[��s�vvE]Ѷ��z%V��
@�R=��4:�g�P������) !��f�F�(>E�;SF������$�3Nt�q�CUѓ�[�K�J����JT�T��J��$�L�®�p�J�xGTڮ,��@V=�:��(>�ѮS����΅jy=y�tf���2T씜���R�xY@�P<{���;��� ��G�ԢOl�p�"%+ⲡh�P�U"wIj��F��z�Ҳ����<��6^8޴����	*� v}@���1��8�8Nt�G�V��UC);6���q���b�Ht��|�΂��z8�Q� L̟�H oz����CD�mo����� \�Ĺ�1��x�*��M;�ӈ�n:�|b��uBS�\j�D0��a/�����1R�t�xP�3O����Y0( �y��@����L�C�����H�R��PfE~,��%�P ����x�)���.�J�`Z��©�(m�M�$�%�5�-�C�O�sr�C12��� �!�W��Eyd�䭒ǎX�5&NiUp�U��7b��;���62T�G�T�I.eùr2���_Դ��i@O��&Z�y]�e��I3�}�����:ڇJǪ��hy��jm��u={��2�9S�G�vVQJ��1Y�{�J7[�ԓ��kԔ��1~��?Z�N��{f����<����������x���]��9������>�����?)��O�����h^+�Q��9���������y�𚨤�� x��yܨW�}LO�����b٪ͺ���HE����|����Ю�B1�JZd��QNK`"�J�x�Y[�7�8�V���^#��50��bg႒���B��EhA���d.AG���D	On�"Z��x¢>���{����n�T�N=���^��EO�-�dt���ȵ?Q-�	��(M0t�"�S{U�eQ�kN�ҵ�Bw��>騋ɺI^�U�x�� FR��1�C ����d?�vY�"oxIj�����g�v�3��:]'�D�� ���\�C���Ԝmj8����ןqv�-��ѯ;r��`5�0ۃ���X�~�{^O�F �TS�)��?=&�;��w�&��%�6�<a4�U� �H��5��|q9�m�J��=x�����Ϟ�>�{ y�l��߮���� ���/P�������s�C��
1J�/b4{��}�C'��'��^�.j|0����t?� ���*c���T��j���2�� �X�:���s �A��=���{���тJ>ν�Q�9�|�1!T�<�
�d�ׄ�%��4%�[�����`�Y�Ǽ�{�Cގ������w&:�:sź �&�L�^������m�X	�m������v��*�Q�f�uOv��Kى�Òsjk�d��[!�:9dϵ	���p�Z�$ֵqKf�>ߔV%�\6�rFJW������yu��C������ǻ?�#�>�ܗ��w���	���~��П|���x�-���pR�N�����P���*�8����\���/��@j)��7��<JIZ��H�0�F48�VMw�W����Rv��Kjx �YB�#�_����#�E�suO��,�����rR[�)��VUc�쫔����܌�� ߴ(:5�|o�P�,�2T��M�RfvK
T݌Jc�kJ��T*KM�&Rej������;ⶉ��iJ+���Ӊ���=z�k{C<sms����keF�C=,�ŋL�rԷ���^�Y�"�yϵ�@XDd�1��b��HA��`���0��ҧ,�[IЧ� B�H�c!dߔ�t��a=&����!m� q=��n�$d�e�䶣�y��P/C)�M?@-j���/B�;��*�$v2��3��-��׸	C����1��i������̰b/���	�,���@>���sH'AB1؟���a��o���?Tv��b21(�����M��w�Y�JEi�j�[VC^�"_Jp���#4�� ��� � St?��٠��Aϛ��d��9�8B��c���?�a��;�C��
�lR<�#a'�+/C�c�C��ئ*�Q*5k�F�S�\��?햛��m�$",U�����BN/�"����1d4X
�1��Z����]0*4ohw\�]�u�7Ů��lO���D�5�v�G}t��VbkZ'��I���a��E��ʘ?1�T�[֤z�{ˇ�Z�,���ˍ�l�X���IY{�_�.�������?��?����G��1��?5��1>tsx����o|���?���_��ReW�&�����+x梯g�����V^krۏT~�c��9Ԯ�� s %Ҽ�B4�E	K�f
]������+��n�d����e8P�q��p<'y�Th��ݖU��d��&c�4K@�fupբǝ���M��͈���<����Cߕ��c���/FuU�j�}dC��Ze�m�8��$�ے�M�V����lW� 펾/fM��J�=V:�X�ߥ��;��M��.9��q�P����cA���^W���q�`X�T�Z���q����P6w�JVUB �U��a!rs�t��V�����H�@Z�=�J��{c�Z�;V^�g���%.A�E�a�SNx@[���L>r�S��)����Y���w��d$��t��A#������r
�D���+�č-9����3���;�N��>�>ձ�\��x�Ό�;W�YjD��x�� dz�Z�р�`�cġ���5#�L?�@Js#���a��:�\�@.�PŇ��{�*clM�<t~.�
�����.۪�GA��G�����h�t��F��j��Q�v'��� �\ν֩�zq����T������T�9�7�")<0!Ä���ꛎ%�p�Y�&㺊���:��vd)w�Վ!����6"V��Y(Ĳ�;3�nך3U*.��`��-��������.�EA3{�e��;��J�S��FO]�T�C�V}���]��B�ײ�n��/ձ�A4~a�v�Z�T͎1h�j*[Gb��qUi���pTj�����.��;?�S�;�(��q���1 ��>����������?}���O�9a:Xz2M\��4)�cOP�J�1���%K𢡒��%��/�����.�kvJ��[*�-���b�R�+����yEEjԐE1xb���MM��n�'��fF�B,�x�������]��ݩ(�cu��n �% �-jI��E��^�l, W�vT�������m�{l��:w����ؑF�U�G�w�m�f=����T�z�ե�
���x`_�YDP{,�,vx��Qڕ%��ٷ���|Wz�䳱���"x����yD�L-~���	������x(�e�h@<�.A_�u�'H?���l�����k�e���1 �\�:�,�S��*͑2��<�2��9@��o��A<$P#&jGP�Eγ����'���H3N,��C�n�b���D��7�`hxpQ��2���mx�� ln��:er�?����*�v�������P���bx�Ѹ�X�I_g^���J>S�N�E�tO`S�"W�S��T���-��ֺP�4Uɤ�Gq_�F�%�*wb�|^�����z�y�������5�wj�UZ��ՠ�F&뀇+�"�)23ON��ha˕Èa��;ݳ���Mj8��:^�J�N��Z�R���;!��&���<w�7F�	�����nЉ�YAŸ	}�Iw������)֨&o���i��8E��t-�wԳA�ѱ�u�����\%��e��ݕj���ZV8��&��P�#�-�{x�0��`���ؘo�^��DI�cJcs�O[�Y������/��{?9�o����o~���}�i}W�\ z������=?���}��~�?��ǟ�۹ҡ3��D7ω(�#)�Qd�܌�˓sk��4n ���C�K�|�<5��稛Q�K֔hlg��]����1����� ���{bTqn8��P�4��V���x��k�n&=�1��!���4-�\$���HYOh`nj�L^4���6�'�V�7��M��֮ThbGip;Jk�V��vG�E味8S��'�a��XO5��2Fz��W�����Ρ���G
�����a`�iJek��%p���E��5pKU��yϱ]<�H?�X�ےR�c����Z�U)�	=���bf���Q�"S@?+��֢�&�*�p�~�t�bq��xK�佥T0ǚu�T�����%��^z�щ'��r�����-�x��  �5����X�;U����n���{i���?0���xé���e��9�ʹ7>�� =� 1%�	�b��h'0���̛��Tԇs$SĞZ��1o�b�0�rօ���* 3Y���Buo��2�r)A'ڈ��`�¨�T ��O�R�ܒ`��&$B�!�����ې�a��R1�eP���v&�_@R b\�f���f#���f�ї�T=�yS[��Кc�L��H�B�d6�[�x���u�L2�a(��k쵊�s�d���Q�� �q�W���*�VӼd=���a�A]�E�8�玧>�y�b�W'���.O��Е��fH�5�uA:��
NQ9�+���ײ$ģʥ�U�c���Zܓ2��:�� ��������o<S���}���?t_���. ]��9��_��3?�g~��_�x��+�b�M�����f"�۾Z,�)p�͚d���YP�����\�]>�^Xښ���V�FM�o*�=���� U�P�xC) ����FIU6��w�<O��9�.|���,��N�KV�y���G�p�����T�8 ��mf��7��\7����Z!.�̥E�u��M��:���-�h��ɤ)�o]ԣ=1ReH/K��bo4� �,*��z�Y��8�8��_��k�I��!�.�R�r�{��+կ�s�S٫���Ty
/�jW��b:W���X�������Yx�T��[�Nw2��x��L��ܣ��Y�ˏ�s�E���+���Q� fA7R2M�>�?/��a�g0�����q��xZ�X|.<�X��8C��;ѽ�ۛ?�h.��w�����J������i0PP�PE�s�Y������R�C&,����p�V�a� $Il�GV��E_������6�̞��Yyz��R� i*�>�A�J��&W�wU7�.t�`�S�bU��VC���&�=��m�6X\zOZ_q����wj+���R5>ƴ���:<D����b�ߧ ��!L�3�:@�Ǔ�i�2����(=+�Z-L���1d��8y-L�Hwe;bF�=����*�
�T��7�n��9�$�qh�����Q���Y�P㚌Q�%����
�1��RF����h����ز�r�r'(��SP�h��
�e��Z����<_���ozzx����߸��W�����o�����ܾ�^�����3��Ļ>���ҟۻ��7oo_��N���J���G��C
��e�Ŋx���5��T=�X|��㵠�� I���`E��;���w�{￐���E[�C��z��R?bʱ�I��6��X�X��S�}�����M�|i-h�^��޸�(�@J��,��8��h�>^���o�K����T��m[;�l�\E�m��9���A� ;�g�~E��T�f�F4�ΏDi��@͜F�j?���m����i1�f���b`�$����"���ô8��}#6���J��Z-W�����KtR�6jP�E;.+���<gh>s�pB���8� ��1�}='��雎Q���o��2�s�讽pZ8l����\�$TFkL����*�/wbؙ��Z��T*v c�+zw�G z��i��gx����Q� �� ]�'Kݽ�0�*O��_Lǜoo��0�38X!	��<�Ѭ���8`k��F�g.�"��4I�Y:��K�xԨ?�kl&ǽB�='c�k�;��М�� W�C������,}ᔰ��G���j׆�;�j@~M�����)�!!K���Y�bq's��B����O�F�BhC���|yC��H�-d�O��̀H+u(H!#�˺?��֘c�;z���Z����_'�b&#]�H]�xp>.
\�'��8,���~��΀�űj3�0�vU_b���W��ui��U;o�G�^6��r��-�~͕=@o�jb��H�IMk�ۿJ��x��T1.ur[�����<�׳�R'��[Ҫ6~���_��O�����O�o���g�6 ��|�j@���}��w�����_\�Y��v���h[�*?(|�ذ�4n��>�'����%�i>���l�C�+"�V��v�'�3�B��ݒ�잫�����WYֲ&��|��(;�罐w�$������eC訵N�(h�>Y0��A���m��}��8���ݘ�T?]�C��b!��Q/��%�l+�(����*Jm� dH�JS�:���@���B�IM���d�PL�� ��`��P���	0�s�(�9��ߴ <@Z㣟���x�!�Nc!*q"�sJ5)�6NP�U��]�����>"FJLU��0����[,x����qa������.]T�������'ד� �:��VA%��2��S t� ڢ��M��Kt}��|���j�9������S�YF��`��Ӡ�Y����uy����{A����{ =�w���t;	 ����HS�a$$�X�9���2b��?�9���0d�����G)]��Y�"iF� f&7|�4<�d(��ڊTH�c�,c C3Dv�,Ε� RMt�X��!Ŕ x@��Xl�����᭓7���D�I�98�;qw��$s��5�[���Ϗ�M��I�/1f65�3�"�Q`e��tH'BUeԱ��<gϚ8��f���٧�J2PIEW��q�C�PT��._^5�T���u���>��T�~���e�,$��
�k�*�,�{m���u<�!_JK# �BML��\�Q�N�}g�c�S[K�x�eZ��*U�u�k��_��z����������/��w�+w-���w��/~�s߳������~D��FC��NE뉒�)��//�HMP��vH{�^qm�����M�5���m! Jd�3�y�@ojb��7���)�]q��R<<i_��"&�".Ķ�0Ƅt�p 5:N�c��&�X�7 ���t.�v
��e0��G��m�uC*.
�ѐ��Ҍ�������uT�L,2b�u3ͲWnQ6V���NK�=�c�p�0n}}��[Ʋ$�.g�ױ��	�"��1M��b��7>R	]4Н�<��.��n�Ei��ZxD���c*���x$Z I-̂b�0s(j�텲TA�B�:��E��?���TYP0ވ+�Y>�6Yd�� �fb�I��6��`�6v�n�zH�����~\l;���pos7�9���қ�iU��A)}i3�>Bؓ/������* C3��3@�*M�;6�0�=��C�q�\��װ+xݬ��pB4���<f��>i����4�Y
Ox��h��@Qa�mwݐH���d[���������A�Mz �<ᛅM"����̈,����6� �)�h���O�1�y��R=-��V%�,�j���@S!61M���:�c�������Z���s�%^�3U���/e�̡���^�d+N='�@���U��;��%>*���5 �g0�Q?u��D���ʗZ?�/�/RK�����pO���Ȥ
GM:SZ��˵���j��.�1�^��A�՘�MJ�M���)m��c���5@���VWaB݇�j3U�v��l�J��*��?��xv����~�����ڔ����W�����[�.�����&-���w{ɭT�#r�E%��N%s��cq ,�h%��}��~Z��^�ቨ��b�5m��g]Y���h��S�Xy�}��G�b
���I �f��BH��j��3êff!�M,ܱbB��ius9�\BY�zr��/��l{JC��V�7)V�T���"E�X�:�(F�NlǊk_?T~�n̡U�f��7%�œ����m��K��6�(r#��B_eפ.!�,�gz�4:�17-���d=#_����K��!��j��*lc�]�V�3/�ip�W�B�g�N��6��m�P�>�j,�Ɣc� ���LI`���p]BaO�V�F����N�f.�7�;<^���@1��m@� o � I{�K([�����U�6��|��+l�x	(�Hn:0�n/*����F��;��k�s�����!���o�"1�gl��0.Ό�9b�;>]���я��jo�U�bx�08uz{j���h���s`�9)d�D*$���Xa���%�R�Ɍ-�mS�R~r����)D��N^2)j�{���$]a���c��\x�@��Cm>�4G<I=a��N�Hqo`�p�ݓ�S+�*�X,��x��$0D�n#��`��E���z0:���f�r+]�6��~���]DF�<��l�!b����q-)��:׵1T�*z�7D�/��������(tD�w�>M�_j~+d��BL\���T�pWZ:�-�b���@�}�j5v��m=��~�#O����#?���ݷ��R�����]���/?s�g��߶�>�W�s���WT��%�y�r�S� j�:m�3'�	�4e*]q3yI9�������˒~�ѹlGJ�m	y.]�R��"�3Wt;V��։�碲g��jC�r��M������q�U�9�-ë��mZE��- _��Ӆ���?�����_�+���9y�۲z��ߒ�&�W�q-V��o���	M ��6Q	[mJn/ކT���z<kmms!��d��Y�O�p S��L�e�fu�����#3���ʸD���~�7q�,V
K�s����X2�XԔg\�BF�wY�u�<h�|��ks��������u�����6��+j���J�m�]L�*u����� ��1Ϩ���3#x����;9hm�;�Gd ��7��]��H�1lo�5E�Yɛ/���^g_;p�2t����qlN�JF��'�>Ɠ �#����!�!��6���6������'O= -��ǵ>��3���#>}f|�~;̐�̂�v7�r&�s���T)�C��&l����x��(j}� ��
Q��
�A�w(�2W�):��Fk<���Ы�/���.��Æ͢f~I`�����iE���0����c����`�5�pUE�l���RPI����R�,CI�o�K޺�t�.�2�_�=��Ns���2�95�)K�jv�k�n��С��
�ϵ>.�wň���۪�TC)l�$��r�2�u"� ��oQrVF<�w�xb�5W���X�V��������M19=M��B|/��]z���V���ܯ}j��������_�z�$w������ν�?�-������r�&���]Rq��⵵N��Vt )�i8U��pi���#X�"n
�M�9iį�p@�H�x*��k�w������G���;uy�S]�;���X�]V�H��
��X=Jo�E�(�@�{��ˋ6X�9"Q�c�X�x�Z�(`f5t�\Tk��=	W����W�|x�+҂F�[��=��wC���iK��/��3^��e�T4�@�VS�E�"����E('�\Y+���AsҵmpT�����iq!妪��Aڜ�:'
�P.R�e#�ȷD��hha�)�J����56�L�B��j�NO`�>ٌ����P����?t,c��v��ŵ&���_,��]���;B%^`�����虖�`�~��M J1�n�qp�H�4j8W&�k�3 ߏ�,ܶ���I�G8 �)N��iƄ'c��f��|��a��E8Q�>;��g��,ǚ �k�ӼlY��(n�5���_�J�dM?;�a&WD#l�Ö����U�?�$ci̓�H�sC�f�:@���@UT^�C�)M=�>���.�&H�G- �:	�r����%4Q!vh�[շ"y��5�p0N��{&�~<S�K'�%癪MƬ�{eY��=	HP�]�5��6����P��܏���h=0P���	�=�ǰ�����G�b�u������Yq>�{��}�\u�-]�0l�*uB�JX�t�6�m.e��[i�3����Oţ&
��>�i���� k

x��Fi��
��Τ�(ն�^+K��:���C����/~����G?�������}�:�����̍��c�����?��^x[�hq�ݒgH?z�ۙ�J1�'��*Y+�b��i���^��`���4�r$v��!<���������v'��{#y�ڟk~���MI')բ4�[? �p�bA���w4��  �T��W��PLƪT��Z�$Tvd`\:�����%�ءn򱀜T6ګ�{�؆Sԯ$��腐	��sq�Y;�:gr��a`� �(≋C��-�
XCU�v��;>��9��
�u��*�h��+/0o� ���ja����{!�OXS��ьF�f�1~���cIOit|  lb]#����kW���t�b�� u�M=p�MyB�&ϕ�Ǻ�q5�|��0f�L�:�D_T�N,�\̘o�=6�����J�/ L��1�?�z��������o�5.fۅ8a���G�(�s0�=�|� ��3SSZ�>�j:?��9>�1�/z~1ߓ�b�^����}�����u}��B�YD���HƑ��Ġ�`�<�򬙿�FN�����'�iI̹^wT�����N.^Ĵ�w���Q2������D'u���
�z[�Z �ߡ鹑VZ*�-74�1(�-cEu�3�d\�����WE�����x7mѹC��(EѤ���7�'':��$2���k�A/@�ɼ2��Nǥ���6
����(+/�(,H�6;�	tJ���8D�X����"t!��e�;�P��cE 5p:N7��B4��>P���R���$?��0{0�Z�
+�T�z$F���Jh�tձU]�\]E��/?<,��]x��x������a%��������ڏ�܇���>����~m��|2�h�9M�,�S,/떼f��SMـ�d^��	l��Â�v������J����R�j�z��{%8S�L�F��)s�jj=�:�o6A����j�^D��Y�����+Z��^�� 1��2P�lP���Ka��r�;2.Z*SR]���w(
�'Z��|�cU£�K�ҵĽY�
�]���n.��J@#��1�x ��MN'ަ�9���\S�� �(�;m����a��, /ݱ(3K�9np��&>���qDU
�:�.��@���W���JX24V��a�����j��ӡ?�����5-n@
�ahH������Z�wW2���^�-=�+�`�Ƕ�t��c��� �ee�dR��� !��.:d�4b��}WcA>�sz�y�餒'�ȹ�7��x}aX�L8�e�{ �Y�;��3��8���tSɀ���Tt� �$���������������QO�\����q'V��/La�h�yb�R�5�y'��E���u	���f���Ųi��pe��t������F�Z�����&+�*�s=�D�[җ��Q?W����f���-"_c��Cz�E��r��26s�|x��12HO�v�"�}k��X>�e����2q��W�z�s��x5����7�v�<��	��^���b��aq"JYG�sW�[OdT�5FC�!B�����P:�X, u�:ךn����<��:���F���>�Rt\4�©Pd4�(�J����b�Ts�4�v���s�͇��_��w~����w���.�6o����w���{?���q�O]y�M�"�����K�g��x��V\�`%���F"�&�]�K�6��)�7Z�J��Qݮ*&�����\ifTD��I�SL�*�DI
�O�
Q<T���� .-�^ȍ��H�J�������YQ�6H�F�>֒���%ћ�sbT�M7ծ%D����]�S��X�
��%AuCqrA���RI�n,�n:.QƱ ���Ep�Z���)K:_�C���6פ��X[�y]ű���B6�J�;=�5t7Eס��Q�F�E^�<%=�x�j�k1\w��J�6+��#|%ڝ:�	�4F��z��_�7i O��-4�9�O���jf|��1W09����X\�&x�A�ڇ�8�����&���6�I�s�������7]t2=����1�~Iq������\1{Cз�U���L�-~a�fl`<$�x?�����tc�dl�9�y=s�ey��1�2��g�k�;��!c�j �nm��V�=�	M%�A��^z'��S�:ؖ�As���@j!����o��� ��e{������A��e[0Mt*4�鮰Ǩ�'H>�42��U�XU�����m�X����},GW�C��7�{��bM�s$��)S�L��my�[�[�(F�}�(8P幻V�(z؅5�bؐ��0-�A��\՜ ��w��踯)�,�Qۆ���5��;�����7�vt�ٱ�>G�����l�
wd�hю]���RG�_���6�j�Ӓ�O�(�!ۯS��yBg7M�(�p�u>�s�*��o�+���;n�g?�����̤�xݡ�9��=��?�3����ɿW�r���Ԫ��T(�:XH�ֶw�FӐ���	+��x����8��U�ċ�`t��bp���lu�<�rV	3�ɻ��J�U���؍e$�Ta"P�NӍ�7=U�/S������t<���X��38(AY�dt�����:����vs����Psa"�v2i���HT�]�*'IE+/��Pq֪�bl-����I�NeTRՆvS�չ<p���S5�p]k	��X�Z$��U򩼐��6TQ�ƶ�;6E����h!jʢ���������iluO(>#���];������:�!-�N�
����\���������8�qԢ涡���m�B?�M{^��FP����^�M� �0	�r+�use�����c�T �va�)~zӚ��q��q�h��F�/�]����)����I^h|�IQ~֩U_����@;vC!"أH8_��8�����̏����;�醚�2d/0hi��y���10��构��M�� ������  ���k.C�^���<�A��1���cvŵBl�"~M?�K����s1 "�3a�� T�%Z��M)�CL��z�P��r�K�bJ�WiʓV<�t��t�,�֫+��*��D �GN�����2VnGkG��H`�k�U���*C	\��2�x!:�+�6���级��V�`P�ǲgѰZ8�Ĝ���{�"��)Å>6su��ˠ�+��I 突�/�vTyf��׹���>�R��)>�{A� El�8+]�����	��n���~Kiq�2`~��C]�Ŏ��L8��=P�m���N���ݣ{ok��nL��?<z���o��?�ʏ�M�:{�u��엮�����߿�-o�t�	�bcg6�j$  !}g�V�y�c�ǒu�K8@��cqk/(�Pܘ,��*y�NUB�v�������{��K�T�L5�{����1 �ᒐ�T~x���_�<rVG�X�ְ{}�!���[w��Z֖�ڕ���+�T�ʞNH�#���I?T�-/V�N-���A�wC�:�r�]]�^i'3��4c�kqa�����hl�}�����V��
] ��\���~b��N;�|��M�aР��b7����~"��P��\�]�:MU��Wޫ,����" V��z���Y�F|GM JU���8��3�`��֣�7�<^���fc������oP�'��1�OA��eJ=��&"G�$�4���A����$qbN?�X_4E<���x�0o{�>r�<����m(�s�68�b��LҦ�=�V������g��=:�ft��ma(�w�[����#:�����8��m�i��H��\��g|-�kʑ
X����V��q�
bU@���}3�/b�!P�@>���G:f�I�6�Q�h%}A��
�t<�g@g�_�<�!���X�-*�)U�������2�g_�v�TiR�;���o}rJ�����Ø��u��ӄJy�g;Ґ���ّ v'k��;<r�����u]+�>0�� ~o*^c1%̅G�}T���Ao�~k���=.v����\Eu`9 |�
�s1Ym[�CL�+IP	�b�C:#��VK���}�[�xsԼhPGC�FK@n��mk|1�'j5�XK�ت7�������w����7������u���-���/<�����������I���Z������n\�Jjb�L�H����"�b-��9����bA��K7����h�#y��[���ե¼��N���ۺy�O>�5Lu5)3%π"�N6Q[V8��;�)�^�!�jLZ�cV_�Rt��`w�i�t�:2���]5S�J�^UH���1>����'b����(j��fuFU)/th�_�Uk�06�ֹ��6��@x�y��RWӖigxKP������E�T5:
����By	M�q��:�E��T�??g:?���]@B,����M�������P����s���l C��-hl����G��](r7��S�00D{�͞��o�e�̖���@�/�zh�\�o��O��f�|
�9���6���\E����Fat�/��I�O���H�nP�m���0�Q�D��㻮���i�9�7�m*��0aX���w\0{�.�Jt(Ug7��s6�Q_3��	��a�ڀ�5�o4�'��)�(�����@�]��'5#�����&F���z9�8p�)�)�bpLu�	4	Pݍ6̼7���ʎ���=\�o��-9��.���(TUlW]��Dt�5��o8�h�3���m���{�iu���z�.J��vt��k�:<<��U�M�H��.���06�"�ڟ���>8V�R�@T/h�^����?��4F� ���x�`B���i@u˲�+�	5�0P���''�l[��T�^�:���Y��O�Ɣ0#�1�9�!�~�t������HLZǽ��v�����'^�����������;>�쯳_^�������7������ް�(]�+��K�4y:Y���pP����K�;ei�:�)�_�#�����0��A�K������)֧XՖ!*���}ŭ�Ҵ/0��ߗb\�� ��`y�cd,�,��@���k����ajIGE��J�G��
��n���;�j5U����5�\X�#�����	��kcZB�9���Y7%*�m^Q�
�{G��&/O��NG�� ^j� @��wB�C5�E��T\�-گ�����rṋ�,���t�X�CY�#��#��ݩ
k[�4W�cJ3(b��)�X�b��,\�3�!f��
c�֚�8zC�5��Q'��{��׿3�1�@2���U$f�WK ��q����+T�9um����a���}��>0�6 @J l�,�_�#?�\E�3��}��3���@l?:���R��Bx��Ɯ�4�T1s��O��Qk�ǱmƋ��}��w�ޤx� X��� [ �=�y��ܦ�cEs���!�w?��f��r�����F�:Y���a �iu�;<�He��:G���Rh?`��FV��+(�hTb�����|h���Z(#e&`轒�"6�����wM�<ŧd8��!c}�қ��е�1g��t`\P���U�T��)����UvY}%ڲ|ic|��}�?��^��*\�=�V�3���mA/`��14��C�T[��8TC�E����X���~Z'eң�J)}U5eq��Z����굱���Wc1���g=s�Z�mC㼐gޒQԖ��1F��q��ŜR(��N$F�A�:�ã�����>���/�����E�������w����í?]��}�\��Cb�ɑ�����}QM��:�HYO&֭&ш�p��:p�`�Ǝ
b*,���Q�#�B�=��je�@���ؗ._u���Ԝ��C���vS���J}��XȈyEM�?`��eW���V�.��5���!�CwdqS���ɏ��	�G�&��D�*�:։�B�HiZ�j�!�|�*��-�au �����wM1��ޮ<m6��˱����+��ڲ*Z2�:��;��1!��*�G%�!��Ƨ�����!�1#�ݔ��EkfP��$����a8,`J;����ТqSC��#(DN��C{�ڟ�%@z ԣ�w^�d ���m�����P�N>���9{�����1zv��X�w� �p,�l< ����s2}._����q��Y��V�;o��8^�i�3c#g&rP���g���?H��8��0ۑ	���*��wE�#YY:O�. ��E.��܈��1�����3� l�'Fw-²�t�EȘ�j/����'��ۂ�g^�F#s	!����W#%�c"�������������pq�	q�k�P�����Q����PV��RŬ֢�1j���h�-�6�V���hI�#`w�_�� :�t���^O s�	�R�c��bJ0>貨�"a6	e�տ����F/[�:��)q�h���	i�^0�	#�A�z Ce��sMAcI����c��Rh���s���F9��@��fu��\,��_�9��
�Ͻ.Fb�p�P��H�S׽F��	�[A�:@��P�Q��PY#e���t�";8Yl�凖��=������W�U��k��������O�ҳߵw垯W(�7�@��1�.�*����vM5��N�`��~�g�3�R]�͔(S�5 �G[�,�x Z���5�PJCV�J�ڭ�����c��� �D))C�R��Yϱ�)P��e��	w!Xʔg0E� �B%�5t9��.9�mQX�n9�jj(���ʏX q2�!�E6U�
O��?)nk�xM³�
@���қ,&��i�6�����x���4��@������wK�KS�cba���^�u��_c�}2���1���9���͂��E�Xx�x`ľa\jR��� X�)B�z�0VX�*�Ff̸u>(α�5���f����M��kI��*��9.��Y�7^��ӹ�����4<}�g�m��ŉ�gl�.7X���>��a�T<'_t�E��v�����]��4(f�S�\ $����7͛�6� ~x�>��`���GI�Vq`n�nt\{���8���'�Z^��m���������ðr������c�(F���ڐ� o�����}�A�t����6�U�a2wC�0�q ��t
#ǽ�e�Ѡ�`���E(���3?���` �0�`*�����Vre:�=�ԑZ��j�Ԭ2G8��i�C���VMT�Y<��'9
.a�#]�'L)�c1o��^W?�� �}��+7u��5qcK -���F��a��֔C��6����Sn�͐��6�5u�?l!Ef:2�[b(kR�;�|����4�l�x�%�uoA�GC3�Q���A�ZI�=�1��o�DohS��NB����vw�A�����k��F�ݿ�����/�?�����{������O?r����پT�ͺ�=Q΃	��{��Ӆ6&^�Ģ	
�F�q�_{Ld��I���ϙ����%Hq�NޖW~�}���s��W��&�D4�>攸X���º���)��W\	��c��.��ȑ;Ȥ�L��W@e���D�k�'�9F@Fl��N�[ ꦧ�[ ��[�ӓ� ���VܠB�6q��$ț]ѩ��ΔkԢ��;��9��[R���dѴH����H;�8����� P"��vϿ��@��x��M��C�s#'����	bԊ�ƽ��|#�9�n��m��<�P�� ƑUDUxs,�Zi�=���,,�fx]�����,޲X*���T,ǀ�c�t�>��ǘ 8����@\~6"�`m�ax#�
4��6O�hF�/��I����\�Ƿs���ל&��r43�%o�u�e���.�c��g�TZ����ʌ�5_��M��D�è0oCx��\��@��*n"�d��1�
���ǵ��I��:�<�L�G'2.y���s�Ni	�=VIXG��`"\��6�006���d9�C���Q�����P{�)M��r�G��\�'o+�}QsZ<�>�;�pǇ���4�{=���c$FF�С��m���Eۮe/�8Pm
���l��iƁs�Z^�H�w�ǔ���]��-9OQ8�P�I1���p��Q�yA-z�<�)�s���?'#H�6RSGJ!�ɛ���RN�$�T�;׶Y�hzU�:[A���0U�L�ikQ��"(k}ڒ����IiQi��+W���×����S������{����%��O�� ���3��]�}ｗ�W��u�	C�����!y���YPnhIV.V�o}�>����BlwJ��^�����qc�w����֬��˴K��Dj���'�A���\MO��&�<�	�W���R��)_�5֦͂�	�&v���	�~%��4D%5-���P�o�NG(���I7m�N���zY>@�+ݴ5-TM�|�჊�6��R���F(�1o!7�n�-�D;������	�Q��e����B�I�7�:�s���HV��Ea,7��O�fwk�yp��1Q�B����5��yX�J�%e� N��Tp�^��+Oэd5y�u-i��u����	���ᭆ@�-YM��E��hX��}�N��DXX��hTt�>K,�6(���cνx������M���L���&8�'������� &ئ� ��LPz�d�m�=�1��N�3q��.9m�^J��i�߅j�i᧩r�m����hj=�A�@U��Jg~���c�y�D�f� ,�lN�b�є��|&���*v'����Ωs ����:�~�3Xyq���}J5��;<ς9��֮�� ���ÙRb�Pm�1�`d�Fx!R9r�1/�v�2�����b�ݖ42y���PO�ky�5�k�:t{�Rȉ&�0�Cf�@V��S�SN�kB�f�:.��b<_{������z��cs&��Ɓ�Ż[�^�Ds#��g.@'-Xc�f�uڲ	s'��Xt;�D�,F5�1Se����P^����js���Qx�F9�YI���i���O�:,KI��K��>3�>��m�:�],�Y��P ]=�����ϽW��/�^���� ���{���S���U%��3-��Dj4�~��e��F��m��Np��B�E�H�c�*Z�
^�������TTZ� Fu_ŏ�%�R�yY�J
4,с&mO7�@�7��Z��*��Y�Y9�
%��$y�^�X���Q���8.Fs-��kBk�ۊ�"C������G	%�AɚV�fT��
�j��D��d�,5
��.�Jj�a��R�*`um�6�Kz^�`�\��t4�Ȣȴ��rHz*R���cx_����nJ)?�!h�((��A��X�R\��o�p�k�p��t�K;J�O��$V�����I�9��q���@-�,-&T�Kc�v������:�H_d]q��M� �QET؁�����ΩE��3�Z�v���܈K`lf �@t{}fw"~k8�<�V����o:W�H����c5��߶:}��c�� *��G���02`q��j��0���mX�Ax{�F�Q�1R��mF^�FF��=@��=�J �A 2�x3b�\�0�l�k׽@�uI�b�nO /O��5��
<�3���R+���0�3F���,�c���}�k@�"�����KB���@�&���Sa�$Q�'�]`��vK>���v�(���[;z��x��]��&�"�\��>����ù�:�`
�
����5hK
����6�Ͼ�Jv��Wq��ơ)1�﷤m��O&�&(���z�:L_��]�#aLDx-��C(vsy����3�@���UI��6��+�f�����z&�c����qƑ�g�&�>[�Ց�4К� �+&Qep{rX�떖�������O����7_�W����_7��_�����O��c�b�^!�9�.eI���Xܛ�ń<P�5{a,(i�aى���`3�3��Op��)c��n�jx��'��tw���"�BEu��P��ޮw�{Ci�����*f~z��#�F`
�-�֦�锆,����+�.Nt3Bi��hI�!C�NI�~��b;/_?Yt����d��!&�c��Rq��T���uŤJ�E5Mߑ���P�����މ�*�q�1�Ay�V��}#~��¦�+�$�11VV�G�ےw��B���V�����N�lDT��Y�,0��W\�}���A���х��(h]?��=hE�y���h,PE}xr��|�gx��s��~7��v%/����9�	l^^)XP�ۋ�۞a��@?o�bA��"~�5�P#��ל���7@�K>�}&'ߦ�L�g�I�
��9;Ǫ5G69;B��&8y3��Mh�� `���T�CtZ��]�3�8E����D�[Rbւ�7ȧ�0���V���63���cq�=t�'�v��nQ��6Lov�CRE�]���z���(
�;�����9r,x��t�Ð��2�a�ub=��"�t}I�dr�Ѩ�5��
����\tc���˜�d�K���,���T�#t +�4{�#6/�Qh*^���6�ʲ��k;j�jnW/K����MeɬT���TXe>��d���H�6�7�q)����|�+�{:�i��� (K����_�T��_V�)�rݍ�j_u��XY�(J.�ѭT����κ~�l63������F�i�1��{�ªf�z�5Z4��{?��~��ɻ��Qy{�������/�������ν�,�򑉃�%��+�@G��pg��ߝ+l��h��D ���XRC`b
:ǎ
���rRP�d]�_�MY*sS�,�� �oM�S�5H��rpg�<u�³��,6ku�ܠ5��s���C��)�΂�3Ֆ���-����� ��o+u)�tU�c[�+7��I��g��Y��*s��V]���*\#AaK42E ����,�ד(oXVIYe��F�gX�N/�<�ݐ��@g xp��e��ֱ�)O�BM���0��k��� �**BQ�PR볊+ր�3Hk"f�g������M�Z�a�S�<G0�T��%$����?��`� �9Å�rM�}䨇1O���d�!�����p
`va��%��e�Ĝ�O<.N"�n�I��m0�s|���V��x8! ��if6^��(�A���8f����������ηf�4�̉��I���w��Oƚx�EgP�Cc�o�MŨ�����:�F!��c���w�ěǋ^�f��)����Y*F��ɩj[���ɋwʡ���b`,8N@���p���y����7��3�?n�0���� �Q�_mq<�L�u��j��
w�1[8�@���!j��{�0����<tG),.���$�J�v��T��p��[Z����Jϟ~^�3�J�����,�>�}��(g;j�ޑB}"p�(�	m���Qn��\u�l��.e��
)rk¤2Ȩ���d�����?<���C�[�B&ڈt� b��Vjm0��4fb+�;��Mjoxit����F��̗�5^Co�. �����ǣ�sq��}ʩV(,���5br��c!��;�$b���x7n��6��5/^�".�b��E��d���B�L����,Ҵ��s	uj��CiE��meV�0*��� ����	4{ͩ9xk���\��������X⩝"ݎ�cɕ��j/ט�(�E������*�c}�X��4��P��+���NU�xS�������ͭ8�X�߉�M�
�Hϡ��n�B8�Y�#���eV�l�Sw��	:5�m� ����b�UhSY庐fC��2���ɫ�x�I�PB̦ҳ��]u��Y��,��5�q�;5-�J|#���,�JhF�Řk��)�@2@���?�����`v�F� ��*�3�2��:m?����9��f�6������8���*0$�ہ37]�!��A�a����)y*���y��+x��� �Q�6�m�`�*=�������	�y/y���oTd�P'X" �۹ګOߩ�B0Tl;�kL�D�%�:C�;��A�]��X\�5'e��ب?9��X�6}�|#��*"�c��	�.�C�A8 �!]��q���t��;��H�����jj|�%�����J��Jʉ�
�v��u��D��iuQ��f@��u��Cy�m�c�q8C��0d8#b�kic��}W��8�g�9;��R�<wE���\{�~a�N�I�*�L�i�g.Z���CL�R�v=�\���v� ��B�#C@�o���x��/��>f�?F���?�,)a�{�91�/��oQ�Oe�OԄ
�䢲u�pQ�#�������{��/���׼@�5�?����~�����z��[$���6W�0(�	qn/LL*�s�ֈ��i*���[P� �,{(6��&��{�qױ��B�*�[\�ȣ#���rC����k� �=B�g�Zܰ��n��R��7�������r�ɱ�6�"��2��5������/�W@6
u���M�
��� *��H7�D��� �Eq�x#E7HA���Zd�Je9��˻*Vc0gE�&W�r@�WU�;�=�9M^(�2���1Je#-N���B�ց����;4��!�	+�]��yZ�ʔ����@��B�-���f��)T�����+�ӵ��Sw<�AQ[�Υ��` ����Ƞ�#�ko� vQk�ך���l�4���1�c+�<n��ɖt��� f��Ε�ӻ��\g���'���_p9_�a!��#W�� ���4*,``�?��q:���@0��%@C(72�Ab��l 
|���9�) o6���q���@�f�)�lx�� �1��%����!�k��Y(���CǷ�2�朋�X<�]$�Z�K�C�����j�P�����A��/�N������E�֔}��@�Fxb�<��\K�T�ݧ�]�a�Чv9k ��!�V�u��Bd�� ����Pb׎z%(�^8R� �������cH�.�S�{�6�vtt�<��_�ϼp�j��2.����6�5�fTڢd3E��26��	��斘�z҉��\u��6EtT�GD!r��V�y�pT��x�4o���{5�G�ˎ�yu�/!�u�k<t���Y[�HbB�eQWի�����^�y�Ǿ���x�5����>:X5�����=��QF���Mf +*��͋��jB��TC���*yi֨�@��V�����_�rk�13ő��!�,�|;;-�TK� ��j���j���#��l�Γ��8݊E��;)��r�`	!�+^ȵ��D6\l�&QH�qs�:Mf�36Vv҄H#�/31��9+*08�³�Գ{un�ꗾ�%y娺�����GzK@~�*N=���LǍK}|������H�Ha�r���hd�ܤ:.���o(�8�T�Bej�,a2 3�.�d�TG��� ܪ^T�,����#M�b��ό�Z��X��F�X3ji��  �nWzc�ii�`2�|</\'^sݗ$|�S\.Ӧ��Q,3s��H�ϸ��@~�~Z�8��x0� &���D�o�E�����;�� $�,X{]k�,�c�[�Y�ؓ�?y�q_Ȉ�q�&�(��B��W�tn��ѝ��m?Y�#>�Jc�q��(s���<�w�����P�Ľ=��颛�#ע���8T]ܜ��0	G��G�ߺ�I�䓧h
?1#�x\4Bt�2�4Ǩ��aC�u&l#����0��8�:[�eO�V� �>�����5͋��u�r�[�&A�X�~�H=ܕ+�U�b�{RA5Ga�|Ji���GKM���^��������5a_Y/��w���37��QW��G�o���A����D��P���КS�t)h�:�_N�I��s��BNkY+f����\aΝ0������!��X^Ӿ`��u�d/����4�u���e�tG�ʛ?�����?y�s/��ox��o{#���|M����/����]��M�vs�� ��L�ΩԖs��0�1���pɸ����F^�:��,-Bx�^�ţ��U�ގ��E�CQQLL�\�EC�G��$q�z�I�CD���+b�Ha�C���I��'p�s�܀4�`q㶢4$V�i��S4�|���oTMN���=1^���������ϸ��v_�=�Ⱓ:��)�JG����'�Uv�&3�*g;�G.�_,jr�z�4	鴰7���Q:�@*�!i2��u<���,Pį$��s��ǢC�|tC#�UΆ�	�7�[��Du8���,���^]�1.\�)�w-���b8��Q3(G+ȝ��k��;.�&m͵��\�>��.΀���l5D]i_?���=� �O��^J��#cB&��c����G���� !�00BA�IW߹�P�d�a�<��b������%>@���l����x7���u%N��T�m�t��j@蹦���EW�L��K�}�+�NS���d���x�̉tL�szB�?Vv;*�>�HE�'�gb��7�󎿓1�����tk'�Iv7v�x�'�ce��
����f�X�[#��ڄқ�?�㣒!D��4�S��qI�0H����SM�{��AᾺ�kr�*o�pƋ{�7Wf�V �A��.F��BM�z��iO���XU]�>ۊkw4ϫ�ܛ�_9�7���k?��
:�!��͛ԏaJ�*J�y�����n¢y ?�����bͬ@ކ��O��i�L]Ǳ);h���=Z����<){f^� i�K�&^C�HԖ�+�}�l�ҹ������>�@�s�������}�b}�[v�v.�Q��ޢpJ-z%�S����dj�@�����`����'"�+4�0F*��ނ�i��m5L`��[ة	�PGnP����;s\�Ŏ�6�7f�W/ܱX�	bB�8r�bĻ�@���^3k����P#nN��n��,]�O�!5i��㚲`8�-���YQ��+���^���ϡ���6mv�,ڬ�8ωJ�SNV�Kλc�,Z:VE`�D��D�wt\Q܂Rx�-�S��(ơ6�zj̼��r��;�����S�4ht�-%-� '�8�C�W���4�Фm#"c�e�#�J7�Ǚp�Ey�y.����r� :?-�y��H�������<Z{���:��>|s���iX'����1��67~�?�;�= :X�ܩ�kvɳ'���6P� ��<LYo>�9ش�����f�u�*h{��l`ƹs=�	�s�7dC}څ
�6Q���w(�k�
�W?�� �c9����*�8�R�а9�ƖcJ��Ĳ�"���rN91u�;zpo�BgQ��>�_[MDh�bFIa��jX`�r��cOۨY�"(V��J��(���םM"����Z�`�HoD�EȊ�X
0wLݦ�Cvkݻ��
ב��	�J�Cg2�g��U�I��dU�C�����[��T6V�ac�Jz�"��J���坏h��I0�����\@v�;��J�.ջ����8T�]�=�C��})ʅ��������ֺ�.鋞G��G>�	���=
-�=�W8d�5j;�in�i�Zl�i������!�Ih#��5�6���cAE��rgX�z�o}������O��o�z������k�C���\��}�*���uZ�q��Z���Q�gSZ}��[�m��&TĹ()i���3�L��Lf�aZ�|�(n��=O�$�"��F�a����Ơ���������nH�050�(G#4s1����b���b���e䴡� ����`�$��u�Y�c���rY�Z��S��7;ݐ '"�]�l��=�|%n�ՊG5Tէ��"�y�̎Ԋ�'ʻ��jص���'�:���-�����,P���I!	R��X���^(x�L�$
��F/�s�k�H��)��PD�����1֢8E��bm�����z!������@3+�U��ӹI;gƐ�ⶫ��y?��'��8_O{���ӢbʝKg�0��cI]�K �El8�)������S�߹��O>/��X��W;�L��ӕ'W�{Yc%*7��&���8�πi$\�(���=�Ca,���Etw[՝�wV�s�B򲞌a�.���GCcAm����|x����b�{��mBl���AT��;�0煈�O`�)���
�W�ar���x;����d��^��2̗�+0Eu��מ���c��nkJ\�yhR�����=[�f���������LWt�$A D(8�b�I�ѿ��(����L(x!b�1"!�á�	�0�h���.��������ogf5A�䈬�D��әy�6�~��]�Y�zV��84ӈ��7��k�m�Od�3JN��;��p\@�ɞ�qh���7�%VQ��մA2����ɢ�u.խ��~��\%RgR���8��(�pV����4�AP2�D7e��^%�y�"S?ʍ����b�:������m{�C��`m�O��ti�24'-|fxOU�p�UG$Gߺ�/�AcI�E��XT#2a}��2;
�6q�,e�X��p�)ϟh3��;�Q�/~�k�o|�|~��U���׏�Co8���_��g�0�oԏ�ԬU��ɜխ"R�H�?��B� ����q�a��W��;�5���#���'�}�!�i6� ��h���0��`�7�t�]�^��ϔ^�W0Q�}��G6�5b��T�Ä�'#X��9rm5`t�����=�붥�1N��"1u>���SZN�t�A��`N��ڙZ��2�~�p�B\".�@�St�ClB%:�� �i�5��O�<Fڇ��*��0�E5�	�U\�Ӡ�(����g��S�@������ ��L�_:�q�-q�b��}����`ۄ�7�׉	r�Q�Z����"e�)�H�d\�ګ�'j�>�,�o	X����&��_�j%��:i���R;WZ3����(p�,yZ�!/��3/���x�=DPb�%�;�9K+�ܚ���R��K�4�
�P�Ƭ�$��:2i3�T����&�m�@,������쁕�s�mp�R�|� �]���$���lZm����b0��H�T)M�Lp)�RP�|��#�����IF�z-0~��#,d�.[�W�u���y'=��M��,ΐ��<�_�s81!!hP"U[����Ùg��@Z�X�����y�F���At\4R����l�?z��U�ͫ2˹�$$\,;��pxC��3��ldOv�tu��^����:���P0�Ym=��x�*s֤�]��b�5�3ƙ�y����������	�5%+���P�����^��x��Bƿ�4z쳵�}gӒ�r���s����6�l_��[��_�`�]�~ww>����t�N����ɯn��j�FC8�M"kBHw$�VF����Y<�����
���o���z�JƵ}�)r��Nf��g�g��#�!����^��� �0�A��9�����d؂h��z�&Pn�@Rf�=�f����h�5�@�YR��F��L �6}�{Hod�2�6��i��(����\?$:�p@#�6
0D�E�>kX�����i80�q�@������9�/�o�^��7�2��PTq\bD�:�$�:��2�}�����\w	/8S���;89f��^b:"�_�T�P��v���u�	>��)2�]��1p?�`�(�����Je�%gL(jeuJBf��u/������$G��lC�d�@OĮ�~J�!9���>ʌ[��EV�|�������{�'�k^WlG���OL*k����{��tׯ�瞱�2솷�3�T>H{��t��$�d'2��)}�e���$��v�y�S�+Zck��y̺��=�<dYS�?2z�;�"�����f��m��z�����ȸ5�	�"J�	��U	8����yA򖪅<>�2M�M�H��ᾐo=��F����*�ljZ$�<���Μ��I,�q����V�8Ҧ��a�,-rmuj��Pt+���$ (���Aټ�K������A��/ʺV�|
�؞kiј��]��C�qL��s�	6jf_�s�;;� 1"��7��3���v�d��5��]"�췘;7�[ڏ�~��g$�$���d�6�J�A
�H�=�޷� <����W�(�N(R#�bB�Yo�������'����Wx����������}��NZ���A�P2�}��xk]�`�k`wP[�8@�A�O��@��
��&j/�Gx�u�L�Ke����vO�l������no�O����u�aM���6���6K��Վ�t|���#���FF�]cT���+٤*�񙄷�9�O�M��}D�g��a��P{��b:$8�"uf�U��Uz��Q����z[N�h����5Y=��]�ִ�3�X+*����B�{0Du+I�6eLZ�5��5���ByI�W�	[��E�k�p�bS��k!d^�u��Tʴ�'h­�ޅ�El?H2⪄y�Z�s�@��Mh�3�o�Э\ 3���f�'J@LL��wP��Q=�r�	ل�s:9��;V3�܇��Å,2�WڴñN�,��A��~������|)�Ē
ZC*����.����B�W�����;���?c�*5��*��K�v]�8��gA��L�ʟ	��֌{�7�1�p��h 1p���s��@�̂5�p95Q�1X�?�H�C��+$�E����\�k�D�}��c���Ƹ������A(G���E �;z���E�"`/$d���LbG��l�c'l���ğ!�s �e���1SuƐ��>��3�ęJ�j�ht�����q��	��l�(��c�\��8�4�Lhh�A K��J��n!����a'�ꝛ�����	��r7��U�T�#,���,i�ֹ}�%A��O�*�Hn�H��ع�,��>K�R��]�(Ŀ�S�
�����?Y�o��L��� 1q�m��gY��(���������{s����s���?:_?r�W�[w��_������Meu�3�}=@�/��r���b�v��*DY90,y��z��hpH0p�ĳ�����Ԝx�赆�O�"�w�	���}�)���O2������y2��(A%����Y��f��x���ߊ�YYm��E�mW�"��� �C�敬��~x�G>��d@[Z�c`�����lD�ڃh��J�*ӈ��n_�������㽭=���� ���u4�����Z�uH�g�@���t�%ѩ%`��E���'DT#3r���x�-s�_\2n�υ�"�J�=�m�"�k�:�2����24�
�%�쵄My����L'��T�	��mβ��Y_O�������@�w�ޖ\��	Q�����1a��D��Yf��B��zf˅��!����w���RTE{�ܠ�V���d��ᓺ��+�����Xa�?s��'�\��������-[��>p�N�Ȉ�4����.@"C����E�<�ԉ7��K΢�8�IRG��:��:&EF�N��NlfyVC�G8���>.PL��u��&:�,XI����Q�IA�B����Rx�d�io%�}�7+�|G����
;b ���ѱ!n�H���$yz��V�V;K`<>�����8�2�>E����ν���>����l2�b4�|Bpmi�{v`���x�e-5�g�؜&~�6�:�w�Vc8�+wn�����r="!ٜ/�:��%�d�[�޺��5Q)�w�G��4�<~�����_?˙�ؤ=�k���M�|���G���hk}_����@[�乔��ys�ǣ���o��{�П1#�^�����/�}���_�+Չ�����\�Q恈�µ�L�W�t��N[�?��6I2Hћ��JOb$����;.v�N�4������6��_;��z�3�]�F�2�zd�n�tm��k�"Ⱦ�548��:&����m��Ĵ1�olH�z|Z�{=U��c[���]�w�]���2ׇ��h@�/ɴ�\X��_
W�����w����к�q	XL�j�6k����%�(�v>Pe�fL�Ù���q��Y3j	H,�#7q�Fށ3#J ��� �a1Iw�!%�ѐc���0���X�A2�9�Y�1FYZ{��0%su,{	���dJII�NԂ�-��dl���X.����#:�QV��������	g5ޝl�W�?�7>���~H�cbj'����Sksk�v�n8�G �N~��詗���p�h$d��3�M�O�8�3�*�%&~����Q3f���H����ɗ�6�_�:�N��9QM�@��z�-S���I0ŷ�w�6�������Ғ\�p�q�R��=��Ĵ4��<�f����"k[3���mj����=b�qg�{�ߵ����=ét��lî�U��2�<��>Ğ%Сĭ% &�^J�R�^1�A'��<�G�ǱOK���|M�uQ�6�v�2g�2��(��킥��(����	�_���U�Y�wְZk�:�����Z̢��%�����������۪HҶ�]���Ͻx�Z��p�;M�^L	Pf�ء�&*A��/%T*V�����_w���&K��6f68݁'_)�I`k�8<g�O����3��0���
q�E-�=�u�V���i�/����~��{���>�|���B�co|���#��?��o^��jݼCFp�;���0��%M����͍��	?x�B��;�2'�ș���#�%j���.,Xd��N�e*e
_���`��0�nF�8�-fAC\{����!n���HO��/�T����#�T�+�jx��ng*;�@uԊ�x���o�ԭl�/���%�=���ٟ��M������ɦ�uN�
��BNщV�u���F&��g~�8a��(lm��͉��?�e���;@�mK�M�{��K9ʈ�Ӥ��p!7o��!ץ`̈́���343D��d2��k�����Ԉ�K��3rƶe���ƺ 5n!`G1���5�ue�y ��%��\���i��T��a�l۬7�N6<OF,��������X�~�4�a�qM2�{��3e�B�Q�ͶH@�2[��e�O	qϲ�E��z�f�~��'ה9�88*|��S+�F�t�R �� m��E�n�2� @�`����%MSX��xOe?˔�\4	��j6(GW5�&e	��oیu���S��$����]/���8	�!!6��
��L�]Bn8#إ��g���B;O�Z��B�?�$�ID�����f�/o�$G��d�ԥ��l���h�+sC����1t�TAׂ�f�em�w�}g9���?�)�V%Q͂�эj�:�/]8o�A�L]; 1 P?�ȍ�`� 7�J��q涜����Mv�S�ԑ�E7|Oj��À����3_VV1:��[�sE��s�NóuX#c}d{0X�Y�#�����Ax�l�ƆK{<�(�?ǽ�E5�rԸq��T�#{�.��W���v�\yW�����l��{4��'�����^�G��Gʡ�}u��wO~��jІ��&�Ƙy�e8���pc�&G-�L��47�S�ؤ�Y�f�-� @���K�:�f�!��P����h�A�8dQ��-8x8���¦�1�,���0ӗҊ�%�mGЏ���1��͐'�Hш!�61��(2%�}#����qp�J���9��t-�1a�����X�1l���Y��q�:gh��G>Js �ɹ�aPud\Py�u��o�{��5��&���t�Qh��"�c>1���}��:��5#��Q�H�{�u�(��L}���ێ���~�X�6����B���44u ��CX��k�lL�p&ЦL���)���O�dH��+.���cv��>|Ydvp�k�q���R��sC��9^+��g�	W��za�*� /�T�J+�K���D�t�˷�!��Q
>���uڡ6���'����Dg,���y��}��-�o���I`��5)&h��3�$�Ǹ���	��������%�"���d�-铠"��GY��q�DX��T���Ȑ���Ǥ��=J�S�q!`��z"&"b���<w2��ަ�WL��<;-�[5\�����qpq2�:�m� �c�>h���;*���#/�>9�$k�[�"�I��5��:jf�t�p�$@�v͙��+Z�l>��+&2:����̹~��O�_#�uƟ�����D8� wv��=:9��톹��*�5����NX�������=t)6��8/���Rν���#��C��Q�rmylsS弮���Cb�s3c���$v�[��%Zz)��di��9��;G��t'\J�>����)�}j�-�2��0�??�����i@��~g"�`�8���8H��������\��b���t��?���K�<����Z~D�~d�`���?����{|9�Lq�uP��U*Թy>��P	�.��v��w�-Ό��mĸ�(�􄌣F�� fp��_�-Ѝg�Z'd[K$��͉��wu����F�7�_[��@��g�{C����_l3V�x�dh����@둙�Q8򵒏�4R@�Q r.�Y�р��hQ������ƹ���O[kg��K��l����4T���f<aA��F(��P�,:�ֶ22��D(��Ϛ���x�Ѐ�)w(\�`k��^ߡ.S.d�A9�A����iʺ̲�3�^Y�:�j��Wȗr�̄�U-Aϑ�:�H���k�<�ᨯ]�`�>>k�H{)p����V��eԮW8��X�Sԡëe�� ���Yw�"fQ�9��4^!�X�f()8I���� t��$���8lk�l~W���Cg�g����V������g�o�kF�h������ɻR�.�����(���Ő��D>̔���>�f�/淋��u����x��)"�'_������(�ˀ�a��+�bƫS��obw|���m�4������\�ث8Z��`�Bi0��֫}��p�ZfwEG�糌��{���*jU�Y�t~H⧁�BK��)�\$1�3P�n�t��X��:Q0ě(O��\+�? r���jTTH�t.�d��\i5��ym�B����>�V���.B(���sb   IDATr�(�-?/ŘU���'D�u� ���Qm������G��Т����e�>"(1@����R��:Z���L5R�$So�gT[�K؏[ӏ�xԔ�M�X2�nXJ���3���އ�#���]���Q�]T^R�B,�̋�j��w�9���?u㛼�̼����p��eU��D���	���2eK��G�T@=1���t���
�$�a�[õ;��-Y,I�|z@%��b�.s��|V�4ř�Ibt�P�zf�佣�%LYf!ݐ�ٲ�xVCNif�\O�w�h���I�����M�K�I/ͺ.��Q������|Y�!pb�ILCHPg�}d]�dU>��a԰��
N��c����6Q�cQ� &3�a-����G�Howp����q��^G9�͐�=AxC���<X��TWT���}�fTJ��mC>�ٻ�.�z��t�d�fd�/{�����>D��\�$����F�1�C�zd�N=u�	l	�=�'��i$�El��3n��d>xr��7��v���4 �l�v��:�kr�a��yw�$�;�����y�:��g�镧�x���}�<�ҮHߵ=+v�cӧ'��C߯'��x�N2?��}�@vYr��� �Ś%�V��'08?r��'� �#�h+rb���%[ mvfV�lb�O���I?k#S��^�)��:D'�y�li���(4����ܕg��X�ݵz������3dn)�J�s���gK����� ��<f�9e(���K�&�D�G�kem������홱�iK�X�����l�!UH��Y	ď�A�������O���R�b��u��њ��=z?��<�5���hI��:z񅾬�4-�G���q|K�۩F{�G".c_����R�b���^�j1˷�03�2��d��aIA�.v��N5��fxE�[���lH���>�ru����'�n����ٗ�����[�W>8��Ԧ�>v�u'R��U�Y&�T��wr��n�����e󸡢&��7Zp
��ښ�'C$va@3��镘�V_���d�E{�5l�E��O��u@�n�O(Ꞷ-���OV3�ԨQz`#�#P�c�:FU8Y���D�&�Qe ݜ�(tʓ���P=�o��#���,^�	�Y��&�9�������M��¼�z��I@*}�^ob�� ��َ��\����t�'�G�h�}�8���4��Nؚc�I�dfp��}��FS���Fh���g�t'���D�"���:�pd�k��]�J�怙8��,.dJ9в����M�Y���r�E�=�;>5K����a����:��˚�W=䱓�ρ;���Ar�O2ޝz�9�"�]`��@�V���y�'���X�n2��������z?��#N��.�Hd�Q�	'��N�ݬ�RN$��ـ�b2�ɘ� c7�6ɤ�)s%= W)K q��Z�>.yF�T�>�{(;Gv<T�.�[#�=ꮩ�m��!}�f�:��s�M����)鼇L/{ɀw�y{ҷ.	-j�y[�p�{���B*��(��E�w*V3 \;�5�U�i��3^CZ9�8 ���;q�J�˷��B8����mN�k��W#�}�=��u�,���k�z1w����"6s�.��g9�k��A1��J�f�}^�:C�
��6Ɵ�Au
,R��Z
)��=�A�s���t�,ي�/s�;���};�����f��2�娬$���'�k�S�G����2;B�s8��Bp"���G�m��[z�}�7獽���W��G"C����������`[aI�f��;�����,�L��f?�m)��ʐ�<	>��v�Y|�Ek����y݁	<6f~+i�&��5���iMȝ��?������b�+Yj�+���iCY'2+� %>��E�&3�iτ
�ٌ�P�Jj�f0R#��" ��!pc���|��tVC^t�|���*�XgS�a�<2�y}!g�툾S(`!p��2=��,����zČt�Qs��E%9^��8�U��!?��aП�`���U������g�:�+�`��kӤ�a��^�f��j�+$k��4�42e�u���\K�Dj���b�o���WLaC^2�0�i-�o�:�<A��7דϦΜh�9R�߮��%~�cE�3����L�Kr�;�>2���?l9B+3J�S��>_��Wd��,��_}�2��캳�?�����|��NAJZ����i0����4W��-}�t�A'yU3i�(��ev���&��c�!��<A'���O����>y_��%51��w*b:��p�d��N�N��w�K��9���A��ּ"�\&����a�٬��A��g_��O�
��n��O���+�3Ω�O���IK�}��rj��C�Ȍ(�3׏HT�=��:����4e��(t�㎡R��R=^+rJ�MK
��5�ܹ��1Aɝ��9ژ��s� ��&�x(툶n�yPo�ue
V"�1�ێ.���d���k��=wq��o����,�&}sh;�S�h��j��~�y��8�ELv3`L%� ��J�v��Q0�P"z�Rf�Þ���\��0)�ʶ_9V�J���ǣ��w��]~�ܡ��Q�w������y�t���r�u��^C�3���d�,����iԣYQ��O8ŹjG�c�\#�p&
Hް��h0���p.�����kF����L �b'-j�a�S��A����aP�NOJ��bHd�ə��}ˌb��Q�V�ӝ0�'�1���s�yeA����5�9Ffl��{:4���7��;������1�أUG��ξ"-�p�x� ]���Ը�.N����
N�����z�%%�8��v�x��Ej�ސ64^OF��(��v��B4��u*ed�>�u�Ő�L �a׫��Z�2rF�	��$#��Q��`Ƿ�(bjm��I��¥�В���&�+��Ɇ�9'�:4�	=	�[�Q��C�t"+�=����ړ1Ol�X�-�m�� �'{ ;0�.� wNO�v0eݱm��b�<e���[�ӳ�v���M��p:���4V��HFW6v8��=�~�Q��>[_߽���.�����^�g�3�78Ol��~����?u�~�O�-��d�Sa�^�F��>c�#�O���u�-Ԯ��d���s�E�}%J'�)���Gl��v��Q��׶�9��2��&gZ<FG���w�4'B�1��4m�&�� 6��y�,+�v`�=(�;�f��"�W��Z�pv����CT$$�$ CP�u�g.�蛝07`���{t���O���P�� ���c�����'F��@[�|꼖A�g�&w�ۓ4<L��u�I���V��C�1ikepE �*F�	��&Hr�����' �!ZZ�mݻ�>�}��e2%@ѡ��r�ܯ���T�����p�]B�Rc��h�S�z�w��}�t�^ݿ]���/:�����˃U�U���Q��lQT�/|:��:f�6�utc���*ZR��ɑ�j�ͺ��Y�lK�MԔ������MC�2
a@����mTX[�������&���:��j�}S;��dq� ED�z��_a+�\)�v�kv�(o���Y=)`ɬUL�XB��.�F&1�ڿ�$��0����k6Vd�J�*cVS�u�z��%600�Z��G-HoH1]!8$���Z��>�:mr� �Q����j� �=�c�Ɋ�X�D��<��鐎8���\1(ejt��j�We��C���&Y�<qO��ѻ�q%yў�[���+��Y�mg�œfd�Q�I�oM���X�]��=�"�-g���z���2�����#c�x�������L��v�mv��#$]�l��k$�׎1��}�����L�U�%H�$_ˍ�Gd!����OSM�@)5W����Ǵ�>4�3��k0��ЖRcw�Y��g4Oו.��(~�Z'"�{
�R���q���W�i���T���EVR�_�f����v���0�B�)߈	��V���f˫c߈ޑr*k�E�Y�i���1�����:;8$/v��@�&���),����������6�8s:H<g�p�񩢉q*d�[��y9�ǌmM.�v�9�"l7q�f��ߌ)���[�G�;�@��cg=t���M��^7�c4۵����}K-���LX6��a��c8solv�}�De�g�S��TH�rt������pv��i*�A�,�t'�?����(Hr�w��� Dnc�Q�*	H`������Pkz������������g��ˇ�j���;������GzY��� ь�7t�cdhd[��L2�kCā�?!Bp�4s�kRq�ñf���?J�^���č���I��ϑ�+��f�I�|�n�[	�	�p�Z�=�~��ՉE�2�d3w�6�v�����8nHO�&/�?gaֈa��&��P��v�����Eɬ�MM ��?ۖgC���Pʁ/s��I8I�,��n��uF�È��(�C/�#�~@���\@z;�N~A1a��X� �e	���RQ�pT�D"NuU3��23��%�$�9	C8T2��ט�X�:}���!���ײ';X�*p��u�1��o &L�����3vet �p2Y\Cj���e����Ȼ��}�7���/֑��6�N|�kԼ˂3�k{�p��-��=;G��*9Qg�D�Zy���~��Q�s�]�Q&&]�����I-��O����e��&2�N�]G���}ŧ�Dx�x�x��Ct"�N����A,�b�9+?����T�tz5�y�b��Nn ���z�Y�nr�B��!���B��&E2���\���\(:{L����(aI�����9#��"yr��ϔB�T�V��I�,\�h��{�x��3����c=0ؓ��!v���%���rm:EoZC�)%���,O�������a��J�CCT��5WN�OE��rm�:bw�k���d�E��5���s����w���x��r��c��$�JUG�z����m��t�Cĳ�=��d}8swv"��ɋ��'�t˥\�Ļ����t�R��R�)��g!�lpE�5EN��рг������%{�g��A �a����Z3Ͱ��">Ǧ�8:���;�{�|u�¡29W��J;��x������_��1_k�/W��o'x�	�!i}L:!rt�A���${R�����2O��4қcL&�O���NG[�;Ϯ�)�qV52�Z���8E�wYu%�}�r�����`����*��T�#ڹ�$���F����9�	�V�&;��>2h-,���$>�1��9�C�u�yO���n��t|�Ӛ�u�g��AM�p�s��[��Fn�1������q���]�]�c�刮5`^w�:=@���ѭ����=�Ω4i8B��S�"+��X�7S'���\A�٬�3���0�ԵT#kӿn}��C^��<��<
�Ʃ��P/$
H���k�Ն�HNN���P�5j��S�#!�!�]P�cf���O��������b�p��	����Ā�����!��ڻى9��Aʻڮ�<ɯ$�a��}��"�D	Y�{ hgA�|jhv�ݽ������ ��8S�����F�V�XA���z�*�x���F��]?}RrKl�X�p�ΧO�C�4'�?j�"��ګ��Ei� �Ivp�Y^h����b�������f�ώ��Ҕ�m�IM-�*��_SO{Zo���x�=�2�|�:iFf�=��22�����1p�=[�3ք๭j@7�&�ȑ(��*�7f�vWgAuc�y��f	J�(���+IEo��h�#��\���(��$8�c���U����`�g%��{*Ji��;��!���8@`F6?�������� B�<vy8��]@Og��洀g���2F�^�O�����>�͔��|�K_��og���ϱ�l@m�-q5��>��Ɇ�����A!z���2��� �u�PuSs����؉H�l��f*�$U:z-�.�GP�|��ܬ꯿���_|���wx�+=+�J;����э|p�K��>A6o�H�rO_Dk��!�7�Y�m*8
3�V�FD�&�I�}�0ٲf��3`�(�Cg�S	���x�X#�f����1��Yk2[My^�ȴ�&�
FD� +6h!�*dP��oX�����S�-d�J���\5�p��N�fQ�JĚ�(�`7��͈$�)ʢa�fI8��͋�zʼd��jnBPalW�nd����_8n�;�܁�r�"A��d����Z�O�<Q/��oY��t�r��'�: �]��A�>���b�xK�P-��!�k�Z����-M2 ��yd���r�4沧��)�{
l��4^��=HNQ���HNl8�K%���m�B�j�[`�<C�5���+)l�������P�LD�A�h����I�VR�����y'ǛО�?K����w�O��e����=�}w�y�\eb�?�J�;C��3{@d����o�0���9���{���C���专pK�Wн��>�gpd� d���>y���-I����R�/I�)c��:4ϓth�I��3��	��l4�ۊT����'���,{:����"Hi��	����5%f����&��x������KZ��b0�g�D�$k��7}�DS���py����-Y�y���2�C�Β,sq1��
��z/�2b��wo@�lk��Wd�)��6]�u~�����M����B7®���.������>�z�-^Am��E����'c��](�֧����wL�����BJTԹ���=HA�A�N�n�&I�پ]^h�*Y6�N�uB�(�|�]h��,��� �/�7�x;	р>!�z��I�Q�O��me�,����K�y��<w�7%�f������[_��R��犕���?�ap��p:��ں]Ԥ<�aTtDd*��B%`*@�+�����#�AjY�-9�9�Qe�w�Iu3�q��%��ĳ q�3v|.O��[;ࠇ���556a�8��^�h��߄0R���`�p�W��	�sd�_���г�͢P��e`*�h�"Yf��H`�V�q�Z%�av���-�5�6a�8'0�JlP�0��џzt��P'W>�rЂ��%��p�;miAS��w�$<��R�:[�s�~ ���X�@}	�l-G4�櫁MjH�A?f�����(UD��^�����	0�Ԟ]��l�k���Sc?d��X�-�k�z1\�TD�$�b&��2��ɹ�	�����1Y�k�ՙX�Y�Q0�#Hd/�:M�f��|'��������X�+�xٖÔ�t�1�˶N��W���UB�<��i=���j��OWÚbr�DD�<7fv�.��3��N9��u˜yF u���x��e�U�b(����h[T�'9��bG���i�B YN��Q.C�vNgr�Q���ᰳ��u��-�=Y3Ĭ|��D�4�K�fܒ���%�`�NЛ�ue�K���:���g'GQ�yk�v�L���/��M\�k�ެ�`6���L�`n�h�dQ��(W ��<n>��J罩�o���f���e�V$c%á�h�4���x\�so��"�-�Wn];�9�(��p�%�n��d��i��s���/���|6GI�3���I2V��H�ʲ�iN�sw�O�>� ��~e���gH&�'��1[�Eݲ}l@�8)���fو Aў��r��[>U����%�HBDX��T&�J���ݿ�3����w������Z�����}t��ş��_�Q(#H�������oh-H3�S櫥��(�-ܾЁqH���(�<$�TU�=V^I��u���L��p�I�ahǑ���&��u>��rgC�*`/o�q56�02N�ut k�M��mV��L#��w4�dv�Juȅ#�����N���F��?ԏ�ٍo��lԍ��nL�+m�g�_d�1�!�?3��	G�Y)��9$����ɖ��ԧ���Or��. �q�3^g���5V���v����EN�CV�܇%�]������A�a�Mi�'9Z���6YAБL3 0�2�
i��$-{�}�� :s�s�{���#��5�(dU7m�P ��ڑ5�xe*g���N;$~�)�y����j`��}�A�$L�H��"{�m�ۍ\���ާ�u�x���e�iV�?�;
^�c�eG���3~��z�w�EK���������ئ��n�g��$&�����o�]FW�M q2��U���T�� &`z3Z��	���|)�E}:c*�g�/h�y��.;����sq��/��{���:�}
�� �E��J;����S�*@|m�-Ig����]�,��,�t�x�43����l�?^�Y E��y�j�/�Ε%'�:Y���!�W�`�U�`��5�Vw�`a�k�9�!�� �;?}#��dȇ�Wl&�e�%�)Z��:�F^��>��P�r7��痹��$�()wF��E����C�!��ሱ#����Up	Եݛ��9�>MMK�ho�~�p.�#U�|M�|$mk f���q�\J%ܹ�S�`Ӟ
����h]&�X��{"����;�V\�V�B3��/�k�e���7��ܡ������;�M���_��dQ�b��ڷ��^9-ON�
1	ߍ�U� S�.īi@X�n�5i�2����!6�t��i��)`cv:�/��s��q[�b�̬{#���	�-�c��Ӊ�>����9pP���8��*�$m�� !G#�]Y�mU�w�a����ԙc�D��y��k3��*>����DB-y��	�	Y����O�ᳲY��4@��v�+���2�9���r����tקU[6{Lߢ�&��\�nG����б���9�1n�V5��{�a�K@UǑ�,�3/s��#�93 &`t��52�vC��1+�:+�|AdّX�w$,��1ȇйG!��Beu�����ڄCR���Y84��Y�Y�5�0�N���"':f���q��V�~�_��":�i-��g��OX������A��:�"Y� �D �H
�T���Bi����g3��}���zS�|�^=!?�?��s�����%�!M7��J0K�̲�6�8�r��E)8ϻWc�̀$ݚ�iQ#hqo����I�EC�1����yA�A��B5�w�ٶ(�bO�
��0�m��+��Z�h�ǳ�a�;�PlB�<�iȏA��O5i��Ndg����E�`"�g��6���ר�Wu�\�d�:�iB�c�SXnp�\�S��3J��h��w1��ݨ��1�jxُ��[Z��S�c<2ŷ<6�%z:|Y?#�7J Dl2����*�D��6�僛G��1��A/7CA��-���B���23��,/(��~���P����@|J94Cv�<��DL��(��heG*WA����A��x���'*��YI-�s^�#������C�3C�� �S�Q��'$hǌ�y�m���&� �Qy4�q�����\Nj_���ɟ���ݟ�Uv�͕����G��GNg��/ݪU��Ed;���j8BE��p|�)�O�bf�2֍��Hsץ;Uk��&��љ�!^b�������0
���c(tS]��1�tIXn����3��z�Ԃ&�1�;�5��� !���i�(��C���60.Y�nG~'f��#j��H�.�
�13�!25C�n-X���E�k�ʢ!IQ��Ϛ�xn�jomf�W�n� {����f?��:����A7�Rv�UvSX�z���P���2f;np8���Am!F#��G�n%tA)�O�4!�.? -��������K�\�Ym�Z[s�/	P����b�.�[��9�C��k�٥�$�u�o�6סg@�����8�ZY����ш��R�g��P��hqs�d�aF��2�p �,�WɈi�8��E@��Sb`i�����fAO�{d
1"z�����x��
�Ykr��zx��ݵ<q�q��K��v3�s<�wMYy��x�~�:�A��,��x���>d���=&�%ޭZ�<f�����`B+d��w����������3� �j�$�9�Sq��|�cc��p
����O��:4���=���3�nY�,�R�w�D�V�uT����P���9���(�"���pL�Ƀ�	tq>�>�@K�l�}�f9��h��������}�N?��5+���i���&)W��$X���u����+ӫ�ŞeG��׎�������d�z��=�S7�9��Bƶ�� ��ވ��Zư1��XL+�4>r��-�N�QQ#�hc�Z-������{0���{�K'½��h����B��/u�U�4����oI'f�
_@-�	x|f烔��Z��Lj������?�Y���K������ϯ�����l�aV�KΓ%Gm,\�O#e��{�Ń�A�b��ѡ5SI3���m&dյ
-i�ߔ���&$�C�_��^Blw��{,"�7X�ϙߒ�(�Qg_��;��!I+),f![�wd)�ؚ�0T��V�,L��AƄ&7g��5�*<�HJ>���M���	�� !K���u?�|G6a;��&����4Y���y���W���w�0̐Z9�!�l����VVe	xJ�6�IT��E��s���8�#mާM�p�$���:�f��M�B>!+���r#"���2�4:�րKW9/׃���"X9�-�;2�]�"D��j��-}��B��ze�����J#}���x��ܩ>�V�sѹ� ?���^�������{�`�w�=���d�[@��+�����bw'��'y������O�Xd�:�ٮԦ��D��^ظ�f�^��c���.K�� ��P�+[Ia[{���C_/�[��\|���N���3����H2kBN�@�c1��A�tx��:�F�(����'�����$ꩊ���J �rD�@P��"1�4L$R����!hɵ@��$ҕ9��1e����}��fBr�G8�%ل�S&{���A�BG^�D�=�*d���>om7�9ڱF�FY>p�� �:� �Y��Ӂ�sk�q�����.��9�-z���\+�0L �\�l�D�L����Y��ýܠ?#X8#��L�AA��(��a�/�����E��@o4���������2�i�A]|��� ��sk�Ա��V-�������O����}���w^9�i��WB�
���؞��>5[��g����ho�'��(���!��*�:�����7:�������
�\���޲�����9���&}T���Y�;���	�#�9�A�$j+0���q"&��,8�:ɏuq[Cd���<�]CG^V����k�?JlF���uy@��K���fm 9�� �P�=�}���R��ĮW�����8�6��,w� ��I��
[ɠj�w�H�#;Oy�3�gdY��xX�[f�UP	CS�0X%k[���Bq�du�1o�`E8���AvS�uH 0V�-2�_K(�X��s��t�2��Z��8���k
�D�{D흈�iw�sh�.��FN��� �Q�:/���!�M�,<��E=-!1�Ev�ZQ/�<r��_�t�����"���,#�^XU��G��:��Z�>u��*��0I
�:�3�4m���}jl�����UсȆv�u2�O l���޵ze&&�%�A�/�2�Ȝ�.��dc��$gr��x�����?!ߚ����_1��o�B�<�Z~�}zl�>ɂS϶�e�7p֐iZ`�:�Z��FQ�mYO���Id�fvL�R�?w�zV��/(V�η�O��4،T��g;��R�rR�^j���J�,�K�&�+[��e_��H�ø�$����bRk�D "I�1��rj�)k��4Q'�i�2�I����y���3QAh�̬��kp�젙�Z˵�i7��m�tT�AN��"gx>@�����y�����麋MLyM�l׭���H1E��p����~��V}}o�ɦ��t	uW��M���f����$�uB'c'�E�o�N��U�a@v_�u�m7��`�κ�H5���u���T� ��jbg�B��F�?`?@$T�g5�F:����&8���<�.�%U(������ᣟ���z����썞�+������Nz?����-{?�VD��v�Yk��m!�Cڰ!$).��yH����K�e��qI-�Z@�s��c�6y}6>� ���D��i���^U/ju4�P��������Z�qlG0�9x��a#�=���C�����ب[�Q�d�[	e
�p�r쪬J<݊ͯV|�B��ڍ�ϭ��\SYUҌӴB%��*a�f+`�5/^�N�F�d�5�kF�B�m�������E_���� ��I�#���L�BK��'ĘN��e�ڎ�5�X�f�u @�b����cTE(��U�F�䔖�s���� {5Q�F�i�aM�l���'"=~n�z �Q�H$�X�������[c���,ܬ\K�9rk'�:Py"�h�m1r��
Z�h��5�2�TވS���@ �O1~�C��Չ�]�e�	ى�+�/}��1%?�:.vl�,	��?ߕYR��WF������S�~�dh�~�,���	=Ȯ-�)9��|"*��
�L� M���C��(\�pK���O���>s�I�5����h1�i"[
,��ڋ����*s��mb7�=�>�u�|+o��H�e�� �:��'�zs3m�,�hy�F��~
��[�\l�2� ��1��n�k��j����=g9�g9�v������ ���NK�t�����w�*и"5"`�,`�,#�n8��C�x=�� ����B/�Z��_'��Je���%�RG @�bp
�	�(׫B����``792ںd	NP��j+(D����?��8�w�T�x2�5�;��,v���S���u;<4�V�9v��k���"XQk3*k�#�~o���ٹ��<�Q��������Y7��'�3I��8yl���OYj%��c�$�1��ֻ���%��)k���;c�EG�}�Kq���z���������<vy�s��1��G���]����T��<d7٫̂��Z�FU)m�^��ο�)Kf�����R����G$�f5���(�?eA��`1�'�X�f"\D��� �mnD�}����~�E���޳Q�7�J��*���ސqx�&º�"X�c�e2z����.�$em6 J��ɨ�-��|�z�l�=�y��M��D�j@�k-�;��S���֩ ����(�8��0Z2mM�$��lL�h�]�${�bP�0j�c�]��6�kZ���!���i����� l��}F��@��`bVό�-u5���tչl�q2Z��gm[T�1���%�6<�sif�IAlK�ܮE,ՠ�"���Lh	yr&zbF�~Z2��5�]1����L���^�\�*�i/��x����(K�љ�m`�����:��t�Os�4�"���&}�׈E�����ݟ,�G|��d�zD�O�`)����}�>C\&�A��v5jBNRvo�j^��4�ҡ{��@��YX�nV��9�46�eH�'ϵUoo��ۜ��^��V�Ȟ�6ͤq Y>Y�2C��r�M�D�L"�cυZ���(��e��/Fa�]�A���Quѿo@��f��q��\�%f.d���q
 ��=FB���^�Ee�4�(I��@��H��Ԟ���ڶ�vj��:�&��8�R���:>+�<|��Sژ��2:p�"�}^������s�Ĩ�zCNN?:.�΀�/�c��*���I�m����S�ĕ�F������&�l$X;Z�gw_K�m
��win���>�$'Dܮ?RA�xa�<AjNheT|�S��h�#��P.�A��Me΄�%�dp7,��������ǅ��DܘRh�%x��O�y��?�P}�?�R���M����e:/�j�[�0C@Y� (IV�
�����M�3v|w�����<J3��)`"F�F�>c�N�M�B�J����V5�cH�?��Wg���^����V��Qޢb�r\�lNzQg�\�y����5�:��l��FN��0r�����48q�qd{"F���<�>7��73O6��ɱ�$*mf�$�7�NG6`&�K�
�Q:�NcB�b��چ���|�3��<�0xb����9d�Ys��%X���)n�y��l��~ԩ��I��~o�V�d4��/q���0�g@g D�F�:�*F���e1��p���!N~�g�.
�$8v�!נ9���`&�����D4%]��G8�J�h��soO�c�e���o�3�q������%�gjiJ���Y6qLshR�Ip�w�1��S�M�\�[�CN��;�m�e���:��!8�A��yďCS�����>ɴ���I�X�]&�[D�8�f�#�=%ƹ	JOjz��dmSk����K���ݠ6�ꕌv��#XpQ%����0�W�����x/%K���5L�HyƬ��HSF�Ï��Rm԰9dx�[Y輨�t�ۢT5T�b��dU=B�i�+f�:�`q�b�uəX��I��Ptt�m2��g�Y�$Ww�Rw��u�.��N)8�Z��4FR��r�f[���'�"ט�cv�D,H���[�ӏ^V5.J#ik�TA�yk���Ѡ-+���<~�-��_�&ZK��2��r��7A�$@���@�2�BtDgi	mD�=�Nm� @𿊘���p�
����GӮ�:aо���z,΀D���d�y�&�7�2�l�w 'bi����앶�=�m6��������}�j�������� ���
��dU{靻?�{&o��[�+E��R���y��t�ӥR��	Z ��{���IŤ!u��֩T�#�7U���؀d�]��9���$z����XH|���`��&F�nk��<~��;~Oi9��zɆ����&�I���p�l �Ld\:���وmq���n�hmoC&�-��<�E��?�Zּ�0�l4�����l���'����ae�9���`�Xqb�� �RZU�N����9�Zn��A2��G�����:�mFYa;1��U�<F]砷J��M�����K�����|=�ꌩk�0�\BԉC����7�p�|X*�	�� hi��kl�խ��x��\��W�`�"�r8y���*�β�D�Iu��<����J���w�ѬQ�2������4�͠I�#9�ȲutOk�)3�*~�@�ps\K�L�n��-����+e�O�xV`y��w���cy�`W?��g�{Z�!=���;�l��P�6��gĵ�糏ߡ��5�x,�H��W�T���p�֔�h&6r��E`�<P�p�Q�d?X����ި ���b��JR�P[Z��V�ǻ|^�yk�x8���"v���8�C�NY1Kĺ��3�3��їP�Y5k�Y��4��BP�t>|
6���{�"�����{�;��a�(���I����Lvp�uJX��EY%��$B��X%��쎅�=ϭ@�R����V������`�[�.b�AM��cd�l.o�Y�@R�񁻐㦖�x�r��	��	�X�2��"��}�rzm��G�g����*�H��Dt��^!x5�	����]2�����skt��_�A����G)3�"�m�-l$6��5�7�n���톢�7QXp=��lV����ǈ�%�x��\��GP�(��k��"F4ݴ�O.{_��h�?���c���]�;�S~a����[��[8m�Ȋ�N�H3t!C|c��*�I^WmV��q�ʒ!�#���������+��Jj�2ؾD���k8���%��
��W��i���Sy��U��W�vnz>�=�Mr{�ʷa�����6�1qT|[Q�o� �N�M����B↊��p$~��f�ёf� �@��߅���A�È�,q��Rf߈LC��d��� �k�W���(�8����q��2��
��2�Xl�w�avdc��\��u�z�mnk9"H!p�=�������	�~ɡ֡�U�|���4a�tؔ��3���\��ۀ�A5Q��,u�}�|��Y���*5b�w8#WՀN'��L*44ד#	��Y�W���݇x�D��VŸr���g�a�ִ��$�pWJ�6G�� se�,���q�Ę�{yY=��r�?|�D'�gIu{�ޓ�����8g��ٷF�@��Gg$������k'����}�d�'������w���O�'��|����dìԐA��*{����Bd�־E_
�#4� ��1>E]p�J.���Þ��k݊ !z�-�	�r� vF:AQ��2�����C�%lG�g3�Hrq/ҢƟ޾P��̹?u�z���L���j�[��q��Z��
z(���
�W1�}[�˸�L�}�c,1�Q�DW`/X�rRcRN��ݸ6�h�b^G���R��}��ans>��$;o�b�tƒ�C�W�r̜2�Α$�xs�B�E^ۀ��������k���q'x"��m�c�Z*��D�_���(ț&{��N1ԑ��Ms:��7����еQoR���fr�1�`S2e�ǌ�@�����x����������O��W+C?��&�k�F�&k�,$+�guc7���?����D�,�V]��ߛц[��P�C��e���������$$ZU�Nh*ʄSBvhKK�w8"��8����
�\	1��j/w����H�M�\�ܾ�ˋ�lV�R��>: �]�[-�m1�Q�F�\�Kr@ɹ%U���g�͎-d�3�8��MXa�R�ʻ)�;f'�����a�8B02���<�$�WB��73�ř�Kt��V,g�����.Qy� GU'���pF�� ������dF���
������D��yX�(�^�ڏL2�r�4sE����oL�㠧�����n�g�!�|�r[�R����C0C
�M3p3���o���*�} ��a�8�O�l��f �}��6�ʋ�:#Y�czz�;-���Lb�k��(>߬���$���������Խ�g���A	�9�q��3e6���x��S����Y�Aiz�g���'j�f���w2E���J;��V��C��Oܵ�'$�)�K������L!�����ޅCM�FYG���t�,s�7�+�j9��H	�``���U�=j�(�������l�g0c��H��'�_beS�s����,�P�T�Ff�Z&�&%$>������S�\(�@�jW�ɹu�Ẑ��C��˺�����G�qQ� ���|�$� ���/z��΢U��aB[hIxI�^1�!��e��Lg^�ֵq�m�d��� ����|��^G o�}@@1�м����d�=<w��,����肹�B9ۃ}6�6c��]��] (5t�����^�,�پ���.5ʠ.�6�1� S��M$�$|@iB{����5������i��{w�W���bMBX�W���;���K��������2���Q���{�!BJ9�+�:9�޸��G�ɑ}��0��謋o=���$�`���v�d�����cYB	q���'nT���;�%���@A��8؃�
U5�����%ؽ�>#�B� �h]�>u�RB���R�jOܭʕm1�e��N��4�s9��kZ�OZ�a��?5�;E-O_�'K�k�k�j�q]����G��� >�H#��=�Cy�)i��^�R~���
1���Km�w���rG��{�c��
\}��9����i��NV>S�B~�DA����CN@�b��eP�Y2ӄڡ�-���W�W�e��pv2���w_�Hl�*��T;�' �̉�[��j��]�h�W8�T���Abx��Ug���Ś�4?����^g�g�����#hH863V�Q�w0֓����w���������?��#!�7�
���/i7�v0����B��S�bKeT��Zw��]��c,�D��~58v���q�uY:�2�{?H�|�� d������jP����e�R����= ꡝ����55�:H�S"Gj��zt
��5�צe�-#��F"<�GJf�r5 ��
��<������:%P�����L\d������Ն�F�N2S����1��>�״We�#��W���X��9%�)5�f�~s�bp�v�	�&d�&�іF��u���v�XhR�6Î�pEȩ��SZ�Bo�[L���(�e���-*��W�i��y �Ah�q�f�{HB�l'��'z~1%��F��pm-%��:fE�8�e�^;�$<��rG��s�.��k�b���a|ϰ�}I)epǚ��O9Ab[�x�g�r�]����Ry� ���2�s����v�T�SF�	���"��9t�`�d�.=���������;wϿ�g^<��7<���ve�`�n?�^[�je<��;�H������V$9�[C �v�P�J����S��7��jܼ5Q�HY�RL)�N��|���qH��>iC��ѵ������@E˖ƘH� h���v�T�l�u����dyt>���&8�1mP�a�ǉ��Y�CV
ԧ�Y�s� �gg������f4�Ѩŉ�J/����&����l����v�S��w�ǲxs{jE=t����3�ѫ@T�ﲠID��!8�s���8�n�wo�-h���%m,�i�O�?!�^,���$�O�GԴ��dAҚ���{8�x,KY�j�̍�%ڦ0�NTV:��l}܀EB>ъ�� k���֢������
RCZ�2�:��t1H�s6��������u�*�y��3���]�K�&�D��	�g1����)�'I'��K�� �Z���V��=�+�!Y������2Dj�{�����G��0鱧v��C�����,Wfb�eӌn֑�ƭN�%�o~�,l[�x��$(<@r�Wf��Lg�Q*��f|�����Ù�y��v��LQo�+��m�n�^{���S�Iy�l�Ϻ�1��?�^q��?78��~�@�
�%}}����lŽ�Ϭ��#Ց j6GY��8+ ��kkp&ؒ@�d�s��(	u@u.4(A6K���SC�z��1��yܒ�"��&�񹓔��5C����(�µ�Ù(���$F�OૼjHa���_/E2�Q' :�U-ԁH�G�C���X8B����D��ZvÖQ�OS�jP��kopb%�⑍�"3J��3����mD&l��hZՔ��>r?0>����K*��Rn�F���Mt>d���?9]4�8c�Æ#�(	�J#WB��kb��V����t�C eIP����I�$�|��
��!�j������kLD=X7��d[��ذ��v$<�k1�06����+�{[�(<w�?��V������:7�,e���p��19i����� ���C� Þ�Q�;��F��j
|�����D8�X�P�,*&�̅��X�Rk+;�id�ל�d;��)Oh �0�O��v����7�n���Q�G薗948A�u�5}��.U����9a�罔��lr��5?��(?F������zR����)���}�����0��s�k�"J��08���b5��BJ���KZ�L�T�jC.<R���O��Ҡj_�ǜ��((1}��Nzva����Bd����9�Q!1&��4�B��� ��0�!�!�=T_��<K���{�k6#�����Ф�k06�Ra��^7+����l����b��9�H�U������6��E�K��RM�X�Yq��&���AdFz9��A���p\gMӿY���6��¼Q:��J����J�p�O������vN9��d��3�r<��կ�2}��L4u?��ߦ����_R�ע�QM<��!�m�-L5շ�#�w(q����\X�HʌuΘ�xN���9������O/S���l!\�k�$����e�׳���u��h�1gpx4�#����֒�k|�R-I3���g�P"h�5 a[�'��3.����8e��g���{��.h�rja�:w2%he�7���Wn�~��]�:f�SN𽃧�k+���>�3
��SZ�S�:��}<k��B��������j<y�9�|ɹ�q��\��������K�'��@P�oV�N�)��N����S�x���B����T�d+=JZ/��E����5�����&̮�k���e�o�ڜ߆h���؀>uw���F�r��g-U�K�4A/ȇY=]�h�b6�1��0�1z�y�{�q��2y!xZ��Aǽđs�#�w=�QC�0��(ߌg�^���6T����y�o�]��+���f�ڰ?E�e�@+���M�C�?mIq�P�A8�N�r� �����aʊ:@S{{d�� �$�,�!�����ZJ���0�*7�mo�Fn1��T�0���?���T�����k���8�$r�)��s�G=��"���乐�1/ᑄ�`��nZE�&WF��v$~��`CQ�����h,+>�sB�)g��(�^7� �*Z��أ�������~?9~�6�~����O$M;�$C?�;���`�;�%e��"6�K���kG#���5E��%�߫�mM<�!�|���D����,�C^��)
�+�+��n:`��ѳf�Q>���Dg����̗�>�2�Z
�:�R�(��*�?�q�q�d_N���:#w��
� W�z�+�8Qt�zi�j?˞Vy+*��k#"u�#��� �R��aQ�)������ǡ���T�Ra5��"¶-��!���Oo"���Y9�_r��C
?��?��G�/�Uw<ޖ:�"�	��#�6�������b nܘf���x�K85�Q�2�D��LC�:�V�ڨN ���C���C#�
Z�w�i��b�GE��-m�Ϡ�P�$3�h�'�N\P{�Y0�7x`ilir�B,k�����U�ң�JP�5J ¤�8�Q��?�r���>�z�-?!F��N|E�G�(q���B�q�&�6�/��h�"ZC�tQF�M�C�tk�귓-�|���Bh8���i���%�
=���aR��o�F�#�Uާ1��1��&�ϱ��h�������*l��dZr!�޸���><�Mz��:cс-"$& A���o���Qі��ǹ��n\�?!�؟���}n�a+��$4ȴJ/+}��A� ��d<߲��֗p�(���FHi�-+o���$Q9bL�QBc�.���kd�����	�9���c�/8��G�l{�I�.#l��(I
���S2��5M�L{��ñ(MV��ݏ^{w0�Վ"���וq���_WnUj�Rv�E�q7��p �]b��*g���Kn�s�f�s����f-��^'���ɘS6؜(tF�X���q@�^P6�� �:�( K�4�aas��F��ڍ��uG��9 7ma3��8����&H��&�ˬ4�ǸT$�E/�A�&��3�5wgSe~�}��2����4�]2�c����qHa�t4��i}����:�_3�5a��22�!&f� ���MhEӛj�b�m�.4��:v�M d�v�p�p�T�.�ޏ�~AX�|���o=H@fb�A��.�d8f���03�[H^�F�d�r[�J�z��8��O�#�g�D�Nr�<Rߢ��~W�pEZ�x5�& k�e���8�+���@���=�f���ȃ��ՙ%�,�Wn�k��Fj�S�=kDc<�p*���@��Dv��b@Cm��bk��z�?&��̫����\2�s^�z�z��V+^��D�3��1�H�Z�6�T+�v�0ࡲ���K���&ym*@J�sI�h�"�cD�Ƴ��#�O~�M���0���W`�m	$�Ĉ��p8�!>����p-��ԇ�g����m�:�M�~�O�2������ �:��Qv�� 4d�F�PP?Qa2����H(S�G�<zk��h�4�4��'��A��?�5�gE�y� q��b�8a-';���3��#+�>P �dB "��b�H��_�&שsƝ�������Z+r�HUA��K*Q$x\���1S���E���6��3�2��#��I�"���uq֢Tul��L3ZH���hM���\CF��~
���2�V��wR�f��@��֯���ޙ�v�d�A ��8c��1���~��;���LNNl�����y:�DE6l"�3kj�A��@{H���E 6����F�a���F�2����фL��sk]�R�P��ER����v;��	6�z����*vMN�A��q��eg@ckB2��@�r#J���k-*asF����^�jR��kWǡÆ�C_���s7m�h��|5���l�d.ڮ��gִT�#J	ϸ)p6���CAbV�v�	��KH$�ǥ��
G���xԬ�Y3JL�S����Dx�
o�
pt���qڂ\�s�8�Gz�2��\k�kY<;aT��6����LDC����JnzM:al�=|��C���0�E�hXJ�A���H�ssF�ʛV��F�ϋ_1��l��]�s��;k����Ug-D&;�B�tbϩ�nF��\���䡨���$&�V��D&�4{�5�Bz
�m9j���^Sȇ��P�w��yK�_��:�)21Ά5$�=��.����U�sBHF}vJ�Q��*4���dd��C�!��ƾ���T�J*�0�B? 4�s�̓�K�i�Z�0p9&����|8��7#>Ӱ��_��˳F�z�l�{�9�t�}����]o��چ�ҦΜ�z3�B5kE��c��W�/������y�Om�R:o����p0+���rQ�,W���������ɽύ'�#�:��x��.7�N��'�5���ν��Qe�o���Xچ4C�7<��Y�7��q�@ؐ�-q��e�vJ�h��e<����*ޚW!��\�-�&j�ؑt��|�Kws���(YV�^'��S�<� �@�����ʛb9y��h0+��Ӱ�?�2���<x�5oy$1�"�1!=�S�
��$������C�6zڊڐ��|2�FG� �1�\��`>���X��sޕi�(��ݹ�A�%���dN�����% 3k���>z�d��8L�*]���c8��1�Hy��~�5y^yM�Տ�!*_�0D��ͤ͠�O���>&�8����оI+5���E������,�R���'4��R���E��4CFK�Sq��v��8����[����h�K�����6&�f�΀H�{�TkLW����Q������ٰ���8!�����b�j��l�Wèm� q��rI#�qHDQ�'I:E6}t��"X0_D�3�l�����/:̅��!�Kr�1�����qFn4�|��CEDU�#��c.#�`���ȕ(�+��~�K%`y-A�4�Z�a���	A���p�&���jY fr�B*A��BƘB(#��!���H	Sf�>>db��*���S� �	]C�&X�>F}w��8DCU��ѣ6�g�{D�s޸YQB]�q����w��ܵ�|dF�Q�LG>��E��������q�f�B��v�J�%y���Ѡk�\�	��%��Ȃ{9���y4���B7#㹶N�3sb)e����)�[Bh�w��ڎ8��k�"%k�
�x��+n���jJ�Ţ�[�{����x@�n�z�к{�_���z|���k��A�6g.ڝ�
�풬{�>��z��G��S{�ӌ�������6��$*������ᇽ������rz}8>�y:��>��m�Y(t�����m�PlwV�bmX:$�5�O#Xd܅�{K@hI���p:�%�kѭ�����ek�[ |��W`� g����$��A1.� �y �"��a_ـ9�0���aB�[�lh0O �P?��1�4�K��7[�*d��D�`_�m�Ir�e��͗��cD-�9�x�c�Ǩ�f0Х��g���@�li�Mx��P�M�,AQJk�e�~�򜪦cgpRsW;9�IgT%������HX��?:T��$���
��Cƚ�U��S�sM��	�ؖ��y�����!	[r��B��|tU#� �Z�p][�$��f8�h���%Υ�t��� �n�>���׉�դN	�['N�Β@_�nzwdJȏ&(�pM#%s-� ��I���x�j�?^^�wr)<p%��L��h>���D���Q[��z�rs�q8
PxX�Ȅ���{���lB!��R ���^�
S��ݹs3�)^TΜ�3�8UF���Z1�u�e^;|!Fq"�*�T+�U(��ʓ�a:���xF��=ER�u���^�|�8.�@VYX��(�� ��00d��d�bK�tʈ���D{ǐn�^a��A3�?��Ň-��5�-�q��%�(#&u&��AO�L(R0��� 5�Fq�p�j2sS�ީ#�TX33h�����Sǀ���$f�� ��҆�r����B���|g�z|c,b����9���$�Le;���_z���&�H���Cg��^��
�Mi	��������8*�b��xh�G��=��^�����e)XC�1�n��������'�v��X^^6��{׎�o߹up��qg��W_�����#����ɮ]�c��]īǰ�b�������k'�Rȶ|��e���O��=x��xZ|��O���|�~w�ǹf$�_��o��6~~?e��w�̃O��)�8;�f��˓�o M��p��H �)/���D�Rf6J��P��^�qv*�M'�lk���Z:�J'ak���c��J�����x�����e*퀽�ڵy\�׮������V!2pj�h�IntyI���K�e�mh�;sl
Ky����1��.sG�>��/\ˍ���X���H��I��>�����S���Jj��굋Rx���{�+V��B�������5ʌ֩'8�����9�Z�;)�ɢ'��:IWԮ�1��.��:�ձ����ލ6C�jwl=�О�)sm�|�U�kB[�jd|+	�f��=e[�6�+��Z�A��@r�?�]=��}�Q\��+��WPw %�e��X��uj��|�ą �,Xٙ� � T�Q�UH�M@�c.P�NVe�z����lz�@glO�IW<�M%ӠU�Vc�)�ʡJKD;�D�(� �!���5�sa� ����E�2,�a�Qc:�C�ՙ��A�٠�F�rIB��C���5n�G�Lz�RF�("o�ѵp`8si�h�?֌�y)�Jq�Ɇ`�5&�w����5wG�3۩ّ$�.�4�ȎS�����Iw����n_uY+�vN�|C,���s����Pt
f�<�����[��d�\40�q &���c�%��s�������|?�kc9Ķsa5u����5^2�	���}9Zg�R�R���%IS��'���7�O����Ճ�fpqԭ������g�vs|�����awI9`��^m])��+bS��.�'������;g�o�������G�Ϋ'�����x����Ѽpm6�/�;�J���R:��-�c=��8S�B��-���	$E�z�8�>�8�~��>�����m�L��ny��(��'B b-p�ځ���:%[]���U̝aJ�K_f��Y?*�hʴ�5-)�� ^�$��ƙX4y�-ә�����a/g��I�[n�4M>��G��[7���ϟ8+�����j���!5�p�*����_�{Nf�`�}��u�ՏAE�f���/��q���g|�P��=MC4V���]���>#�ɔ�{v?�t�9���g��g	MVEj��|���T���J f]$Ӧ�.ڷ4��Q�grμ-op>��'b	�$�eyAؖP�=��&3�/�d>��5�}��2�O�Nl����R#��S�s�|<w�?|�f�m ��-nm	G3uH�ɳ��o'�ئ�f���(���2�9���Fo�m\ֹ���p���)�jN]D9�]6�����{8N��`{��7��s $pE Ɉ�b�q̫Y~��Ȃ$��	�6^+��zg0 ^�תuƖyl�0H�ze[���܉���Հ�/a��RW���������CJ^��j<�A��>[^��)Y� �I[֦� ���4�T�yس����i��)U�'���P��_�;�'�`����� .i4+7Ӑ�VcMyj�우r�X�}�8��;�T����U�AN��=�3�����f�n��(�9�Za��1�εa�Q��EƮ-)�3 ��(�����d���VӋ���޽bi�����
���?��Ͻp�����~��^x���������3��3�r����~�q:�տ��y��Fo��F_x4>{u^(ߨTZǵ���ͪإ��ܮ� �f��UK`��`��z[;�J ͗�8*����g��"`�<�C�(�j�H��QڒJj�'.#o	�FO�\�>����/��94�_����^��2п�9K�ӂ�H��o���f
�QU3H�.+ !���r*'��&ț�Pd���27ũ͗)�����m�S��ߌ>�������aS���Ȼ\�d�=�u�r���݋yl�5�ǈg���T���S�|�|��h��NyhF(sy�5'�p��OCx&���n��G�]Eʎ�9���9����Yu��E$,�'��}��~Z;W�*��v�e[���Ea`���?�ل�i'SPf�0��$xU�wDD��49�[���4��2&%��\�J����wE��L���ȇ�ql�0�"C\'#$,�~Im$�x��;s3���'���hqI�\ҘB(���T��b@�(��םP�oږ��p��RKWՖ&aX�{{A�gq��*��A"��X���Ų�}��X�j�1���";w�=�{��q�Ȁx1F�#@���Q��V�DN���'���Y�D:eU���l.?_���u���6�A�"��\c"��������I��G�o�z��'��
my�X�b@�
S�@�;k� k�c��b2���5jH��ٚ2֩���u�CwԪ�4ِ�砟�[�"H�RZP���u\��)z�3r�x�rȍJZK�';���Nw�2��m+ ���|�ZO.s���|88����wj��ߨ~���7�F/��_�ݜ�ɗ����ʭ�����.���|���~����Ea����k�����hsg���(�^(��G�r���X-���!�#ÐuK�$��"c���Z!�ݠ;�;�{ΕA��P�
b%8���X��H�h�Lv싨��w{������t��s��0&X-��5���"�0�Y� �D�M~������H�~֚	Z�ڠ��fvo�C����gp� +3�u��ܚ+�J9 ��
��"�=cRr���c����9�m�T� �}�3��`�q
��s�4���˹����D[ژ,z��{C�8�:Uk�/@~�ϚyG^T�����#�0��9�"���N,������Ic ��^K�}���߾��#c��$-2r�YTD�a"b��M��!�}��!��Ǆ�R�!�"����CG`�p=�6�s��Z���Шm��ZG��H�X��T0���mc�%Z)!P8h{D�S�f��h���Ё#��ը[�L�0����[yE:z2&<Y�r��,�����JE<����P���oݾP/��&��$��>{��9h��d�%�W=�n���:�2jن�R�[_ظ�����LͰF�Z'h�E��%���	pJG:�QR��J!̤�u�q�X��4����t�ƣe�Lr�{[�8�NU�Ů�z�Ȅ��x��	M�{��L{d�m����%�v��"@o}�%=�DA��	JN�MT0���)���UU�Z�pY_��IsY��"�?x.%2&1/fCȅ�,���vyڮ�u�V�˟z��ݗ^|i���ٯ��s��
ء�K��v������o����ރ~�Ï.�=x����۟��V?3)�V*5o�.�4�����G�����3%��ڲ�Ϫ��0�DJe�\�p�c�H%R�BŲ4G@o�;E}��Q�!7Cƺ%!�Z<�rMȖ��B2���s%I��wE�մ*{۳��93:`Q[8��	�d{�NG:3u:��Cnb��[:�A�C��:6c���!<o}��ǜk褁��=��̓V���bHҔ��U҇O�k����u䉳�,+j{�F���$�]G<����N� %�&1`�o����$5NkU4�T�s��Hh	r���ٜ� �X8Q�fݿ`��!�jz��n1�\��q,�A[��3x��*f�����+}=#�,C����D���z=�.�ٰW���8���5��_Y�b���'ID	:��������*�E��7y?a@�m!8���u1�LG���c�Ǚ�s6�l���9�Q�;�f������=犡D&l9�v9p6tԌ�h�L�;����-WQ��e[����]���:��J�a�́�m+ �"���\֢���&�QsF���-�NIL$AOέ�i~t�.��0/̨"��Y�ލ���|��CW������
2�^F�h�YfrCj���n#YGP���݂���$��:��j(c����!Z�f�11�/'2U �pH���6ر���Zk�?�6�
��q����c �R�J��/�D$�ٓ̽�l(B����z5{�[Ot��Н��Q���W_|���_i�⟸��dd_�3��2�V�_U�)�����{�>xt�{?x4�|��<x������e���{{[n���ܶ�%1�uu&A�L���,;#&�FΈ�L�
I�&��)�<?��M*�9���Tl�	�y���Q5�%I��L�i�����5�_��l�����=�ł�-���KO
���e��i4�η T}�oq�5x2^�A��$��x�]�����>#&���&�*�����piz}�t��p-0������{W��-ȭ��Yȡ�i����q�(������^�3r��u"F�Ҧji�'�:k[̰�"#J�**&��Y��
�ɅZ�A3m�z���,��8�<yr�bL��UG�|��n������(B�����M�7��la���N	�(����<C��3�0k#Cz���#�-=�X�&���'l{m�
xE�&e[q4�r�*E�v�zuxDۚI�c�z�=��J�S�5J)�9hF�U2׼�Z��89)X�R������s�x�^�Ō��2c=��C��*Y�duW��+h���
��O�0��u�:��h\}��:D���ZSsLi�x8��!��T�N�l��Y��#۷.�a�-���=�
 �\��k3��Q�8���k��0��4��G����82��j��k|m۵&~ɵ���q��=�fׯ1E	��ބym�{ЫJB6>��3���R��j���vu�0�_jtR�t�:�z�K�~��K��$E�&ȭ��6N�|������W�{�Ž�˷���~���dY�;���O�X�?��5Zmy�fo���G�����'�w�;�s���g.z��Mf��&�7V�k���A`�9+���lhUd���sX�����-�e9�H��4v�HR5gS�6��NTG�3�Nzk�D�Q�Z8�� �ٌ ��2 ��(U4�:�͹:u��\���o�D}p|H�҆&9e�Wq�2j.�>H��[��p�ɶ�Q��Z0ڭ�)�F�@�}8�@ǹ�pBY�H�CP�Iu�u\�f�'#R6V�	[ef>Pޙ ܾ~�5(T�����"�&k�� m�5�e~h`�I��Q>Xe�Qo
�C��R_�e�w��2��ح��(Mb��L)�8��B�JS;#"�D��,�&Bb\k8~q��w)��1�|]��C�vӗ���9(��6�N,�ϧ�,I5y�ń�u�KpbUe&n����5������h��}s/w����~�H�<Fm�#3S�3 3��� �������f3qkY��+�b0��hh����86
�� �B�FǼ����5�(O���Qac�D�ʖꨭY{}ƅ��P�vb���L����#2�9��!�âxFhd��kF_lb���
�(���e���:5�eΛE��x�Y�$m��7�XH�[*� �����Tq�%֣�Q��8`D�c�,j�$1"�?���C<��6���ˉq0������W#�Ge��a<�&X��j_$W޻(����+�k�����g���Ͻ��;��z��fg��k���_�W���^�%��~�l�὇��������=�����/�,~|�,^G8�V�X?([m�k��9�Q�)��	��]�J��:	"y�\�Egk-V�\��#��h��y�e=�JQ�<�!�%�Tv������&�S��B�C�r����*Nn�����1�=��4���'f�x��f����w�}�첟ۀ&T`Ëޭq�s�t��Z�R��.R�8sJ�����ac��]��K�i��-�	�s:�Pn(BE9�N:W��(�u'f��0�)�D�J��xU� �ltȺ�A�|&�=��M���^D�P�~s����Q�[ �A0�ҹ+W[�sٲ+���&�#�J�1pI�-�H�t�vS%��`�,����ø�%8;ih�a��W�V�"�a�2A�͕��Wơ�Jd����J=�?�D�֑hk��j���otP1Y(����t�@(+)3j[�D-���o1��O�鄳ᥬ�Z�`m��mO���tԲ�\�7P�6�\'�>VQ��j��C'�l�I�AiM�Ċ��)@i�x�}��s�@�=3]������ۧ*7���!�����T��R3
�G2^��&�)a� �r��8V�k�F���錑ٵ��f���գ]]j��B`��˘��B�nb��ٜ�d�{=Kd=�I�bek	�9�0�<w )��V4�^)���B�6$:��1 2�����{aD�o�k�ly9i+�,��cQ����/1f����,���*��?<>���k�u��S?qx��+������;��.�_���7ӱ.~�h���x����u� 5@ʿ������'??�4?�^�Q/��T�����Я���#Y�J��2�+��$����p�pf�f~� ��%ʙ���C�I�1�eΛbO���l���ւ%��GNR�$5\\LP4��N���1Z����1��֘�T�tZ8Yf�k��I=�%ɥ��g~tc]x?I�����v����|ř�^.�r���:p�����Ѿ�89!/,#�a/pc��,'�Δ�˺�p^d��S�k[���Vx}���.�mg�3��x(���/�=�yk�;�,&-	~R�K����=v�*v�Z�ĲG�JdD5OҴ|#���������v���w��\��ZȰ�w]�se:d�� T�(�T��y�.��Ft�,>#z"�-�:���0	}G�"7ad���pe��F���E�e"�kD�J�%����l�C�`l�3��-�Q��Ӷ���W}j����]���`Y+B#��#QX������Z5�u��|n�h�]$2.���O.z1�y��U�bcw���5m#ɌQ++>*��N�W�����������
�����&�+��4:ԗ�З�M(��+��d�+�SG�
�/��-A����"j T�54Y�=��@���ʠ�S��}�=���P%hi?�8$WB��@�UApL�h�2k��<�8�������byv���u�z�^}���?��}����go1������wX��o�!������G�{o��������}���.Ͽ8Y_Zm�/㌮��U�x���������Ԩ�U�&�BK����q�sߣ�'C4xM�_G�e�3Ź�!U�O�Le+�D��8��z588�*�}�{$T'Uh��!�p	����Lc#��J���anqzA�K�����Q��#���5m��S���}>U���l�z�c^#!��b꠷�-�`3��0�pN@���Z���k�����)t��T�_��M���T���	heH�y��y�)$5[	͇��0BX�5� H�v�رd�E�å�f��ðuv���m�l��'J�<vD�ΐ�$�������g�����x���Ʈ�וq�!����fl�)�9�}�Nr��?�&��n6��P��k���љ��3�GN:�H
l>�Xʒ����m�fv�z��	c�4�q����>7�é`��a#�=j+1���T���)@��P��Y:�X,�d�Bf�f�4Ig�D�5{E����M��\wGj�{�'���đ�2�y��llJ���*�a��`������?h��qΡ�^z}����? B�,�8XV�����b}_∅%�z	��l�/A.�P�4������z�8�.��^/S/�g�I�=J}�Q���ǚB6	�tA�s��-� ���1% ��3*�F����[�R��_x��[?�3�~��W˽_z����+b@�c��Og5��ޝ|���ӿ����=��7{�����s��WK���R�ޒֺL%X;n��X�s^��`T,4PvD�֬L�&t�LQ����a̐I��nC�7[�&H�N'bZ��le@ )A�`�<^�N �:���w�h�����b\8^��)=��W?�u�k��������ƴ}��P�H�g>(aW8�@�!@�t�4��:H�]�d��FQ���$�@�!0�P�K�Vr�Fi���a{�AJ��xp��ge�|�1�I�����;�����8y�j՚��O����V���RK�Q"ӟPJ��ɢ�f宱갣��)���j5
Lx"���蓗#��B{��I��L��i�*3��1�r�3�6��?���>M;��{�3��r�&�9��À�%e	�Ԉ���R���d��^d�5 \� �q���f��> ��O�t��)V6���g',6:�s A�!��a��I���掉\n�h�e�s%�(�q�ړlX��~zB��E4C�Y�����zj�<���B��hyF<� 4�Y[v��&BzzO�-��2��SDc�D[疔e����G\�(�?1J�>�AP!���=�P�uψ��8p#Y��*���v3w�v�}�����!"W{��]��?����m����$�1��y��nT�ڹ�@`L����Q��ݝo����?����_��_:���p�W�c��?Ǖ^��~�a�����������sv������w���xY}�h���k{�L6is��"x��p�f���i�@����4�d#z�uVi���9�,�d�jҡo��qc�pQ/���y�@b���s�Oq\1��;]Mn�f1������0W�S�;��q�x~��A��G�{���R���ҥ�Op�����Բ=Z�t�j�O%��0�cۆ=�b3d5r��=�0d(Jr]�������~�c�S7��}51������1E��~�6c<���56�C��co�$�:q��<��'-�2H����E?����&�����q�:�S���G��G� �ܮY�%�JV��������L��mW���#�
ز.����t�Lq���W���㣃�{w�����a# j뽪�M�@�?����Ht+�l���(oj6o{C2r��x��à���\�B
Y#!)��jA�� yyv��w;�ê���)K��	���I�Be(Y�ѱ%-�_r37?��&ￏ�C�J��lLϵ�8N3js��`�_��/��Io��$-ǨJuѭ��d����'���r��M`����8U�^y:u�Ψ�EE+�4Y�پ`�2��B1�f6���&�X�7xp�i�`�MF��a1 g�0�:/����
��Hvk0����!�<AP}���y7W^��#�������廕�����o�؟��O?���ɫ/5z?s�~.�rU������?ѹ�c_�{1����淿����o|��g�>���`�z���R���vS:(ی���(�B���{����}�Kx>:t��G1g>Q���#C^R���o�ξ�h9SsB�G	c#4�H�f7�V������dc��r׺D��؇{q��LމڲdS��3J�Ns.���,n��/� �a�48�-��g��Ӄ�8aν�����Ga_zH�8�4O���7�9r�"v�
� ���Z�.qЪR�ױ�2�.'HtB�2!A�WiN��Y���5����52�!���+8�Q�H�+�O@d'��ML�L�m���_>w��:Gݎ�GDT�� L3�r�2$>�L�32]ue���֢���ťj��DK�!����l���T�ūxA�ZO�G^���dk�J ��r�|���a�c�8��� ���Qi�^~� ���z�A���2T��\�-PZ�uj���0��_��v�����k�A�ѷ�z�m�)8�86G9�Phk�'l"�p�\-۷.� h��Ȭwt��s��0>��G���jd�d��.�C.�bm�p��ǘ�I!��^N0�Wj�,A	� ��!� �5��A.TrEjUե3s�	T��xp�-�wY��'	�ry�aTN��r��m���ȷS���8���D(�r���3ޒ�頲��w�;���_���_��7���Wgw���C���#_�x� �Z.w��������W~��o_��o\����������E���b�{��I��nX�;ɭ��--i�+V%�v��P��'��G0)k�mv8/�%'A�hY�3İ����5���:3��`܏	�y ������G�@p�����N�N�ǌ�b�140��Z�=v!W��� ��@�Q�{�U��oIM�,�5)�;#�5��u	D��)]����6��\R��ڬ�_`3������Sĵa3����y�	��ڎ	�� %�0��VfZ���w���I��_�QqX��;Z�g)��������&e7��wz��̚�{K�\��H��!�w�8l�i/�_��+��"X�++:�.Q��)e��9#Aۢ�M���6��!-��z�+���nݾ�F4SN�Vֳ5j-��fq&7�-�mAr&����ы�V�9;|`L;�(H�X�a��(|_�Q�`�룕r�m,@�D�D���O��`$�x��֬�͚���03m��g4���U �!�=�"F��ȼ�/'½�͍HR�8��x3_^��8Rޯ�b�)ϫ)Fak����*A�ױ�����9G�Q	HE�>���U'�UϩM����x�ݸe�˚y���5����)+�#�M�hF�Wc|�2�_��LP��S�^?]@x[������L���W��/����̋��7nt��Ư�]x~���Q%�����ͻ������o>��}����lr�m�{�a�,*���[�U�A����k�٢q(�znԼ�q�G]ޏ�"�l��%Em�
rDr�D���3�����*��e"�3��7o�:$@�@_R�T�I�|����m���Yb���rl[�׬6D��\��Ǌy� �#�q�K�i�3\��Ę'�m����q�Fԅ�_�.�Z�ϱ��,)� gˬ�@#J��\��s��Ŧ,�sşs~��x=e��M	��o?�h��I��mN��¾M�1��*fq�;ov�4,_�������b=����FgwO�{�K�@%��PT�r��:��睖C��וq��FqE�|��Z�c�17IG�� ����oR"�y�8��w�r�����n���Y�%��N7�O�ٌ%u�ݸ6�A�(����p��f��s=�|� $��i`�N���Ԥ�[������3�F�A�y�����^WH"�'h##�t~�u�嚚�h�Yu�z����f����~����s�c�`�D�K�f:dM��F�������Ff�u��L���-��#H	 ��u�#I�3搏�����!�	�ۢR��4�dED���i��~F�l�`���R�e��x|�2�Z  �a;]��9s�1(Ó�l}٨ξ��?��[��?��7>U8�L�����0ϯ��v~���Ϲ���壯������������d��J���u�y�T�6��I���T�T䫨� ���q4q���EǆR�L�U�ගv���&#c����U�;Q&�G�u��4g��_�N����Qǡ)��Wf�,T�
5+�k�`Ń�E;�>M �}����U��56i�#W�m��gv���R�Y�,뾍=�|�º����͔.3������S�$hK�8rb�P�&O�B)@"�ܺ>��z%fXT���mMǮ���/t�X'����g��)�C�vVRS;D�d�Cb�zg�5�'�ݲ���&ozq��D[7Y=>�K��ą g<�X>��te:m��Cg�����3��w�-�u9�%��yai��b,��v�Z���߃�x�s%�R%�!�\hI�T�3�\H��Q���Y!�b���w�(�@௽t#z8�]=��9�v)���1���9�9���]��j-:��ټ�F�LF�F�A�q�|�h�c�(s�BUnʮ����ԪgҴ��T����`N{L�S_�g�`{�9(� ��&�F*��y([�!0�#�RƯ�Y��Q���|���<T}F����CP����&Bi	���S��-��m��:O��Q��W�2ZE�1m�!i��9KQ�ҵ�Es���F�?j�W���7��/��/��K/W�������+��
|�vy���l�������}�������毬f�ۍ�R�����Y�Ru�C�ZiQ�s�m��'�tDq��)c�<�{@�f�C�Pz���8�lu�R���J�OO9��H�ȧ�`kV���1n/ ~-�cNEUw<<�b�'�'����}p��JxZ��6B���)�ڡtx��=�}��S���X�v�J<;\�O2ћS�����g2��R�X���Th8!�;�ef��� G�ڶ���o�Ơ��gR�ݭ���ѱt!�:��+�AISQ�4�\� PP�%��a]�$8ʌ�F�D��\-uP-���o^?|\*Z��_WơCR=!�D�W����bK[����zl��}������G@%d��L�I�B`_r�0�����Z��9����~m��zD��6�Ă#|��!���Gg����F��V�9�h�0�Ж*M0�vE�éŰ�Lz6F������pm
A;�T@����p�L�^��e��K3�+LN*��s�5�8��{Ѐ�A��8�uވ��Iy3�
y��Pw��m�9hm��q~�N	��3�ʆo�B�:l�D��Q����YU�X��C���y�.�
F�kb���v{��Kw��s?�������ݯ~�FU����+��
����������������>�����3���b��B�P=�.�t�%�J c9�,X����(�
�ކ--#Pf�Uބ���B ����M&�]��Q���y"b8�9��2æ��Op�+��)YPZ��>��>]6p��u�/D�|��r�h��d&�r����Mݞ`ݶ�}P�Cj��d���l�i
io
"���)�R� 
��л"NՏ�	$B��OM�4�� }X�H� ��H��-� �R�$k���k�3�������tJѬд��%�4�1��u1�6es=I�z��Q��$>��R�Z���ȺU��_�y��tB���2=?_����^mu�YB�V.��=�k�Z�>;lRQ�-Ԟ�W��K��~�anH�^��d�ͼB2�od�f�FU�P�g�n_$���UZ��n�PL�����>������{�AYV&�(,Æ^q8�:��E�.[.֩;�Tt���G��u�+���m��a�F�����3��&?��j�>mJ�:�i}���S��=`S7�d](t��3�Q�z6�����:%�\Ӣ~|�W��9m*u��� �jor��'=�4���ɼ��əY�\����0C�o����\�k��l�����3HvΏ�U��f:Z�z�����{���������{��OWd�?���+��s��\����'�k_����叾����?6X�d���4�j_��n� �?0S��i��z
|<�a� ����Qk�p�ʜ���2���Z�����y���j`$G:�ݮH5$<�+��dT �q�Q�8b�1� ��;�]BhF�F�g��+?P���_H����PZl����)�V�A�ҖZ���u��31�blK$:8I}�f�r��]Kd��-�u� �s�9R��!ΚN�ב�s]j�N�tl,�V�[#�	_����6����2D=��q����N;M[[�o�ȶ����M��h%��
s�C4��Fk���*A���^�˵qq{]����2����D�ԸX"��'�)f�����P�X�W��4�x����^Dk�ځH��*J��w�C(E�^x	ߔ�d�ҟ�m�6*�(~Pq0u��O�r�%~Tu(6/�EL���zD�D��&ׂ�v�ړ�I��"����r�W^ը/b<�H��܈�O�O=�ɼ��,�Z��8��s���{SmQ%��\d����n�� w1D�A 2���7|�`c+0QWJ�:ʵp���<�f���zC1�5)	����~B�S١�­����2j-�V���;�'�����M����o��O���������߬`*�=_�?^+��J�7OWg_�����K���7p��)���Խ3̷
+�Y�M�s���"j� fꈓl,��
�-am����;����	� �2�y��2���gG$r)s���l�|m�mË��-t���ހ���̋���HdKj��ػC'��:P<�Z�T���u�w�aL#��	�^	T��ͮB���,�e��ɐ�~C�Ub.���eW���W~��{���J���gW�к|{���H[�B>�e�n?�"1"�N�3��0�G���8��n�#��f⾏eπ ����0{��J����
}]�~����*_ا�=Mhﳍ�l�)��5mл�,ۣ�8k�c�2n����>�́~�-hܴ�D��n�;\�<�tEOwd�D��_tv�y�y6)R~�uʯ�x�CG���(Nm_ v�_g��D����W��d�/l��+����e΅*�9��LlD��m+J8;Xb��yƐ'8�9���r��c7g&e(����iI�pXzԂ��<FD c6���v|�M+Hn�
{0��)� �{�B�u7����vc���X��}z[;t+B�Nd�5���5��nW���{/�������?�՟�u�g>3��=_�?�+�㒭����hy������������{��/�*�����SF\"���d�S�ep 3�.�3���8w�Ԥ%����A�����C>��[� ^l�*aG
�%��Z7Нd�6A����K),:ʠ��Ճd��W�PuȮ=C.���w�z%��
�\v9:����J�j?*�ː�J�Ř���t�Zq�9&�r!���,�^6�D�`kE��ʓ3w�6:`v7��l��.Em���'��R%K[�]9gE�V5J�9/.��P�6t�jE�^���d�;!������R��a���sٯ��߽��C��'������J�z���)�A_���+j ܠ9��Z�2�E��7����6r/޹�����ZO�zl_���,7ll[?����S��c^���$�YǢ���j���~g3��Mm��oA�����IX��X�&
v8� �A��m+�n^�H{/dfl?C��E��yv��]�P��8S�;����6;�V$k�!#�h�X�@b�P���lM��ڑ-o"���3�i-�q�y�cz:/��u�nx���2�1J,9ü�G4�5%JFC'w���9}���'لu���T��F������g�E�~�0������/���~��'�=�?��6��?����W���)�}�d��/�O��?y��{����\��Z�y����H�r�ȦJ�/೔��v�a�����AѦ}Ԃ���S�.��6�y%��,Aek[��QNkwзP܅�@TS�RDX�d	{+�}N�$��(�.:�`�cC�8˃5r�a�!�bfBˣMf�Dv	G�s/��Kj�=2�!Lzu;���:��T�7�b$@���W��50�f�U�_%�@f7�k�(v�����{g�`��Yy�k21�� �5l��Zu���5>w��"Y�W�y/44H�D]K%G����<I���-���HW؃.	�Zju?x����O;_7�
��J8��{�y�[��j�6$p͉�O���I
� 	��I�%�ܔ

:H�d���-2�r�.ٴ-j*J��y��e�$����C�����%C�����
X���\��dS��A+{��&�Y�,�_�M��&��=\`��dp���4��!XB�W����<�`����ۊa6�Mxcc��� ���D�cg��NU��r�%�W��%g�t�n��!,c�[�,�Csr�d��MJ	3t��Ӓ�D�/qX�_���F��u9fC�>�	�gj˺W���7珋���v��?��?����/���~�F�	Ͽ������V�ǯ�'����_��k�������_B��O���o,p䪨eR�xV��z5&L��&S��y��I%�Ji�V��
\��i��Uk �8q����P�$1H������ �Z�;�$c�].JkE���t?��ߚ"��֓��׼��ϗ��'t��٧r$J�:Kht�"�v���p� ��Mˡ���/��$y�g*-Gy'�]�m�d��y���QF�33� �+����;eY�t�c�a+خ��4�1��*~$ƫڑD�P"1r�K��7;7_���Ko2�@H�ʖ����Ѳ��o��h��9�������/;Ț�ʍ���\5���Mu���zF�yIm@���/����u�]ʽ��ٽ�����=�	�G$����,����%
y�4V�C� �)��6tS9إ��1ceuA:)�u�{�/�n�P���
{��ö�d�U�� `��9��r���c"˞ݱ���)�UnU����F	�����	�Y���f�R��x�_�h�dod��,%nֺLW���M�gD�p|ć�π��Ǭ�k����}_�w*��K���j��^ʧ����~+:d]^?��k{���K_�g��_�������|~V���Çs}�{�ƿ�����Nk�V;��x���:h[��N���n�ٯA���`���Ʃ�����a'�Kv����,l����q!���`��#Z ��_����Ix#��.ކ=�mБ���>S2v����k�B|AyO�> :wқ�@��$�2����ρ\<���m��U��]V�'�ՙa�Q4V!��E���;dŐ߸D�)A������E�@��R�Ro��Ժ�_]���w��]Ag'f�
gU��.k?���3yP	4�K��xAmm��5(قT�_4��O|�{���a�^�mw%��������q�J�ڵY��
�� ����ٿu6Vr��S�9�n�8�]�)u��ˇԺi�(݌6���Y������c0��j��Ʊ٘ݚlu#:m�їD��y�9W��_`�ur������M �)��-�E��5�������w�4'�3
�K4�sv�����瑍[��3��8TF���1��Zx�6Qu{F��H�&M��mIQ��̆w�q8}�lb訊Z�0�(�LGr���JĶ��i������N���9�Q?���:�����8aJu�?�S?��3?�y��_���~�V�O~����m߼������}��䕯�i��l�����rX��l�}�\�۾�dC2r]T�2�4N����[�vȓȜ�Q=�r$�*-����5���{gUW��٣���HT�H��pk �N�I��8�m�9����8gr$��t�%��|v,*Y���c#'\�#��Q�U�N G.�b
*ʿ�؝6i-�\�%E�1��۔ ���	��v19���P�J�oLRsX�v>2$:�B�k!�Q\L,_u:<[�Da�'J����	 �ng`�r��,��X�yv6y�o���_����������ң�_�����~s�*Eԓ���f�Ʉ�b&mm�A F_���NdE����ҧ^��{tq�{08ɝ=vh=m8S�~t���ޜ�mkd�y���[�����x�<�
A�A��B�%�;f��r��(~�6�,@�EvM1�b�P7�8���H2k0��(t@_] ��5B��f��=����F�Y�cH)���Y�^g�1��N��⌠�O�z�C�F
���⚫D�%g��<�{A9X޷D�]ktB�b�1�'k��� �����=�6�����P宴��%�\�3����@3���ۿ�o�������/���>{�E�����
<_��
|k<(�������G�2"�/�*V��*S�6Ls�X?'#G�,F���E�zC�v�Te>�|�C&MR���5�Қ2�"�ׄxF'����:�l��Wxg'Nְ�f�Go���u v�n�V�n%�c�CZb8�>�Ug�X���A\�M%���R5�7�����*�܌�B;�(Y2���\HP*�k,%��f#U9T�R")�R����	t�H,�J���$5ۓ�8B�	�5���%Wl�m�c׾�>�qy.���@h?Z�d�i#Ӕʠ���TN��\����v1�yM��L������[�4	>�-��;�w>�u���L�x ��̙aE��s}�	f���ݮ����T�0{�$���i�h	�^e��3�
(	�QL�4�Ԁ�wQ�ϙ���L��b8-�����\<�����7�H��ן-��P8L6̫7i����ݻǄjG�������!�Y���y7H)lnþcEgP98C�[�=�x��lŰ�c&�]Q��Jv�v	^mٺQ�; {�$�v�cP�Ǽ���(�3�ycdwZK*��@G^ԡ�Uɼ�D���������&���鴩�9��ٚ-}!6��b��k4�������/���?<�ʛ����r����;/7._l������
<_����7/V{�?�����������*?�����:_��q�l�5;_�Nk�A��t�����vֶm� ���R��>5i�dp��^7��ո�;���IP�N~lb�����joMlm�wA��uB����QwD2�b2upVj%s�D���;�d�n;����F0���^��m
��<u���eT88g'4�l�{�;�F�8Yj�N�P�� �=���"��r��I�Ҷ��1�L0�c��>�R�ps=�{��Y�%t���d%��M�w��Ζיg�;��	�u
�W[Ió�r����<�\l�{�q�Io�Oܡ?��5��j�!��8s6���2��k��C�E�\VeA�8��}��˶QՀan�p����<���!����:+��@����$ H��qIU����l�`�@iI���#3Zޱ.����N�{'��sj���u����2w���v;�3���D�D^쵏I@8Gg9I�0�^Y�!���w�Ҳ����v�������� %nY7�yƕ��!���{x)�G-�^��7Ȇ��N�� :��n�����&��S,P�z�C�ɺ;\�|���M��i�JS��;w^�/7�����O���Ͽ�������_��O�؝�;7�._n����ҧ���b+����������9�����x�l���xQ{�X��J�ڹ6���e{L�:��O��S�-5��2�ᾷ�Hb�0��@��C愎Q�9�1����1��ἰq�?9x���~A�I�A�Bf���Zwf��0��2NW�'�򛰻��	p�j�P�4j���Z�1�<�fLb4;ِ��<w��ԭ�����$V�h:S3|�s7K�����R�Z]�D_[wmC�<*b`����.\4׬�u������~@��hԅIM��۱�N��9�zp˲����Y��:���c��|Q�V���'~���<z�7�~�ϽB���������`ގ�zŅ-��3G9H2�nB�Y�mg���q;�e��0q�'�"Zjr��̝�b����fpˣȴ�*:��� �pw�:D�􀶅�����4R$��	oPpS�@)�_��~ ﵁�_xAV*CMW��$PR��yX	S�FM��D�%<o�}d~q3�rf�I�ӌ�^8��/�L�]-G�E�,�	��$~o"y?���0̕�t���*kY��\'�EX�[���45�9#�o�h�Y���S���6Dl�l��:���.��>��,Ē&�/�d�7n��n+�z�_|��?z��������|��տ�O�y���{o\����y��g��[�Z�\\�޼�����k����ϝ^�؟�_]��^/6������t��^܇ς���Z�sQCK�@^��[�2��a3j�u�������#Jy��q����.8��v��]/��p<�ᑰ�����!�ݬMv~G�$C�5�`2#�ѭ$��'���9��$gM��j[�����f�p�]/��$f6 �yJ��Z�y�����ܛj�Nu��<�^5�2ɩ����;���2���	BL◎Ԇ�f９���t���0(P��3y��ZX탢Z�̃R�S.R�w��dd}�e��gJVv���5�8�Mt���{,�������5�Ce�_�|у��	�C���Q���_�e���h�B94Elu��,��e�����ր���]q��ȩEl`_؆��#/�n�D�l����rZosi�cO���˨���.�1%:8s�ۯ���RGi$�F��U�C%���(;|��X5�\��k�I����=�Q��]�R�aY����I�3(P�`�@�LR��F��F���h18	�����n�L$AR�mn����P�D�^[]`$#ay�Frԩ}M�ul��8Pf�2KKS٠"_��ǵ�s�Y���������ٜ�JI���kO�0{��z[�ME��5�n�����ԇ����o���A���^�Q��?�Ç�޾�?�oU�w:�O���Ⱦ?�?+��p�AXe��O��7���w.?�^�^,o~j[8zy�hv��|q|�#�̩�8�F9�AX<���'�ehך�c�`~�Ɋa���l6R����o�CemYp���9&Y�d^�94).U�����,N#����%��q趐92��|�s��j�iEb��q�s�d��@�W�0�Vn�t����\>����#I�3��&lzg�]�TS�1��"[~)PRp\�Bc"�ی����1®��ێ洶��G߸	�o�P�K`v�s�G	��`}�^�H�Μ��OU�$ٗ�&�&����xm����(��(+��������o�~қ6���+����,pt���!����*lFn�hFO`��']c����1GFĹU=ȞM��k�����s���pn���7F��_hF�X% �~H���~�+��T�@(\/��tp�m]kǤ*ʂ��r�-67������9N�`�C���8���Sܬ��Bx�(g��׶mP�ip�u�ʺ���h������(W��Z�:+>~�yID!����5��cde�/!�My��	���2a]��y�[�4��������=�5����[���ku�g���Y�&с�� �pzL f�Z�޸Ѭ7��K�[�)̆?��<�O���[wۍ�{��s����O�{����_��������+�#��-���h�}��G�'ӣ��o}��Ͼ�����|aU;z��`8+զ�:�	<�9���X��Kϭ�iY6������+�c����~�48�)�!�'<�e�;ĉn�*N��㶭����ծc�TS�H�c$��8�)�M�+�.4ܵ�����s�����3��,��}������t���)�m'�aO*ι��X�O*`��A0�1�9��5bo�6�p(���r�$�����f�M�;ۓC>;f�����B�Q�z��%�D H������Juvk+�%j*�f-��̶�nF��s��?#�` N�����}x�x���'�}?����p�x�֚r��#�4 ��t����7d�B�Wsn�uEb��9dbҪenZ��L'z���ח(�=hzJD�x�`�u��#�	
��a7�����ÆW�X1F��(?���=��d�S�Wg^���-0�&��x��S��K�����B�������p�V0P��}Ȫ�����3a��$�o�W9xB���W���_E&�!���r�b"j���ڧ6�U��p�.e���Y���T �������<H�M�΀��N'�����8����(1{H�:�ib_+=��^�ZL{hOBD�2�Z��B<��ȡM;蔛��[���|1��t=�������G���{/����������7���Ƙ������示O�:<�?r��oZ����|����|�7Z~ꃻ?�ش^�o�/���*����\^����8&c%��n�g�j����D7��A�:f?L"(������Y	{�n:�p�kB�LN�]֝k�l�n5*�dM:R����&$#�Tz4��3��7�z9�©i�d�_���ɉ�&x�mtʺ`���zV�)eNɵa�!확���P���d����ߕ����->{"o���J���# p���̞#�A�����Ej��x#�2�f�=�1�t��x��֦�j!�9��>$^c�&R�S�];(�av�zh���a^����lh�f��������y��>�c�:��xY#�9���t������[2`�D4����3mu\FNk6mL�A]!:*�E6Ɉ�U���و�\�è_/��L�!���E)���;�}]�u6��:�1�-b#p��v��'�8X����d��d���z�D�`/ߺ�fr'w��q�{��P�"��Ysx�8��rH�PQ�CDC
q�i��8E���HD�!* �/x�ka���L��x�;9*�9"[i��g�y����³�Bs1�h��F�v�Nݨ[ �4�ZFq��:��?���@��Ԁ�8�!��Y������6F����TlO�R{/c�5Yx�k��������~p���o����Rav����Ν[����p���k�>�یA;����'yX����xk�m����y�~����_�o������/��OZ����|��G�i�=^+��q��RGZ��<%Q���,5#�kR�s�Wǥ������S�c���y7��~����8[^�cp3f	OiR�ٯG<�x�c�G
� �K����[���8IS���ĜG�ߵ�!��]%fɒ��־u������^�<#�'�.Q�S[�S�s$_�q�Km�$3�/��#�4� @濙S^pj[潽�i���rpy��]O���b��l�o�6Fj�c��ԡf>�EMt2�]9�.� �j�v��8�-&{��]O�@�m �2�f�L�A��)l�"(�$������jk0�|�k'��Ե�'6N�v�x�R���l�����}@*SV�l}6����1sz���n��@Ą�qH=���d�:<��*� ł��X8��}���t��~��kL�~��lty/�G8�Ly�j��(�fC��	Zo�N��`���ʺ��95�e�o��UZ5ZP��L8�����q��^���ڤ�#�?�?�Hw+4�ód`;Ċ���U&©W9�E`�6T1�5�9�ɩK�򎣎���z�#���'dݜ/����y�(DY���S�\[f��:8���{�xa�K��U�<1�0�58T�2��8K�����A�;Dcr}�[N��P�۰�2wϙ�:�~�:8�JZ�:W-Е_�s�w��}���b9�����G�N���G��ѣjy~��.���{_������u��Z�V�0�]er���+����p����~�W{x�k��h��_�w_��dZ��lS�3^�_ؔ�w���e'�\L��+:o���+ ���l�þO�]�|fY]qav鸪Tr ��i��Lpb)��\�B(vv�B )V���x�9ޓ�j���u�D.��nK.͂�d��t��_h��s���	'ƌv�-*@�+��Z�[a�E�����m	�m�4�<+���$����4(��4�ېh;M̐�V����$ap�����ȸ��{|+-+X�H�1% ��Nn�/�ڊ���\s��M^6�" �b{�0�I(t�2�ݡ����b0 �Y�˘&BIH&i�[~LS斔F�38c�N&�V��Dk��P��D�U��l]��xdQ8�G?��Oԡ_�g�u����ʆI`n�r��Ԉ�pA*�.ㄱ2��3��vT�Ϊ̆���{����M,Cf2�Z�a�}��**��j�����%�����uȢ�D�F�1I��T�#�|'�EU:�j�_3��Ћ1���C�"�-tj	�����\��#�Q_�v�P��u�rg��N�>H�A8�1�NEc./�M����Ҍ|(��8��s���Q���^�(��%Q�R��k1{wZ�T:��T�h:�5c͋��W*OE�jznյcge���a�d�z(}����8������$�ݝU#�j�����]����X&���>�]�p���j�d���eS���bes�}�4e��j9��O/������=a<�o���_��?���;�/o�O���ku.�����7\��/�G���ǽ�������[���@_)U�Ǜ�ዥ�u�X�G�M�u�4�������â6K3C���J�M����w�8���B�YPmiʹ
C��LY"�"����6��ʨ��^��<�J9?������L�!q������Tb�����j���+P�p�2��"e���f�sΡD�|�rX��9������@B�Κ��8s�jk��d�kb��oy�2Ɇurgo�!�m%c\>���w�PNU�Z<θF����1��C����`?��kg�$T}`�䪃�K�U�$�'��VK'�u�SH�~O͜�:apQar?�5�l��5s[���/	t�Y+��FYe8��%�C�{�Ĭ��kW/a������7��y�c�/4��ʵ^��'���:��dv���K_����ܡ�D�	�JH%����@�j���o@�.�0r�゛2�ǛЪ��.K���t��Q�h��;?~�O7t����I� ��	�M�c����J����$k�����6Ï!��:#JL��S�a�C4
Z\������_������A���򈵄�q8�D]�8D:��ᜱ�j8�&B"��cC+��0BF!*�rR��;�y�vzP���T�3���C3>s�ֳ$~�NҊ�i(``� ���	�>���Eyd�a��<�'^���̾ⵃ.����5(#}Y�~�%p�$�9e�	�,�+(�Biު����®�6n��hL�F����{8<}�������'�F�޵��7����{�o��۵�SJ������O�=�O~޼\�G�u��w��٠�������];�>Ky���r'W:�]�5�WvƓec1-6��me0�qk��k��{uӻ��j�B��nC�U���.�;d�����^d�"~��/�\B��$����Ѵ�U���]��$��:9g����ψ�7�qc䃓ҔZ�����	����;����/�(iK���z�`�狞! ��`��tL������623�8��d�t[NІdkm?9׭���钭�،��=��꜒$�y����e��9 7��@Ni}s����23���y�� �	�KX�����9x���t�$2�B7aE���#}w�
�GKax�T�}��9�&��E3�:�����q���s��e�xl�ʅ6�����'�������wp�mk:X���J@��t�:��9��� ���b���M�ү�kUT��K�*EX�S	�-?So�֭#n���=n���q΃!B�Zz��\7p0�P���Yx��@T��uu |Ej)-�]T!��+��2�%����9��\J��yۈ�����rՃV�����Ú�pD�#�j}j�f3ʺUōF��V��,T��e�R�)� ��v8#�T�b�plR�/�T*����K���s����֡�MZ� ����9����~��E����q=�pW�0�ޘ�K�IP[��l���գ��V����d��!���@PV�����1��H���@�J�ެT[�r��!\�W ��8,��G�g?�{z���Y�>�~�����ݷ��߾����5�qT��~f���'fq���wN���d�x�_������у��g�����b� y��M���:ߺ���k�t�J+��qi��S�dR&BgP,�@�&��G��XQ�E��¶8������:qKh8r�fagϗwÛ�1��q���e�7а�N���k��|O����E�]A)���:t�)�Z蜫��u��sc@�����D���!�����7D8k��$XR�]n��{�&���wL�V�̉�[��7��T�wTt]�ާ�cHH��~��
l�Ȟ��9� ����V���Q��^Q ���нYBNËF[�ķ��x�eT9W�v/��X���TX!���%x������S�3lQ�զYz5�ѡ�Rt�e� �� �9�S�{�����b����u�A���R�6DT�q��*Xt
��C���,}�� ��u��2:4jmRk��Lp�8G�R�U���ad�.��6�?��nX�p���ED�sZ�.9l�G�-Y����?��5��;���;�3�ɩf�H�Ss���6<�6І��0|e��d���d��vېa��e��rk���EJ�T,V��U�Yy��#���g�oD��*�V����ɝ���{��{�5<�Yk-8�ۦ�T\�\Kl� Ȗ`�[7�d<Z3 ��, ��JG���eȯ"��`ųXֹ����w��`�?����������2�ĝ� b$���L��3nn��d᜸�dƆ�5��S4���<�лՌ�lĠ��}���oMZs<�7���q*�L5�nܽ�m�j]}�O��U[B�{y��[�ldm$�g�!B��k����.�l0�2��\C*�Aбx�̚�ܗ�)DA�>�Z���������� B� �࠮��_��;��W_e�RI���������q�j�;�bJ_�m���1�ÿ���O�{�w�h{x�xg}���������o?�3�Ͽ{����b��`:~��b�������7�p~������������å���Y��}pM�0�����pv1_>��zr������M��.`@�*m��1��Zꖳ��ၡ}�޵~�d�Os���7��č�1��%c�)E��u��-�N&���U��)b�V!�x�R�����^K�H�ɤ\Y
�P��x��^4.�OJ�G��:�y�`즚9V�L�l�^~v�bT:C�59P��x��<�ɦ��,�*Ss�,)�G��� ;(�G��c�\������������!��נ���+��x�7)�W).�Wn�9����M26�~��0�p��>m+ A��T4Q	�o�(�;�##�XYj�V}B�A�^�
׳��u�ѶL(X2�o�5�������y�VdE�?��)k� ���f�C$��P� VXrݠ����+}�1~��ع��oZ�uˍ��!���Se3� �M��U��L��&���o�SM��;�b�H1�{\�yj�{�*uב�\�m��H��ڴ|�@���w�m�4�æ ���<$���(�FcY��1����O��h������?jp���Q�u�����/;��o?�+������jވk��*J�=T��_��wa�]a��i�kQG��yG|�#�0)q�<����X�J�J��4�|z�n�eb�*���]��5<���)��Z^��?Wc�Z�I�a�vP�H�)B����"脄#]H�2�	r�o�R���|��C9��p������������{��������`z��������G/7V��Q1�C����ڷ?��_z�����O������?��x���M?�̿0��_���������^M7O�������=�\�G\�����[��[��V>�m�]��6)ѩ_��,�^�+a��3�2�C���&����e�d����1{I'VA�l��F%���ƐOO�>��5~��65-U#���&�M1Pgژ�lŬ�/��gC�J	h�^��e�u@0�h`$�X�{�2�Q��^vkS�Ȩ��;�B�/��8�g*\K�aJ��\��4�z�)7��ظ�O'`�C�F�Y~��e��ѧ�ŭ��ca����}��8h#<t@��w=�-ꣽ�Ԡ_��`�in��ΐ�'��%�s/a�����M9�b�#�ډ	� ��O$��Jq6��e�s-��T6Rv@3*���BfSm�44�uN�u�$2s�T����-r�W�Q��_btXg���$eE�n�"����v���C���2o���:7m���[���Ғz(=�Ļ,���AaF��(��Sm�عV�fTHWxq�b^ �k]�����oC���;�����?x���%Է����q�Qn���w<��R�Ӝ�,�v���Lw�]�{�#�����l[X�("��S�.�9���xu��MbD�ո�q��O�`Ll�����pH�:�!!�����< s�d�/o@��E6��.�1��e�vE){5����1ř�!,�e���Px���<6�A�<�;�����d偫Й76C�C���̵8�A/�!�6�2��
�+sN�=׊`�D)��k�W�>�A���Yvœ�c+]�9Ġ�ZT�Ϗ/懃�-wk�A����x�ؠ9�dI�5��=zi~:��P��p~}���_}p�j��� ,�|�`��g�k����8���tsc���̀ݦ[�K���r��������͐x��������w�<<�\�m�o��������,�>�]��P��)�rf��x���5��5��=��ɦ�Z$�֟�)�m}t��.��66���UV�s��yS��}'Fx��z)�,R�b��i�R��*� (�K�vc2GR�2��)�5���x�!�XO�⹷{}��+%^m@���r!�.F�(���2A���܌3�KΑ���yS�O���W�b�i�2��:�9�<c��g���Ƨ7�1"%���}z�,,��ù������(z���1�'�O���_�qs�%�O@1��弌�B[��;�\���42����ɡ�i���|vŐ)��GiI�~��lJ�2&,bN;��6�2�Єf��ETX�B�C��/S�l�}JMzm�!���(~o'�K>��^;^.�����6Ƀ��lu8z#��S诎�P�����ުMA�eS\����ƣ/�%5G�e�B԰�p{j��X���s���ɦ*)���3��l��jK��X0�����e�:�'�(�� �ailcQ'W�����Y��Ŗv�q�[26��bem��_���2ga���ل�ٲ�1�MO�S<�U,ĝ�}�gڳ�N�H�;8��xC���4����<_b{*�U<y ��k;�IA���ՙ| ������Y�t�Ka��6�ܽ�R�ث��B �?�uI/^@Y�	���@x9���h��� ä�!D�{n�+c��S���Ž1�1�Xx��ד��b�̦d ������x6�Dۦ�8&�3��xZS��^�W1%~i����W�^LRN����"��L�lcg�4}���7�����������{�WG\��\�]��A��z0�������of'�ӿ�/_>�>~�>y�p{�Iy.�i��O��v�}���������z��[;���=;9_&�hx|6ѽo������.nޥ�c���l�!p���xoc����ߙs��(�5��[huz�X�����+�:q�%㺦,�K�n�;*70���(���af�ng�VJ��67����xzdvJ��ܺ�*Ӝ���Pf	��BkeJ�mK���i�h����~�_!CQ?E����j�ʗ�u�-Q���K��OT�zᢈ�*�l�'�OA+�G��Ҳ�3�Ya�FxK�L㺌�B��4١�p�����`ѥ����Ĳ�`�->���6)h�(5!	ne�B����~3�Nph�M1��~�s��'�-�N.��Ls�SsMPE�YR��{u���j咞���,�����!��g[���i��8F֛�v�-��%CS��j�K���5�\���$锍���������G�Z�i<�E4�����p�����ۗ�g�^�o]P�u��:K�= �S�����\�F�M�
yD/��L&<�Py��Z��ǴbM?��H�̀z6�5U�F����~Jԥ�'�?��G0�A���f9=<faP!�H�s;;Jݘ�����64��75�D(,qu�U=�ĺ�[�x�OP�ԇ��s��C&h�?�ucuVJ�ZۧZ�Z��)D8[&�� ��d#	��@��pƸ�"��͈�K���~�9�c����e�My��m�ֲŇd�����)8��x���b��I~7Ֆ08�ϥ��ƘYF��}� �bT�	6w�}A��wB�K���3Ka�L$�|������DcfcDkE��� ��8����3�(���ߣr��4���,1{+����Bqc�����!�k�������9ߴ����p���px~��zNj�5?���?�?~�{�@x���NŻ�9D�+������"��b<Z������Rx�_G!��ܬ�dV�^����|8u#z���r��t>:=�ܤ�ɣ�����?7[��E!���Ž�cM�J������>Ya۔��"f�~��:�\]Z�/�������j><c��O_�QG�G��a�����6���!T��B߼o�h�h���=�_���
�4-9.���fK�UXj�[���oq��!�G���8��M����s/,ڽ��2���9��`r6����։����Hf_%&n��}�~V�p��*^Ε43���2̢�:�A���@�/���r��������BBso��o�P*�YA�g�̔;���� ��Δ6QZg�=�����3���#�����D���7l�V"����[j��z����-�큑��2��)�C&�İ�����2NI3$��5��jM�a�d��aP�G+֐O)��c�t��x�������ZU�$f�| }���~�Q��)UL���Ͻ+��G�Kd���d���+rۈ�	���x���p����??�z����3<8�P��r�1E��X<;�NR:Fa/��v1��M封�eC7HZ���u l�Ā��V���T�.F�V(]�M <xL$��)id�=�G�A ���O$%�����i	ס�z�1�-�X4�YHZ~Vbڟ�w�ۉ D(S��aW��t�X�#v�*͈si�. ��I�ᇻc,�G���u����KZ�DA����kkBa3!��~��%����4|�u+���N�d��)z�Y�U�����g��O�C�i��w�\�Ƀ�������&�6?���-�}|v(�N���c+��d��G�v�E*4j%+�'s	B!�l~��B�PR�$�����ׅ3e��g2�9��p�)B
"�(:�H��2�zD!Ǆ�aBU*���눋��K�K��n�5:魬�]��0s�UD�NW������tvv�rv>���./���/g�7������?�.�=]����o��̧ 'ӽ��tgmH��ќ����5�S�D���ͅ�ע	���e���AZ����'m{�V�8���$h�"�Z�7�S�CTT*7�����DK�@�����׺D�c���k���x�X��t����������
����ԣ�����je����%?�W���l,��o��w7؏�(�0!�liCnB�2P�
�aYO{>?H�l�M���8s�����%�j�	s�"Y�~��E%��=���]�[#O�w���%�:�=3F�0<��T��U�rrOk���q�P��2�&�&Ȗ�4��W�}}�yw�U�%�5J+Qv�g�+��N<�=U��3'�~���[�Y�!���A�iY	�\wI�t������O(B^[�c�,�U_q=��	������^�܋�b\�+���J� v��1v��l���`iÌ�Pn�����A|{#��ؾ좞1��;�k�Zp\[P�sPG
�\�����a݊&T��!�;t��`Ϫ|�H��ܢ3k�ܨlI���L�x��k�"4*��cJ��zz#E�~0�9f�)�4 X�yE��9X�_/����S�y���ͅ���w�V>o�_�k>�d��7��7��N�4�c��	L����V
��[��u����p�xX��o72�#R���\���փ���oa��e��G�
���� k��7�O�7ʗ��������Rx�B���*P�^*sS�)xZ	Su�ZV��va蝦���(��X�c>#l��F8���Y�T�;o�]�뽂�!d}�V�ƿ� dbPXLBxI8��F��Kc��M��
Z��٦L�%'��D�`}nh/�Ђ�	��֛��O\mM�o�N"�d���XȺO1��b��e�1QJ�B09�J߃F(�N%l���^pC#�Y�N��twR�ˎ5]ζ��|�:�	�/C����8�*�� +�C22���fgѢ����\��%(��@#Q����Һ�WvSQ�6��+x���愣7�[�2�����6e�Q5_^����pm>馋�>?�>&��7w�R�3G�[�����V�ƹ�%$���  �_���m��˰沢k���eb��/F_[
k��G҂�O�SWkCH!��Q������1)`c�F�
{hyA�0��	o~��İ<'Ģ�����i������G7��}ԁM���F�:1�(�Oz�����?e�!��4
CrS��.cǧ��}G���R�ZH9L���JAgA�ā�-��m���d���X���M�*n2��"��o{I,��+�ALcj����-Đi�R.Q\Α7����6O�ZYiq�u#��@"%׺�ۇ�6��ˊ�9���sѳ�C����`���F(ݴc�f�w�����.e[�����x���ޟsV�ma'Ȥ3ba/O��Q�Ǣ������	H�mdPf2�k�y��å��vJ�������|���dD;D�`�`�p[�4�c�Cnӎa-��O�DJ�j��99���7X��8Q�*�{_��g��`�=1���hH9�8w��g{�������(�W��;<9~�J۹bt�؂�����N*	EG����"���튖�&�>�D�����5��Ǝ<:߷���Z�I��(yW�Xm�,��}:�]=�b#��WV�)c�S�����Nn��ʅ]����e�K���,\Wg�E������ܧj�3��B5�����X
7�����_o[���T�ۀ�f��S���6��0_�N��5x�^����E)��T��U$�1]��N�-�V��a��E9z/�\D��	��G�O%<�[��7<a��VBR+�k����?S�1�W�_V�-]�#T�k ��XpcyD����c@p�6�K�j��Jݴ�6U��j�������y-�s����|��d��5�q�g�X��u����!k�q98=<bJ�r(���%ǳL����/��Q��D����b��X�
�gh����TZߠ1�=�T8��d�.0�^ޏB�(�<"L��� Ze	bY�ZݪB�K��
i�]B�³z�K�'[�Nx��e�K!�[���z��͖۬�,�� 7Q��P��W)����~�u_��uX��A��t�0�Ʒ��וu�m;����p�M���x�ޜ�Z��+ʍ�����	���θ*>�6m;��qgٵV������f����G4�t=<k@��ظ
�
6�$�j��+[ �*�!s�'ה�%΃��ԍ��T�x�Y%��u^d�3ޥT���|�f���+����6�L#�1�i�½��B�y�T�����,wQ�[��MR�v��-��=�.�%�N=�s�n6~9�^��� ^��ٰZ{,9�#�g��"۴WQ4����Ey$+�����z�75�hINoz�d]#��B>B����Y��:	N4ûT�hD��#�D�s�׽�~��9)Ҧ)�,�Mڟ�ը��p�����������F�w�w�1Y,ol\ҥk�T��Y��t���hȑ��/U�� ;�&R��,�b��X��9i�*Rd8�ٛW���mr� rњ���yE��m��'{X�׃�}p�CIw����z�W{�o�*�%�]��n��v���(0:$���%d�"�ri��p��-��r?ϒVƁ���͘'.>[�x�R�`��=	V���F�ɾz�*�ix6���Ǒ[J���'���/��RJwi�X�l��I��=�RPv��<V��^ĭw�X�^���#p+�-1M��l��^"�:���4�lU��Ԕ[a��k�Zg�
�����`)��[!�����`�ސsp3i��r|�J��=J1_��`���K�� R�b�
 ���t�����ޢ�����:>%$�S�#�����
��Wp�G�:K����|m�Ό~w:5tTɺ��^D{ԗK�9�
�0���N_����,ק&����{��W9r�Db@;'� �(�L��~��2c'�A�M�3���Ճ�׌�jC�)hN��T��DṦ%�����Ra�7U����ɦM�J���\����YK��r�����}��s�7^빌Tф���{hii�֚u7Q�)�Ա2��;@T�f�U���_P�[�z��'	��;�(2��]��Ƅ�Ҝ�)%d��&
�<�1O"��ɚ�5.2���`E�MȾ�T��lZS�"���˚�k��v���.�����֩��7���I���a��)"1e=+o�`���
�Q�x�wz��r˜ǉXhW�5�g-����	����F���+g�V��}���{�_���Z{�X�^"�%i��	k	�}����U���s���$�β���r]���kZ5��P�D.���Oi�M~���G��/�O�Ë�_xw�S�ȼ�����)��hyx��4���e#1�B"S6�=q7�m�aZ���p*��0�ƟO��˪����N_%��9���;ػ2�B
I�z��[К��jG+T/#�bO��=�x����Ʃ�O^b��R����wv���d��������ض��M^\!��+���o�t	M@[�
*U��	����l|c�2.͋cE����i
sL��/^e,��16̛j����skF��Z�%O�7o�=�}1@�Ʀ�`�kH���b��7�e,QCDe�F//��k��@�w��+E-ݸ�M��^U|�GЖ��<�0�K0��-(q_ѫ�3� !� t� ��En����҅o�D8��S���ǯ^5]MĽ�����
]�tkʌ(��3�������ى��<���@�%���5�hyT������p�����(��͑�ތ����Wj��Qlg��>R�����z%,ާ�i�A5�J�T�M	,�"
^�T#CI/�ˏf���HN�w�zb�(古0����V`���ڸ ������C�"��g";J2$]�0i�K(�\���Hit�-J���0#��05���2bT�A�\�ͨ���Z+�ݶB�nT�S����S\���}�'wf9��flQH����:��s�u�|�$� ����̀t.Q�)���c����
J��*�"c��
�_X����`�Ɂ#,O����]I��8Z�rՄ��<��!�Oz�9���j�ȣW4GQ���꾡*�h)O��Dw^2�̵��͇�(�ה��,bk�= ��5�6[$�Z����m[mY\�FZiԆ^��7�k�M��G���y֐�V�3%��s��:=::I�Mxf-�[��/�^�$O���ɘ~����??����r���|��O]����������>���!���pB������ޥl�*B@���G$��7�en�L%�I�C��d���%�mLΣ�u���Q��ػ�__�0׷���&�����g/Q�"�(f���u���T<:Z���w��*��)��XT�	�\�E��H[���
�Z.����^�J�?����p�i^�⧒1ش����������/�����T�b�H�	���r�Y?���0����7;��}vO=����TQ��(ίʈK�8S�(D��O���8��b��]�y�(�����Z��LA�&��]h��B����甼ihA�]��^ao"�O��(�L���>swE�\E��w���3P~+���Ƽ_��
]�2�Q�*�;E�B:�u
J)��c�0rOD?�Lǝ�P3���OE{�P���s��ϻ��~�XS�7C�?,�,��֧��_ҕ2�{kh'$�Ƒ� iA!b?=��_�"hb��Y.����z"��}W�Amf�C�;�W���k�\���P���n��fϞ׹��Y�Z��%�2�jݦ�J�o��)���k ���ςj��z��{um�5�#g)j<�^$�����{ĸ��?A�a���*��3�PT`�������f;�h�'�O��f�A�:�Y��N��0N���v��Tm�|�!��l\'�����M?ka�t/9����zn=d�	���Sd�)_�SU:(3FVړ��g��D��-��P�?g���M�D��gN:�����@�����AQ��)ǺGїMK�j�0��a�rōykh[q�w��;Q�h�e�U�1l���Q��Κ�Ξ���GŹ�=!�0�m�:Z{������+����W觧W���巯�W7 �dA���s��u'����u��	�SӋu�}�5�Q�ae�,U�C� ���$,wf4�h���eX�)�/��Ӎ��M�M�>ٸs�
]��TqSA}��s,Lkǯ��s�������,0�*�iX��y[��%� ����:��D�w!�)1&�y�
�X�%�\4i萔0�0\��hDnd��a�X�J�*��Ǉ��%��TI��DN��A6az.���[@���ӑ�/
�s
�t/4e[��UJ����J�4ޚ0���P�"�9Ԗ��<�\�=/�5��5�X��&���u��~ճ��i��lz+�鱄��F��<\��lt�Z�L��Z��j)����%X%�)}^o4(��ګ�^g����UP*��3�amＤ��1d�ә���eV7�)0�'��wqQ���9�יWY{�?4
�s6�o�2VFA��]?�pR
a	¤Bgl����U.��I'�W֊��*m֮u�*!����ó�{�}�?�����[<���S}�}vN�0i%��}���qE��g�Qezjޑ�Ռ(�ANQ�5o�[�wJ�y0�I�F��PΝAU���S�.�����i�tr%�m�	l�0���=���'�>7�!:�;�^��Q������_�o�<��X[J����1�}��Cd��6\��崁��z86��!���Y�>�X��a|G��	/1O�9RN ��g/����$gan━(㫗�!�#��X�\ �i:����*VI|�]AI���>�!3aI��^�^X��.x�{f�4Be�קs�р8!�IenuPE���ה,�o;�M0Hg6l*�d�O��kY�M��f��t�s����i��{�T}�&Z��L�T��
��&�[Nr�Q���؃�V���]}�RR�γ~��H���M�I�V �"�hO,g��w�K��L�9���D�6��G�?�M-�3�OغU�ŎdG`+#r]��Q��$��w��7��sLM�����(��0�e��Ucj��/��%�g�>��-d�7/�K���.�؆!4`!��$t�Qn��cA�Ӑ��HU(�o��0�
�I(�7牃�T`Jt&�� a�����-�*4�F�Ý�V𫋺*�i�)���zx"�#�y���_
�+���&���z����4Ӌj𾞴y��E(��\�xt�b��6n�/$$�p6�Օ��%����6#L���+%��@kF#�1��WP4�%ׯ�ټ�D���s֗K�ʋ,3.�_���niQɉnJ/S���I-����7���|�De8C���vg��[S*T}�̅�iŃ�ך�M�=^�U⛹���3,7&2�q��e��� ����o���2=�����w��e�٘�W����L��-͋�q��=qj���^�8��4�"uJҔy)|M�Z#�=��2>ly:��-�w�֌T�֍_B04�J�3�JK���vL\�ŷ4��z�q6�5�pD�8��˦�R�6޸𳗓PPP$Cb���"� �����E���l��y�s���
7�!����G�@@<�>�98j���|� �C���|	ex.墳ϔw�z��,*���d�n�{���ڡ��>���W�I�mƺ�m�����A���=e\/��O�x�F\���H��}��Rz2�	ň��:�~ެ
+M�L.�����z�j�N[h���"�%� -��g]�9T�����L׵O]�g�$����Ҙ"MZ�Ƽ��h�L���e%��oP�6��&J֮8v@�k5E�Xz`=�l7k9�4�͘I�D�1�@^%���	+]�lJ�1W����@	^/vY�}�-��^�B�*Tn�k�Bm�*��h��NBܰ�W퍬�i�%,S���,�<�+gmѮ�tfW�'vv+�J����j	
ŧ�s%�Q��M�l�9�&�]��������8�α�Eq�1�zc6�M`�����Z0�K�1"ci�8�0�����U��M&x�Z-gӊ�����9ZPv1�&C	����s�Q2�����A��"����gne��:
C=�sy=�nJ#��:7iy�uN[�[C$��R�)�ȿ<z����	������
��~�D �\d���(���}����:�y�o��w}��=�-�W4X����Ԑ��46����e������M^ZL��4<�kZ���7���519�銶<�Tsu�o��,%��l��k{���̅L^!F�ԉ��nBtӋ�bd�K�!�)��
]��y+��L�����5�<-�(w�C;$���7�c�tʜ�­s)�e��.���B}�B�m�w�ǈ��o�8�M�[�m��l��ӌ��=C�����}1M��:"����%T}����X��2-{J�Pã9�Q9z+��:��1�-~��1̶
�AF?c���eW�6�2N��K\�`��Q��ѯ�o��$�Z�uUe����D
F�Έ��)��b3"��ڹ)�T�
X"��Ù֠���`{�����d��ݫO V�{���Rw��K�ֵ��&j�q����r�"T����S�Xu�~��E�\ofNS�{D��5����i�
B\e^Ό����l�5�ݙ�P��<>u�N��գv��nV`ZiG����2�/6�K�wd�`%r��Ϗ>b!P%�8�������!���F���8�J
�مR������$L����׿��ZAH�����qv�0�>f,�Y?��YN���j5e�z��kޢ������a�E���8=���_\c�,¡!"�ǔ�_[]�ux9?���c���-1!�[������Ɓ6d��Q�s���=�;�/P�v���z�+��5v<s��AL�N��ï�U��A�j��G��w�J��1�o�bO�Q%�OE"� �0�����^���h�������^v��=��0vB��J����O�|#�#��1/7 @뿺(��twxJЉvQyW�J��^'.z9�5����QŢ�ex����_�DZ&��c��ѿ�5D�q{�W����4ٽ���BW�����/h�ut2s_��2�p�!��}�JY���Ƚ���kN�o 3�J�֣��N�ǋ�הrb�}��%F~7�����Ļ+c!$Kw�
�B����ș�p��r�F�l4���d�4��'̛���M��ae��>q�/_�+Y/œ������(�."9KkVBo����.\�G�'�A!~?ǻMZ��ɽ@�mo�F���q,R\��S�m�0XD��Gf��C�p�hr�o��:rh�z��}ݭ�7"��2���h���N)�|�,�/�K�
 c�԰�����v�6��wx�jA�t1>b�\�9{�(���1ǹ@Q�(lt�(���+��>��=�?ƙ��!щzD����̈�@Z�(�z�3ݖ�/�S?������e���s�b~DM��?E�S]4��qkPa!PxB|�±���y�=�S(�%\6�K�~\���3
����s���>�_?��� Va�oA�*dR)�N����Iȝ+Y��
gE��{�F�p�BNl*� P>��x��i�ns8�b�Ƌ�s����hr,�S��됦"�ǖz����bŘ��/=��=�p>b�{�3鹩�vq�8l���R$�f�ڍ��է�0�Ʀ�<���|ݪ�y���U�+���Ji�B*�Q$���D�,ls�ӊ���Z�ħF6=H�˜���V��\�%e/���f
H)��w2l�2�C�~�Qu#t-l�]��r����@S��{�?*D����D��=��Юݵ�Ii��G�ƣ=��{
By�\��y�*�84�+����Ӑ0��\��'��O �>��������z�x�Q��sl6���٭����Jf�t��* c��sύw�p@Ho��Bu��A6S0�E�*�<����/k$JK��X�5����A|jFɸ�ׯ���m�� 5�<��y����7���v��6#$��:ť��ź9�t�)�~�+���k_��ݮ�T"ǞK��9ȟmm�a�'٫A�l.W]��5��{~�ɢ�_;V��G�b���^�N���8Ճ�/et�$��F��PT %mͰ΀2Doz�uc�Zd�
�=�4J�Tb���Z�:��8i��V-�y�j�7����$�]��+���H�$仏%/�������?Y���,)i��B�R�P6�Y&�onF�׳ft�!a�*qv��b+
W�98&vM���v
�ļꑻ�t�����"M��%�������5��0W�����Tϼ��Lv��+Ua�7�����H%�L�O����%���6���Q��fX��R6��{(k���nm�qN�n�5�xz�����ɱ^a␐t ���,`	A:����+�S5!L_s�	�<��!�}��[TYk��%c&�S�"
�P   IDAT�!�����֍�	�J-F�䲢ٜ�}�V��h�q''&�����z�T5�q�6��������NZ�	�o̕4��E#��dvH\��R�Y�p���%�IUXaUj=�&f��k�)IiG��MF´������+�T3�\��u)l䰯%6�<Wdc��P��9�5�r��c�U�A��"GH~��P�:
m��=%!�6��x���W�%��X�nHY�Q*|�L^	u�������[��`���'����b�(�r�qW�ԁ�#�+��~o�j��z$7��/P������|WK�`���=�� ��K������,���_*�����Ѕ�G�D��9�^'Mu���I�sk\�3�k����E��?:�s���&�y�����]Z>�)�W)z_K�զ C��jB��i��N��3\k2���S�2����gx|��s��LX��nв���{��K/Z�3<sb���y�m��j���o�}	aVE�Y�Zu��î�"����x�Ep�����OsËe��溒ܒ���˝s�ʡD��%��J�j�;O�6�1|������(M�Q�^�V�0*  �y�3��"+�5�aڤE�6L�#��	n}�Z�1D�,�%L�;R\��b��w&���v����`B�1BP�~뙽x���}����h��	2��(�]�êmz�*�X^�bQƖԵɮ�:iix�m����f2�����Ǆ έ��M��v�K�7i7�26aCt�5"rn�PVR�'��:
�_Ih�cA����Pp�sk�`~O�y�S�}��AiF��N��,��.'l�(�*@(w�Ah�a>�XD�ž�w���Z�Gg'���c�b�5S�T�Vc�X���#6�V��&7ÎA���ua�����e�Ǯ�i�7�D!I�B��hk�ͼ�4+�_gql�n c�F�H"�q 7�lI�#e�i�r�>�[tn�@��Rf�n��("�8�J>Mh�t%�qnҤv���z��0��BT��PB�h��9`|�S�H�+o�`Ea*STRno�wg�u�
�)�{;ęli�����lR+~��WKK9M�ӹ��7vS�u&�^a=��E/z�B�a�[���d�rw~D�R�Ax���Ϧ�Z7�����)�E:+��=�Q�]ŗC*<��� �h�-�<�t��U��m(Go�N	�۝��A�P:��$��v�@^K��̺���?�UH�����w_�:nUi���X�=�ڽ�ױ���XqQPu�R�5�~֞.�F��_q�5����=<~PuM�6�G_��e)��̔2��[��^���B��;oGP/a�0�!�����fy)���Qc��I(e��2B避�!Qʤ�V��IS��u��_���w�p�&�	
��.O@���rQ�,�y#��_��)��R��~4A�EQ#kTލ��r���g����%(�99$�7��,��u.�\��זc4yL*�5+fS	Í�g��=��F^11:���U+b!� ZW�^>%V~�"�9�F���>Wv���o��7�Yb����,v�=R�4L�k�w�@FOP��T�Dщ/u/��O�p�����2�:B�ޟ5�x�g������@C�l%�xt�<�O�2�Vu4�.p�ƆƮ�@���T����d��quLR	�<���S?)�z��=�T�;7�m�Lqa�&�#��f �!M+��'�����`JLc��Gy���V�����-m�e�' s9G��#F�&[�ݼ ��j�rㆯ��g�ٺMX�|Vf�=s}��lL@�����L69✥k%�s)`A9�#b�z�+B����e�^\W�m��¢/nP�%+�F	
:�b7b\�V��,*�@õ�u.�0�y�}��-��[g��yB��tb�|zA���O�����t���&L�
ۚ�M`*�ld��9ɂ��q>��V��D(LP�S��%���*D_�چ#Ko�*r���b�r��hȀ�y@A�)a��Vj
B�,�>�u���lF��/��\�.Z.��u�޽S7�-j�+ ~��`qx}Yt."�[#�{@��x{|2��3pv��Hb]�+�"́_7򒽮����۾!l�Z���v(Eܽ�>�9XY*1���kY��،�5���[��"��n"��\���+(�ӝ�c����bL�`epAW���=p	4C�#Y"�2�E#r;ːY�b�9H�\�q8 �a]����z�U��Ս�շ��JeL��P1�8`�����kʧrt�P���n�5�%���8VЬ���"���[`G��kZn�Ư�2U����r��YO�t���.հ=>G[�̦%S���_�q$����rʇ�H��7P4�i�1`�-+ۄ)a����� w-03jG!�H��Kf #b��V8��Ld*?��i-�k8�l��w��7A�Og����³?�h���g��פ�Y�-8���:�K�s�/ۑ���*��$km��f�́
۪{�	]�	�b�Ef��8M*�HIZ��VI�3]U���G*4W�
'����70�vv�*��?>u�N�Ƣ� j��F#�pPr}����a-�)���D)���W﮿|O}L�����b-
~�K��(�A����S	������v/탑M^�f��QVpѫƏ�E�xl�=�������%^��޺�j��a1���"W�{,S��:E$�������$�p��.�SA���8�]80GՌ��e�od��	(pTp-nYP	��P�����Ҽ��i]v��벾����\7��F
,hv�(��2��ԏv,�x'
��ob�4|�ZV�2�T�+-v�[��T-�ޟ��P*֘w'��^���^\Z��o��v�w�҅¸�ȝ{��߽.�on���6fFC�./����Z�JX��'�єqW8��yS�k.���z��v+�����ٷ�"@�?bc!���ֳŰ��=MM��n�)���f ��.}�+K��9@)�WTS��ϑ���%ٌ���10k���6 ����Д��B��|�)u����=�צ�YJ8�>D�����&vl�gC:Z�Ƶ�Oy{�噷s��n��nj�!/aU��1ߚٚ8{O%���*4�ymh�λ���(�sz�Icz��N׬tf�bҬAe�"[��)`6�a��V�ٟ&��r�ˇ�2ސ�L�6l���-ZX�]��y�@U�X0���3	�y k,�F�nt��>H��(p<��4ۄ&Sҷ�7.�b`��
	�cR7C�ߩ�>G��җ�kO�(qx�
4�:� �Ɂ�霷G��<��0���&8R/O���Sd�nm�W<x�+�ލߗ�%�X٭'�g�:��vsc��)�A9���gȘ�P�,�>���`��待�%W8�]rb���p�rFҳ��z)뢏k�78&6�"��$
����V�s���*0�dˑ"؅���.���2���88|~8��z1X��=A��kuEf9��7��
F�wZ_���D����e}-�KV�k���\�)/j̋�u��r�rl�����jeTH��=�br/o�An(똍dAkXo��6�(?�H�myR,��5<�k;���(Q�(�Q�,g9B�d,C\��L�B\+���
�t)1�2��k��,㲴%:�6+2�K����W�����4LE#9��0�c[Q����J9��\a�h��X�Ȅݠ��I�hhC(l�w�OKC^USՕ>��3ji�L�5�Ba#��	n�A�������aT�ɮM�Ƣ.�Q�ՔKI(ث�\yE>��{�{8�EP��r:w�|�^tW��Z��o�=�ލ�{��įw�ar'���w��Z(�������G��9* R��{���0��u�B�_oS��˝r�/�����X�h�TSׂ�-ϚR6&_�~��%��������P���x��=��ﺘy��\�wA�U��8�f�*��<���Q��c}���i��Zk�H2���P�f� kR����'�&6�<Z�_^O�~u�o�����F�qO�Kd�z�$��t�i�Q�+��^��r(5ɘ�&��3�ډ�"a=�[��s�}+�,���;e�(�쓰j��PwȲ�1K�r��<���]
��o@?[25,:��kٳ�>ї�wLE��	Ye���o�u�i�{�9^��榥͸���H�
�휺O�[��t8t�}`��S�4��밲�r�{?޲�ߥ�w�Bt�4���y�'�5�ŉ���z�[q[9m�k�6��vڦ4^��簮��v_T��m���w>u=��b7<"���0�Pl)۪����X�G�IK���+,�Iaۅ`�x{����.KT����[(���a�uy~�
Ƽ�=��餳U��lou+E�`��(�X����U��6��EwEm�+���Ѣ�����Is	)��`�������p΢�{����2�B�k��n򲀛�`
,��諾��2��;n,7M�^�UQ�F5dq�&$�b����"eJ��D-5 (�CV��0/Ed�E�|�I���T\K<�<[v���r �<����e���x�������7£$���B/am�yk�g<�h���ͯ <��b�����赃*��b�j���T�*�N������%~2�m��4l��-r�=��]29JQ��`�����+�z��_yM�{ǟ),ģ_��o�u���}m��_n��5\��ꚽ>�c�SC4��������EC�,)q�w�zVj�y��� ��YY�rz3�������g=��X��1���	 ���=�H����=�⟇�û5H�X<N�G�+;�,��/����R�>oM�$i�X)P��SZ,ט�����0��ȅ:�τ���#���F65V��	��쫵�����]F��{���s"�y�QI�;y��-�!������wo�i�N�!�➈�I�����4���H6��>�9��	�%�S�[[�/Yѐ���߇���qr<�m���-�6AKL����'px^H~È�Е�׭�9-g�9I&�+���a��u�M�Sy;!�9>�s^g4��8��AI�e+��zlN����d�j�庽�PH� ���hk��������BG��Z��A``b�3��جM���N)[j�Z~�!�$��Q2���t��?�|���[_�I�N���+�"�:u�YbQ B�S��8�`̇}4xHg��U-�v�vɄ��)	D�
2X��6�Q �́�P���VP�}�U��E�]�������̷�|Ϭ�~in�w�+3���n�9�洇��ɣ�;]��3΍�R�z�(;��(A�����J�љۯ/�N2s�;��(�T�����F��5�?�5���.�k�Gx
A��MR�UaI��{?���.��( �!�զ��!�ֶ"����7�<�$�dE���SQ�g[��²���{���8��I57\���!W���yK}�J�x�&@�2i��׊���V��*Е|�B*�i.����?L�������}�'����Ϩ[�y�#��9�k����/bGjޏ�W���+*��\Sז�7/��3��yT苆��c��9��fH�F��L��(+��f4��B�Lt�Gg@�5c�!I\,��yY1�n��x'�%#��,m�,����-.x���t��{
|���ڜ'��s�/�
�KV����=ޕ4�T1=x�F���F�"pp����/�H���:q��P刌XiMGD �8�7%�م-{�����'u�h��*rSۦ t)��`�����^]��ʸ��h�H �:(dI���m<�%PS�����Ir��3��������H�[#Ժ��3l�4���	� G;��Q�}(�y�n*�,�3�
)n�p�/@F8�����K�øy7���تj����.��\�i��	��D&bL��{o/����o�O]��y�����0�Y6�1�꨻�8B)'į�ݞ�&�Z[,�1J�!Uٞ>�|�X��g�>-Г��1m���*����x�fa��;��R�U�k�����b�k�;�Db�r��=�'p<N-W��E�ͬ(�T�b��/8J�ݮq z�ƴ6 ��/x� q��*qSB\WX������b�E_)w
P7js!�H��d������t!�d�ʤ��1#�kR삺�7屗�luS��
f�@�*tc�����-�˛^�pc��x@��	/�e����-�ߥ�G�`1 ���G�'&���g1��X������5�z�T��i-JY�K
GXk�|Z���/M�#��α�_�B��Њ=ﶔo�C��U!ٓ �$$܅zˠ�'T2	=>5��y�?J��W�~>��g-����^{�t��^l�-��n�)�㞂�1�. B#�#e�ݒ3�B=��]��W�	�x(��*�5�`�]HYW�U7޺6@�z�!��&JAK�tE�Zo�&�W��mj�u��Ȋ���ۛ�B�|��eo��Lu�Sf-�܋*p��	&$Ÿ�/�W�z�!e�������n+,RT�j<jfg�<d_V��@鼗,����y���X�i�R��<��l��J����<����Ж琷d�8lx�={�m흮��/NC�@M��C�H���z_.𜍑�(�R'�C��̕7?B~�s�춆<C��ۦS���m�8v��.�k��p�����^�6\Xe���?"<Z���sH��~C�#������;��5-Β���)H�� �
cQ6J�S�ؑ���Y�Ϯ�n�HwD,$Υ�P���)c+\�^�߅�ޕA��=�3���������A���9�Cm7v����,��l�w5D)��_DA]S�E��p����y2�����/Qc9���Ko]��
���N��͋V�R�唢�z�*�흭lk��o�N�/,Z����換?��0�q����aAc
�	y���MH���N�Z� ��]�Y$��d:�O��)`��%����T���ؔ�w����i��U�I���ܥ(���b=ƸT2 M�&��Wo5��B��L�`w�*("����5Ů�/2�/�ى���bT\BLE܉"7�pU�He/<J�1E8Ɩ�d�~�z�����e|x�8����[��9O�g�r̬1Y��*����yΪ3/���?�A��)0�N�jQ���͠�5g�oC;W�<�W��M�1�B��ꐄʻ�}��tB������|�H����������͟��G������9�~�=�su��^G�9�f��n��Ȋz�R8]l��W�sG��ii_��K�{����UdM��԰����W�&&!��|]����ȿ(`~��%��z��D�L-5l��YQ�2�<��h����%3vKƊ0Xm0���3T,����t��F6�����90.-���=j,\3��㪷Q�� t1j
��z���0���n׳��BM��ͩ�'+?7�H�:>�*JR��TP� �S{�B^�kܙ����Ȳx��1�̚�C��6����]B���P�[T�5o���N0&�o���1�g��ƀ0�6��9�S��ғ�4�{��O^��N�O���̷���Y��h_JͲ�l錩_\S!�r�O)rs�U�w�Z#�6�����uAjQqǠ������E��⡘
��;���M�o��7��X��Inb�x~a%8'�I��'d�P�8��RF�&� ���+ܐ'o?|�������������w�ǃ��7�*@,b+�]�,��,�"�d�^�IS�^<;L�L���Q��Q�x	L-3s�> ���5�)��O�'*K?lS�^�3~`��h���A��#�q�l�U)+`�r�N�j�Bk5C�4n,-�,_ݺWYI6X }�v�k|Bֽ�R��siG�fM;�Ķ��
�(h����JW�AʽS���z̶Z�j(�j5���ֳ9���ȭQ`��T��5��5��o��
�k|�6�X�|0�y��(�U:_e����W�7Ew+Wض�Tp}�?��-�d�y�&���]l{-��-���z*)Ѹi��W�ۨ^�w0�8���޽�w����yS3Υ�2U����t~�ƕ����-�p{�y�kn_n!�(L���v?_��;�^�)���F�;9׹7�K➾��*�
^-�nm�ڃV�~�R���0��Y�R�LT�I���w�|y�-��������0CCw��*T�^���]��k�:ry}ss��x�ӷiG���J>��U�g��v����]�\k�G���*�#~*;'Otl�B���o5�i�!����YU2�0D��f,9O朗,�T�k�y�|r���۔� �h=5�璸82���z`d�Z�2.G�rlɩA0��ш�=�p�}�����h�e����o����U����5r�9��?��y�R��O���2�:i��e�x]�y�=p��R�=����ɜۉ�4��p�̨���ߴ�ܴR2��Z"}�yڣn҂�d�ӡsԑ)�����̃8��`.�a��l�z��8��\�~ԟ��SW�;[[s�1��e�uٰ��`7ZuȊI�8!�1�V"�t�!�XX#&u��ӓ{/��Ë��>zA;���*PNʛr\�!�����Tx���b�.�j|{�l�l�Kc+��U�2(�/V�S��k�jW	��\DA$s^��z�V4j��=g�ɑ��B������~��d��M��#��_�RV�ҙ�_<����g(;9.$��pR-T���v<s�|HJ�T����ua�
4(�/P~���?r����knE�"�P��+D��-�=T�F��+���i	z�I]�ϋ��қZ�N��@�\cY��[�BJ|yC�;d{O�7�ۂF�hɣL/S�s�4���O!9�l��ӕr�K�f]5%�扺���ħ����:��бEj�<F]��� �6�`�qd��B(wFAY? �7{�X�k����� �=�.e]^l⿟xtc�#��5X�d]J��SE�T���R-E`*m�*�Y���|�pV)�� ����o�P� 2-P��Ze�<��&�sPɡ��ޱ�͎�U���Wz_f�Ę��_��*�C�SƇG��+ʢ&�ֶx*u���Q$�1:=�N���p�ʛ��2�e�R�}�O�\𪼔2Tؒ4��~����I��D��R�
r�an��O��p���p_{�2�r�/���K�
����n'5F��Y�N��T��=����Wp6��o�L�����)oCvۅ����
��5��0�	�`¾6_���E~x��E|�`�Z�����HN�֠����WnߊMd�'OӬFMy{j�I�^)���A=W��f�ZCYa��!��B�˄(
���X#ί��N���*�ɭР*늿/��H�E����N>س���������ȋ�ksȤ�[�8�c:�x�ԋ\�hV�
H�}DΆ^�L�?��{�>~�G��=c�<�>��N�ȇ�m� ��Mq�Z"�'�MB���I����z�>�ML'�e��������U>,��oii����,k�M�M���/�(\�2���/��we��ۗ�p�qA�؆OvB\H+p+�|�5�{������m
�!u�(
�P���<�w�B��xc�._�5ww�
�q�л��Bn��J�*���5L�fe<:�fҕ�R��#�m�M��ӽ[s��/_�	I��''Q8�0_k���P��H���Lz���a9����ՖA��+rd���{��/��~ٹ��ȔQ�W!�|)x%fwik�ʘ3v��R!��U����M��W��ިm��y�F�ajL+�{� �$���ݝQ�e�J���b��z�Q��=�|�
��>~n1�[l�v%����T���f�4I��;�^J�g�p\�k-ِ���j�1�0Qy�)���#^�Ϣ��h��
�t�e�޷��$V��������u-��U<��o^jƜ�r_T�$ר�蠊Y�c�R2r��v���pOJi�HAͽ���&��^o���Q��b��|`y�r>���V3�:��B��ء�Q,*�A�ᔲ�3�װՙf�Ua٥�
L4�Pņ{p����8�h�ao�[��W�����|q�cI�o���|V�U�|"�cp++NX��4�:��v�g|B/�����7��u,�_GA.�m��o�*�t��&���>��v�Tk�W�/��U�L鋣g%KC�e�9�����q*|�5rW�k>&�{L2]��
q�����g/�jyi��^���lx��=�_쌾�����'SS��\D%5n��3�87V�D�;����|oN�������<������_��������ކ��c69�
�yV;�T�S��aK�|v�R��r��a!�0���H�L��&�#���&��e?��a��15U"Y2���X��l,�;���;P8�8��amq�嫉�]�N�7gx�@�#�*�K$Ӳq/�e��-	����̯-����Z,��O����A� 5�Yvw�Y^�U�7G��g�����t~�p#��8���8��WQ�)���( +?q�� �w����p��_�)]F)4�1���DGnmg��чO��#C��� �,�	ͣW���c�2�0���d�����k�dx�U�(��
_�5�y!1I��&�W�=��_�Y��YT9��Zn��'��q��;�f�7����9�S�^g���1�+Μ�1�qK�|}tC�:�/IG�FK!�1��J/�tE� Q)sϙJ�>�n�6Ϙ��"..�$^��r�+��ps^��=��R\�ĽU�����rY�d&�1�|kt�q�Ls��"Gq"�m���m�A�B:���%��c,k����[8/	�0fa_eCdT���q��k_:�Q�*�k9�&�Iv�{EDӝ�r��_�QM6�����^�%Z�����"?�G����O��9d?���ԝ��F[5�\�i�I���&ŐB4Vuۦ_����������{̴V�(�)1����|1xIV�u��)�jUi����4��;�b^��^���vC���J�����7�'{T}��ye]]̑���\ۅ�IܑYڐ��Wd�Z��8?�ɖ��E𬶫�6�`�n9���#\U�������s����p�C9��P��j��z>Y�:�h{�φ���mL����^NO��.(hn��ac��y�saQj<B�5o�cgv"bQNym���x�{�3xv�|O������bq������ְG*[n��r
�Bp��~%{�cyǇ�����;�i�k?k	�T�!�
�1P7q]�Z�:R0�sJ*)�R/����˒��>��/Z��&�;��5^d�b����ט�i���/�Lm�`L��B��p�M��k���C�+T�b1v]r��+�^%Ӝ�"ՔPW�OUtM엳��+X�7��mg���D�#��l��lJ%Z��
t��c��8f���Cm
/$����`��������%D�����k�;,�"
W=i�NT�.����^���M
SXA�k�)�N��)A�h
9>�EV�A���Iy�
}=�Xox]GҞ�u�Mz#�:��~;�w���F�Ջ����UQ4��Gʟ+v��3r� J�X��Z�^�� ��xY�3~�+�X�B��t�=0x�$��U���qR�4��mu�k�U��y�H�`X!(ђt�J��
�%�����>��e�_*J�;MN�g͈�8��ߤ)�[kJ�u`���P4:%���%奤E�D(��-��S1�+�c��y�?l��"f���F���R����g���g���Fmu"��m��:��,�ޫȒZ�3ɦ��!��k1pLIb�̚jv����"�f)�U�WV:�&�!�T�k��䐞aȋ �P`�Hx815��_���+W�� �mAe�C8CVy;A��<?�<�}�(��vj(e"��Zc�����ЫȨ���ꡛ��{e�����:���M�uh���=��>����g�Q	��h���C`�ԖW��� D/�
T� B�����+����qm��k�"���k�H���)?>u������}6{vy�^]�\���D%d�?S)�MYR��j�oJl�pb�\�,pى��]`'nl�>���N������;8�5�}�˦7^�MXH��v��։F�&c��ia>~A<����C&{�����Znv�_����6v�m,s��������Z�3'�[A����Ū2�Rt������}���5��8�����V��U��ɀ��X7��'ڏWag�_� BF����o��f�)�C�B��H9N��{(��3đ�x@B�3F,Ϫ@�:��^�9sS�gA��:k��Xנb=��Ơ�aT�$?�U�����\�K��x�*���ve�S���e�jIk$�(܈2���S��˪ T(�bl͓�OH��V�*�6Iqltk�[y̞�����Qel�e�sG���]kC��Gb�mNr�9n
y��$ˇ�o#�)�y�����h��~F�4 �_72?mhc���/%輔�7�Ga-?A�0Z�Q�����������;�k�s����x�G<^fC$ ���ڗ��rM�ik}f��:ͅ.#%F�d�x�E��c�|�pL���Me��)��4���[#'�"�Y�jѡ)�P��Υ��iZ0����˫�����z!���;�+9D^7FzG�b�yC��]L5Ө a�x���ϵ��aI ��oJ�+eP�:6�1�K�&����*vc��.�mov4p�n��X�$^�����O|�m\~b9�s:���������x�T%�i�ΪTXbU���mK��m=�W���08q�W�L׸&�5B��c�3�Y�>g)�����p�e��_�a�H�KN��C�)�WTǣ�\z?���p=I��P�EF� ":%�Ǜ�����;��)�'�/}�� ��ݞQ4����Ԅ/�����J��4raZ}D$Yb����n}�����	><��E�����4�PRX��EE���F�K��*R͈�%�Ն%����'B�pOl�Bm5ǣ|t�X4z��0�:��Q9���WS�z�dk�P�&֠^#�E��T,�M����jM�c^��	���Ϩ����O��u�)p���uCIZ�̮���`W0��ƈ£��5��!U���d��>P޴�Uf|�G�{�{-��c�$i¸,�[�7��
>ʷ�ֽE٭n$3�l��𬩼c�/s}��41�U�MI�X%^J@EXHY��-si:�JZk�E��������!�B���CJ����1�5!�F^��Sco3����a/�}d<��
������/�S��s}3��O�{���(��?��p��0���#����@� Jo�����m���+�_Ӆ,�Spp|A�띿{�{���'<�$�ލ8�A���Ӊ�{.4��NjH�D��sg�(�o�e�1��ү�c:��z��C�����C%���Z��ݠRY��l�����u�T^2�SD5� rPL����g����Ņ*��&k)e.��������4k���
,1���5F�ې������V��x^JPf�*V��$�SH5a�o|��wq��醶M��UK�"�,+�����M]�#R��h��$�Z�GYW��:��ø����:a�c
sA�"�������p���",J����lz�s�N����6�A�r�g.��R���x:EO�����8P͸y0OkT����Q�� �����������{���r5Z��|k�ս�����F<�w�޿.�{gW0
VW���Na�eG�%o�i�L��
+�5��qBӓ��E�ߒ�(w��v`�O?��|D7���)�F�/�j𬖖�j��?e�BR�}�M��"T��_�1o�n��N�Ш���/�n@�vV�;j2�q{<K��V}Yz
FA��v���կ27>o� ����-7�9�K��қ[��e��\��&�Ǳb�ݢ�����Ҫ��N�%EҙIx)�)�`E$�U�/���g�b"��G��`�
�����,�)X�\�W~��v�~�}}��I��9,��4�)�(�vo���R���su��|`�oS�?l鄄��`4��@�K_�t�-���Ox�B��ʂ�(Q)zϔ��$ju��24�5cm�K�/+���^Pփ�F�?o�����:��""-�z!F����K��a(@���i�U��22�QyMO��
�x{W����d7���z�d`i9��k�34U��O��;fo��A�5
���>+6�jj�A��g��c5�.�U%�Y1^�7W�.Ť��*7���OJc� 
}E�>΅�SB�=lѕ}P�̥/ 6Cq&Tt"�*n����81�����n�9�+�>�/Ah]Ҩ��)a�@���*���0�H�&���Ѕ��9�Z9BeO{��n��A	Q⛛��d�u��]m��[Þ���߿��ڔz��+�.� @�7����Ͻ��oI��Ͷ�H�
���L���	�|{��?<x��=�b�^�	��!�����!@V�apà����g����KR�a�[b���਽�Ծ K1���2n�4�f��)�����
ԙ�6���b>Z�~����7��ވB������ꏩ�~6�=�L�����6����;�?��ɾ�[�D��N6���;E�TS�VQ\��=_x������^�`�)�� o]��,ذbY���85�Ie�"�s����&)�q��d1M(����8nAH�rP
شT���!֔�\Of_���A,��`T��$[>��cT��j"!ĖEUZt��i�=�x��3S:���lr�y�p��}��M,L�o2�M֦���5�V���ήh�P�7�hd~�ЏP-A�R��\Q�/���ע��D-a�æl`�{JB��Y�����{�y�}����:�% �s�Y0�-s��7��{<5c���ҡ:�\�4(� 	@��}	u�>�X��Yy��V�k$�wC\m:BN�/ǽ*,�SyQ]A9�d&�R�Q�΋��.��NQ���3�hjsY�^�m6��q����{�Qw�=�*7���ʲR�ի?rܺ��v#��Jij�Z\��� ƪ�m-����
�u��o�h����;sŸu�rW��xJ ++���|���Ŭ�F����V4����n�{A���ʗ�����&(�����:"G�����&jͪ�M4����ʽq�W��k�ҷ1��]�.�L��3�X��E�@��R��,��	��)��3�&�� ���w+R�"2[(��v�n&,��`���TC��y�ɘ����ʭ}1^'�E��s�q#W`�Nk46![��ypf�zh(�7�1���:��w�ŢrpR���c�L��)qv���ֿ�����_xJjq5���� M���ٯ�/��D�iU�uN��D9:8<�*q��a�W��ǵ����������N|��[�,��-��p�,���*�"#t�M96׮��`�8��y���x��o���G�<y>����οqM����D��'���a�/s�«� f�pB�6��meHD������go>��*r�	���C���hwju{\n�)bc��k�bL�ǒ����Y(=���y 	���ͣ�J=��l׬Yܙ�~[v���h������
����GaFh7ƭ�:�)Pkc�5
�W�#��"�#�O�K��c]sW��1�W�^3O6���a6�径�1�.�7a��gxy���6T$"�A�uC�)�X1��=ںKS�1�����[Q|�f���C�}�w��p����J��Y�~�~,�4xyl
�"���v��k�B/�z���vxoT��1 z�"-��Y�{W�z9w��IK�R>��V�m�#��ki�]���M<�>�u�)���4��ٸ�I���~G����m2l�
��#�m
�W���Kf�����+~���޵����7+�U�9������	Jэ|�����ss�D��K�:��Ұ:�oJ����(P���c ���������0ݾ��܋U�ٿky���^so��{,�T+~��^�>צ7&z�'j�UCB�"�!���%��x�i���4D����i]�w ��4��\/�"��SoQ,�����Z]�؆P�l�{�Ҭvţ�$��B:�;v�OҾY�`Q�n��������g[S��E�,������_�k\e~����9J�B�@B <��4	r�(�{A4}�}l��a:*J~s�pm`��ω�/~��ާ��:Ȫ��08��tAV�]�}�X�Q�AP4"���z#S��#�d0c�@V�~��Wr��F�'��[P�
cd��6���lo��`�/��V�����N����y���y�g���7������_��_��_����.]�4�{�b�-�uدK$���B�E�Nen6���d���9�� ��q�q�Љ�����/�ф�����(�rd^a���8�*����m�2�{���N�λ�mζ��i�gXg@V3*��a@�r�-�[)`ՠ4�y�@!��j��w��� �����l^Y<�b[+i^Y�M����V�sU��l5���lLV�V����S�Yr1;�'dx�f�[Rv����v�����BK�F�Q4B�sOB�Q�x�Ƒ�xC&i9��B��m�몾<-��=ՈΦ�g��c��n��(��T�Bl�ܝ��2#*�+*�)�BJy�O�E���ౘJ�W%)�.E:j�F2��ˎG͵�P����[��=�ŊS�)j����Jo^]K
mh�vK�]{<�3��vR��t�c�*�6���feԾ�ZW�M�3k\n�홣ys�VK����������p��R{��Z4���������mו�Þ�+�|>猂�����%CO���rv�yKDL�.���0Q�:�n{3����j5��F��w����7C�֡2�e��C���y��Gr��^CA�c(�ț��ѵ�������MN|6,�/7�\�_��*�6��w�41��l�(p|<�b%�KZ#�fv	��K`z|I���\쩎򐲭����-��x�*,��&�Ԍ# �sfr�/ �	�G�Q��G�VZqy�\��?l3��#�Ѐ�0�2�c�����0��y�h��ӝ�{Owa���s��k�%YMz��U:���/�#sY�~׮a�U�G����T��X�n��!b8%�{Ӯy��kz��a�oռ����0���M�N�[�?����']z}�?߈B�"����'�����~����������ۈ^��L�Mj�h�4-H�Ǫ�ee2*���,�0��؊(��%0���{����4{�Q0]��@���.���wmd[��5
�V}2�K3M��UP)M!5)�5�� ,ұ����H/�xT�;@�I6]*&'?{�v��A�H>�� ^i6�pTR�R�`�U�{U�y�>�DD�l��)/�dV�Ⳬ0=-أ"q�z�U��+�%4���
���>�XK���,� ��8p��8&�#%qy�'Ӿ���_�ǵ3V ZD��)T��+�"e�ش���X�X{TgA�n��Ċ�E�F��Do�"j��4Uc#x�Y�r���)~'!פ��Y��5�<%,��&��UB�{�a�N(n� ����b/��1��{�A��Gb�����]��X�q���5��ax/!�9[̽s��̅3�Y����a���o(�{�w�T���fB�F}����[)E}�Tg���_�?�"�-��.߶���Gۚ�ߔY��F�1��Z*~j�&�K�� ��Q�b>�zr_
�����}���ᕬ�B5����VM�������W�w��n�ϓ��>�Ӭ�*�����3D�1�C�7��e/T��r ��8A�_F�e����2��m�^�EL%oEL���_�#u�.g:0���p8��c�
�eCm��M��u`��e(�m��-�rK�1�6����5N%�Q2�f**t�l%�sWD>i���La�́�򦅪k�9�5Y�>�A���b�����ዏ��`�>��/��x���^��y�p����3?�Yr�2�C:�I�[NA��0�|=�&�ɱ����Λ5U���|s��!������.*+^�V�c��7G��N���)���!"?i�jF{��|ao�������7���y�~�`{�����W��߷'�-�f��Yw�\f�%JpALW�;0֭7����4!�:�arc"�k}ko���'�6�������#n��bS��)V\�qVڪ��ɱ ��ɃZ@���������+��3Hz;ԁ�����3]�$�I:�_�<w��{��{�m��P�����J� �l
����vl��[��1�UHj��7�]X�V�â�Yɵ�Lwe�$�:o5F9�w	�a�����M���G���9�,����kJ1�]BQ_'�>ȃ��pq)��q�zYnޔ�mם�s��Tt���^���Ԕm��O�~W�<�a+�ߴ`��iU(��D^^~	ډ�	�mPq�(�x_B��y�(F?�Y�h1�a):�+(���J���{�U�����}w�^_#hB3����(el���
�x{�k��<g�Ap��G;O>ѿ�F��䖺��FT.6�T�q�)THO�Mʠˑ*�Y����Q���Gҟ����P�0�mWE]z��j\){Y���d~�}Z�֧03�I���@��#�ߍ$��kc��0���O�2���sR�ߚ��)k�*�h?1c��hl��Q�3��9ETj~��D7���ݺ���P�� �I�u`�|Xe�Fe<����x.,>Q�I;�29$bİ��
}�R��k��%O�L�%�P���NPhgTw�s ͐�t�r`l��cQ7�=
���=e�4� ��*�s)��x��11���.A�/����~�ele�QM�99���&�}�.r�E(�!�^Y������q�p�b�9�g��ֶ�[��_�x���$�R�**7�b4����Ԅ������N�	ɚ��У[�� T��Ǐvߘw�hߘB��/�L����?��ǿ{����ϳ�wc����Uoci�x�B_��&,��,bB	�X��x�
7��U6���C,�����)7���17��l���,�e�k�R=sY��j�n0�H��>��êu��&��y��lu9��}�%�	o�o��|V��z�9�EHλF�6���x����G��VAzϽ�BJ��*hQ^d���!I�(Xw�
Rʜ�V Ŝ-�.�4�Z�:2;;V����x����z-B�.`�د�@��N�ñ�Aڝ��IJ��N�@\��I��}!�4^/�ы�T������ރ䣸����1'��^OV^~��5.B�S�+V�&�W�?~�|���J�k�cޟ�Ns���m�YH鮊&�ś�{Ԉ[�n)�~��p����q���h�Id��S�M�4K/�eW���dr���݃/�7��@�G'ʼ�vw�� m���|=�֝(�U���sFM3GUE-,�\_�F�f2dL�VJc>[�)~�
�`eŕqẋ^�x�_�t�Z��Ю���PԫbЍP�{�Th���h��*:���)0�����.�nz�퐲E������,�k³ň�h�4�K��k2X.QL*�\��fz ���ly59F�@겔��PG�ir=\ ��֭v/���.�鴶/E��F�\�y����q#��:�ehr	X|�z�Ŝ"g��Do��j�=�+�� V'���ʒ�2�_Ȅ&�$󧒜qM����i���<�:G�[s>�W���}�����~��t�S� G�,Q�~'<:"�?��V�C��Cq2�c<Ʊ;�m��{ِ����/�r4:8��� �Y*}�c�1jt����B2G	Q�q}Dq��.�������λ�o,~�zyc
ݓ��ϼ��_��������/l ��#hަޱ��_;��(������˨(S7�Uij�R��p-�����o �ms��o=L����=#�B��<p���;�R�,��%*T�q!U�`�W��i,h)���T�,����e��~��xx�t�MHs�k���F7�	�Ք������p�/�FB�5:d���a��^F��Nr�#����𽊩)?+�6'��".��z�(Y��`0]ːMq\����YXS��)�Kk��"*�X��O�>�p� dU��x�r��Kr<��/��k]Y̨���[�����4�ؤ��.A�\;�"Yޭ2���^-.[��{*�Fv�B�9l�2��j�>����Ֆ���=)�*���@�I�jFA�_��DX��3.����_g+���uod�"��X�������z�����罫�x�5�R?��j�G��R
�����2n�U�s��th��S���&���#�6�ħQ�gp�z�8ϫQ�~��S��M��z�M�gG�,���X��/�n}/4�CNz��Sї�N���4�d�e�J�2+=����VFxS�����@Bd�k\r��Ʌ���֤�9u�1,vd���olյ!*dI��j��Y��J��%h���9����p�6B�+f^HrL����08���V�]��ő��79�h�
�
k�Y�������_j�s�����xV�<:��vJ����{�>|	��-Ҏ��M;A&ـJD�9�G���1R��-d�h��^�b��cu|D�w��fN��4���6���8{���P�w����+^$���<_�|�������#O#��!ۆח���ww֯~�����g?r1
o�Q������wƗ�s���e�b��r����&2�ױ�ֱ&�W��S���Nܸ�IP����9�2X�K������=x�ƫJq���$=f��j�ysb��y,��M�rO�/����֛
�.�+ޓ0W,Zs�ݐlb�]@�*�D���z7� ��͜հ�RX��^X�z�*vIx+�E�=�Fت0o�.M��0�@.��,��UM�*<�q�ě��6܍�V��4�^��M�*�����-;{j�����H`�Uzm�r���_����B�2�2N�?�sD*��&`U9��N��R�*����&��{i���P���q[�OekHP���A�wz���g2�Vk^w�L�������4�}���<�sV�z�(>ʻ�s}2Ɲ�k���M_HB@�n����i�P��a�~%����*��������3��e7�/׸���ݸ�{�Q�?�A���^Q�8"5V��9�,�璇7Ю���O{G��Fi��I�0������9rj�{��$�v/���V�����{SU!��B�Oh@��.��ww��\��g��,*�L�#	�U�^%f:��ɹ�
s�=8C��x�(�+�
�S-U��� J�\����"Q<g������O"��6���hq�y_g�!����y@��9�c���XV��M���9cS~���~6���О�"����v^�v�(%OftO[!vA�}2;C|fY�˓�����/�����O��_s�/�����X��ΐ��W�L�V�� d��%������#�d�)�Q�.��>�^�_s�� �ܯ��bź�sN��5A��4��K'yϊ�WGG� �����Ú����yt�||3;���}q���6���*�_������?��~��7��f������6��(A��^�U������4�Wѭ!Eq	�2�Dqؙ,eQ��#*��J�� �b��E<}n�����,N���XK�M:�I���V+Y��j�ź5�U��+*���{{���wK��V����4
�lB���0����w�B�R�8�0��W$���`����*�d�
g<|��Fi��_av7%�k#��
�JK�\7�L��;F��;2���ld� _*37�)�'Q2i 7�P�G,o��3�ؾ��U;������+��Ni���-$�eU�x�E&���"�`�Z5Tjn%��趇qi����Y��~����˹��AS���`���j�����W�S��cv=�ɐGTWCJY���A\~�v�K\ʸ���)>Qv_ѷ��w���#����be󀻛^�W���#������k)#)m|Ew�튇�N%y�~�9�U<�����5R���kIcu�����uWC��㝚�V�uM%��ײ��b%�j|�O?�O�bN"Y���и5�[��4T�T(2���@���<VL[��ꦴ%�Ƞj�d�@q�W�J|e�;��'��%]��e���@��=3v8�䱴��0>,�Y��I)S��׭_;>�y������OKt��jiX��y)xރ��dndӧ̫
�c��9�$��!�x��j��u	�)�,�}rl��	�/�����{�/������Vj�+of��!��#*�=C~����Nwv�k�=��4��0�]������/r�2�Et���[�s��f��7�?�x��͸��;WYe�O<p>szB76��܊�R����M<|I��t�Y�/�C����?��Wm���oT�{տ�k���;��wN/'����������% H.�u��"������Kn��2�o���
�(����(|����eb0*�Mn� ��W^�p|��h�E����Q�d�Cm)l�e7V>�,�%��e0W3�c1(=|ٶ�	_J[F�TSR݆PMҼ����LH6
�j՘�bj�
"*%+^���b�o\�n/{�� �>MaF��'S)q+M�\B(��t�5s���/	9H�I꟡��]�0BM�#��|�H�1�e����-3�Ҷ,��+��R�lUgjW��(~�6�y�еCe6��K^��Ɨ�*�.�"-�F�#T�B(~/ex�bj�w�ZSn��R<��-��wg�h�ŝߡ[��?��Ԕ���=��aM�y�塽�h���%AW����:n�	��-�=k$!�[�O��V����[%�����[���w�
�x3bWd*������cS���Q�*�~�:'b(��J?�oH9�J�lƄ�|{�b�Q�m�~:?����B�hFU��r	K�*�?���t�-��P��c֖���5��̆���"�:��z�_E�{7�qi\��V�?�Q��f�r�'T�z�d�Y��@X��#r,�l�Ժ �6s�e��9'���d��f6���>�HQ2���F�:?gx�YB�
���0�C~U�h<�)����p�k&s���98�W���87�pN��k���eڪ>���T4X�,�̶���m��c�H�` v��LT����󙆋��1�9ohv
,B��D����'1W$a��82�w�7��-�+g�Ba�q�G�)���U���8���AR%on����ﱍ��9�:���������������h�ܻ��������?����k�9����������5pȄ��S�M8���w��?S*���Y�^I�r�)ԭ%�x3)
l×��҇�vk{��p?7���>�:�s��6����`��)�<��y���F�q/���A:�{���e�[k�CȐz��3���|j#�%�B�kJS,��/�5��J�i�5��Qb�J����p�Xn��
9�F�1'�	�o�
����]e2;�6��lU3*�.�PqH��o������nP�lK����Ϛ���*$P������H��[𑘟�/�o��@�B��evb��kC�#�3���3�\�����BR��;̬��؉i���i�D���#����2ར;߶��ͣ��KA�[5�y����.X91�F��~A��u<�&�gɁ��{��q4���}c.��Qy�����ش��Қ=F_�"��A߇�}=Q�#�K�cA�m�5����x,`c�H�ˠ���c/-����m��W�`��%~�x��}����&��]��ٽ��
�O���j�Zʷ
�C���;�P��I�x=�=��7׽9Ё��X�$��Xv�*e� {��
�X�_������������������*뤖T[#�Y2�8�u٧�.}�n�*��d�_��v�Dx���MXQM�4W�Sg&�� Kx�F�>!47��
���CHlo��~���i������:��tp�g~��z	��c8N/�bZ��u|���OR[8Źo�6��4G״�3C|Lv�c�! "j�Z�Ro~�+�!�;E.��(��-��Ԛ��c�k��>�V���Y�1J_�N����;�����]��|k�����_y����n;���޸B���������~kiy�' v�Req��4�z�2I��bZ�,������ׄ����t�"�b�]�wt�}u}v���6����wz��&�t���-���P�U��=�K9Jʰ��;���9���o
=�޵���v��Q��-��4���Flv�܆\��ט��^~�^u��M��<z~F.O=�'TVZ�����OO��r���,e��^��za��Jh�VQ�6�1�M/E�8�Jv���B*q�&� ��R�B�Q(iQ�(kvߢ����9�BZ�ɓU��W�ϔ��O{/���S��<�Ook�,����y����%�(�LK��w�8aIa�@���o,��7C�N<�BiR8
��V=�s�����*o���GY_�Hi�G�=ڭBw�T���=����P���·�F��1Z�@kk��z�]��y�Еt����,u�R����w1m�n�H#6$I{xg�j�hhȉ<�c݆Ñ\'Q�Y[*�R��W�J�?�N-�,v�^�S�Ë1��=U{�P��=�k�a�7^ǰ@�E��+�b�є'�b��ҍ��?T�ًd��Y�+�o�5�S�ąP�*UܼIz��K烱ٜ��8�����>�3K��������y��c�J	�3�v?S.J����q]*�����R$��Ekd��S��53"�΍a��jWJ��S z	u�������}�5x��[�/��h���wo��D��[T��sz��d�B9O�1�̓��Gצn&�g_j�B>e���s�}sDl}�f�P���mo�)�:��&�a�Q;�l7���2%��x�?\ي�}����\�[�r��qF��iz����l �+��x�����0���������c�~&��~������?��G�~���o�7v�.�)qa�k�:�������쬕Ȳ�;�"��!`�c���N�&&aNKw�����ǏӃW���/_P9���bg��C�!6L��[�P��6פKリ/sۛ�!N���b��e�%	,5�ab�Ѯl�I��&u"݊�2�ӏ%��vc�Cr��8/ff�g��P`uqj�,�Ü�V��y��BڳK�NDR�&��%�����k��Uo̴��
Eo�L�\�n����Q3��Q ��̩�()�)4��a<��æQؕ�cn<����fc#Wl��v��k#XE#$���^z	��V�U�S�)6�(q=kW[��G/S��/��5F��q�|�zC�����xl����O*�;?J����~���k?@��S�H�����ǺU`�����#�u{��P��۳
�?�Bj_���	��pN�ex�l��Ё�X��wŷ��wg��٪�5cK�}��x�M�g=T�[���>��{���p5������)��`��hֈ}��d�g?�y��1�WiN��,���0eݯv�]�qO�_��WA��˝Kc��>tmc�h�Q����FNh�$�'4{�M=�p^�w�(H������e1ԋ<�w��[ķD�b 8��O�-碪�I��,b����{�����_��у���{��@�� e�WY���ꂾ同^�^v�����}�Ej�A�|%�,��9��-b{F��3������g	�kݸ9a�m��%��Y�f���i8׹c�c��:�kLZ��2���勃d�T��=QF #��,N�o�N��/�ԗ>�S�ާ��gB���۫��o~�?z���j���Kk�w��������YXcn��6
d����%qmn?�<��ã�j�i6��Y#e���z�)�o�o2$1�o�^u�W�vC������nD��-�m�!�X��vS������˅�2p�H$��B��Ά����~i��Ѓ �R�`A�Y�-��I�D������0�2�k��GR9��MW^���Zȭ����������0qG�5e�e�~���aG�1n����oM[J6�`��)vsW���ě@0���k�`^�XW��`?��Fbi7
�8>r�L��9���	�b���j��Z`�ټ�"�OS��K!+�Y���ͦ|E�����	V8���N59?.�$�V��l�����2����Y��)��?��I;~_�X���:���w�?!B�C�{ݕ���?��]~)�i�����q��rW�7H��!��.�����Ve��sY� <b���YÅ)X\*�A9*�U|���s�Ez�\��)�z�U��I 7��������X��c�r0I^�s�릛��M'3�.Y'#Y1x���]K�E;V�rCm"@6W�Lh��̹�	�'�Q��~
�M��.�M^�[G�1�1���5��y�2�a�Z�m����2/ҠYE�S׀:"��9�H����8*@{�Y����p��g�/��m3mn����l~�K�_���nc���LlqJ\�������nhu)!�=as�Q�xӅ��ɠ"�z�~�����d/�N�ГF��	�˘H|~�#|k�s�Ó#�L0>�7G���*�޹�@q�d-I\"��v����u�T����d<8�͟}o�����מ��Ė{c~&�W���γ���o���?y����wV�{�� G*�7��;�1�|*����������S#��-s��n�L#�j�w�Rһ���F����Tb���w�!��qM9A��N���<xO���-�r�n8n�V�^ 0��c���f|�:I[�X�n7@5pY�+w��u�f�z�j���f�uә/i�5�[��;N�:�[��7�V�Ҕ��\R�#��̉�V��{b������Q���)�����ĳь�'�p�`J�=�UѮBU_���K�Ak� "_g錰jtzv�ӳ���������UbS>��Sy��}�S�z� 3]_/Ң��dj��|~�����7ǊqӼ���:�m^sS�����E�\��<�kkX�?�}3��x����U�3
~�Ǟ+����*w�:�����nS"�`�B�P�Ա��^�����$�h���|TE�:l7 +�)l�H��WZg��*,���2�T]󂆵yJ��ܛf���5t(3���h�
w���������{�a�)SJ�u���fC$�WCQ�����nmz3� ��B2�Y|�:��A��J)�6�O�Z�+�`peJ�� ��S�&}*5��O;�a������k<�m;?�A�[8�s�@� ��������:�E�"m*���a���\4µzA����k�.��Cj��������l�{۸5y����Ū΁Ǐ��)���-�o�����[.�S�Q}���̝[/�jq��/Ďm�R�9����<�ۑ|���p�0�S�������]��)ykm�jO�Ϟ=�VcLp��4*�r�M�{�+������Ճ��+?����oK$|&�����o�����������&�ᧇ��[v>�b�Y��{���@1�u����w�78�����,f��@��-<G����%�:\*B>���	����8cُ��>�srY���ø��UM��q/���i��}=�tc��c�iY��ܐ����<�e6H|6�ǘx:�	#��n��)L�5�]�ց�T\��h�ڦ/��YC`ܲ�UJ���L^-�-�.ϳ������Y)̶�]�1l���2V�PR=����~�}��8hh0tVz`�^,h[aeU,Y�z��������
��:z-M)5ѽ��c���0�^'��z��6�)B��(HYV�wΧ��&�2c�9S�������vC���깼���}?_Qd����I�A���T���b����}�ӟ�����+�y��E��x��]7"jq�{q�73��:U�}'F�
�)l�OUR�Zt��A��QƵ�|�|3r���W)duL��D��˛*�[W�k/�+W���J�}���Z�]J�{�_k�o«Qq�|���v�υ��Ծ�3ҳ��|�t3��J�TR�Ԑ�ĵ\WCT^"d	O1��44����y���Q2�I��P�N>3c1��3ʀf��8q�3֘p�@�ɛ6.��ɴ��t�"'2-������b��6h�\�)�eW8Y3�:,擿��������G����6���"28^x�vI�y˹�=��i���y�h�h�$�s���q.Ɏ<�+��3��5xP2�W�owk8�G/l ;� ���ݭUG/0�$��QK޼~�/}�k������=�qF��&�w���@�}���p�|�����_��������Ol�7��gF�;?�շ^|������W�z|v��hu|���=N��)�|r����������@�����1e��X��ȫn0F��	����������R�vv��'P��-|
�b����)ؿ����,SR�F�U�o	b��n_`��%뤟q����� gV�Da�E89dY�.D��q�x���l&ٙ
��uc=ש��"���"����T�{K�al��5�Eǈ��#�dT�n�F�R����҂O<�����TĊM�*�"T�	Yi����&��o��x��4!�&�\c1��F�O�`��*�����A=x�B)�u'~YT�>%2�Q��7�i�.��n�ċ&N����n�4�je^4�L*x<$����&2���Q"�>Bv�=.�w�Iw)J�yY��ތ���T��?>���0�>�����J��������nyw����w�{7�* S�B�ڷ/Du%[�3�R#V�4��uiո�UF/�9���ÀM�ʧ�cZ����������]�ʏ�Y����R�z��i{��\�&E�Y��9�K�2\�@�s4ԃP7��/�-�<v-MS�4�{��j���(.�-)ҙ��Sҗ�Q�2����n~����ǹ���ۗp?b4�z!Au��Y��w�~�F�]PF�7�ص&�""���k"W �p�w�.��%�@AJJ~ Z�nh_�����'8D��m�j�����k���0z�2?&�\F{ڷ�S��/!Xc>dYɄ�r|��	�=K�Nl�r
���4��'ǰr�������8 �u�Ω���g�O��90:vۛP1sɇ��΄�=^�']���ޣ�~7�A�kjT�T�bS8@������?�?����k�����R�����_����o��?�W�77��
~[ot���D�������6��Ͽ�����z��?��R�X؆%!	�����{�<O����g�[����/��v�c��.bh�rnc����&y��4u����b<C^<�����ݮ����e��d��s�w7Z�K7���l"7l-�t	K��M̃6�"e�ܞIM��!e�c*��uk1W�����v`]:3�Oȭ��x�w�
�M3�A	�t���\�`�	۱����P�tЂ�ߊ��BtG���~����bα�*W��eC�smIGXc�G�kD�Bg�����P�x�b��OV����C|ھ�<�����5���e5e\K�PK4""
#s�=�
{�IV��g	Ȉ�� H9_����*���`�N��"��n��'��� ��2����l�K���rH����^y�k�YC���b+�nx��-T{��/���Ћ"	���\A^Ja]��t/�y��x��ī�j�)��Wp�_F9rY7j��5\r9��&��F�X5׉�p=ܯBN��+$lC������G��5�S.e3��7� 3*��"1�'O�׸ߗx���]����7�:�1�?���r]1Se���T�	=���=��������;I��\�o�ۦ������wۗ��$�p씛6��=�I�
�[U��c�R���}�#ZG��h��]JkC0޲�<��9���/����2E[ S f�f��L.�\��Z *��vG�͈�pi���0 �?F�eam �X6�.[��_�����x��v�J�3V~¹�ALY֐X�d��r�f�8y^�������̓�e*t������,��f,��=����r�t�w��>��^x�����?���������?���H�}n89�Z�������/������zw���'ϩ�NE8{�ºY�/ؼ��r�1>��Fs:~U�+�E.��7�N���$6d[Gi� �,�kfZ�x�S�.T�z$�%�$
�*Q%8#4��yS�Z,�w����_,.ܤ�J�*79�-���0UB�����*]W�,
��^�6��"�$�p�:8C-v��S�E*��|��u�+�~	�4����N�9�!�P���a�@����R+�!^wZ8&�Z��ƀ�%����!¸b�
���]~�p罓�R���tg�Ѹ�\�w��g

׻�`3�N��kDO�<{7q,y�!ʐ�
^/|��V�*i�^읷�Y1�.b�5eڈi�=O��Ž�t�o�8��#�mz��
%@dK�G+لv�z�h�����2���{��o��������g�Z�MW�yCF4��jo���i�!�l�Dg9�m�#�d�oQj*�@��u����<��1SJ����7֝=�gA��:w���J�tZ���̫ͨ,l��~��W����rJ�"'|�97�K��j�t}7H�O_�T�x`����M�O�$��]an���]詇;�k��[sAY�}�j��3�!�X
[R_�e�֘t8�Ґ�f�˫Ƙ� �H|\كW
(8xH|�1U5?z��L (d�}�� �͹�!ub���S�3+f�l��!z��ȩ7{�Њ2!mn!�^� ����h�a�Ūm�G�:R�~4�m/1���گ��mXVΥ��]�9�lu�If�C���G�3��q�W�>F^&Mn込�)C���0��[��i�c�������O��_�����/|n������ϜBw&~��=���?��o=_��	����XV�E��`��S������ӽ��w���W���.�ij
���q��G�'�Բ�EdUT�33e✿�2�j
�8Ўj1�b�955+)��������hBӠT,����2�J������w�Z�S�P"\�Ҭ"F_~�d�K�����=c���`�d����]��=}�5�Q7�Ƈ1|L�1mNb��úհ�/���r���Ŋ��N���Q�%0|���q���S��7��Wش=C,�7���Rf6���b�y�l_�M�`
���/�i~��"�֌��A�c��jwV���
^�$(נ@P�c(]5R��]�k��2$$#90�U�>���|zы8�*4��5� @���(�Eɰ;T�s��n�p)�R^u}a��w�����Q���=;��FQ�6OŹ���C�%���u���̉OUŚ���0�e;�����M}���C|����8�+��tkhxo���VY��I�c�Σ��<��UfM��~56���2F�����e�w�2�
3\�l� �}�@&rT���N��JK�����U������S�h�ñ�e��zuW���$.��2ã���VGU�tD�B���XNϛ�M�
��M�s���=����	5-xE������CJh�nA8#�ȴͨ��8_�pF�rd��P�gTa;��-�]�M���� 
�Tqjp�S�ĬW��ƻ!�1�IϨ�.�Be^�n��4�Z<������Hpi���V��bLc��S�l���we$5���3��&�է8k�5A^[vw}ydf���2g��s�S�0�W����ş�ܓ����v>S��ZPI���=~�����{��هgic��ӳ��heeEc�z����3�{[���?�dp2?|���, �x,7F\�����5��b%��P������3,�Z�4D+��&z�X�,p��c�K�� ���&rZ��Z�W��8�1slHs���+����:Ʌ�#$�)l���	z�Vċ�,�5��B�vd�y�Ǯe�8b@H2�tj9�mpcaz�c����W� �_�A�y	WSj�\�j�P%��CeV����S��֐��q�����2�[�8u�â>�Kր�:KĖח�Tޓ���G0��U`�J{"�;/E����~˰VXF�k����r�k�j��d-�U?�iлMӯ�cN�NȚ*�Jz�͛��>�wJ6^`;��C�߉U�O���s�]#�J�jBT�Ma�y�tw�S��O��+lR�'�փ�i��M�<����Tk�	�S����P��D�[�ǝ��q���>Fnٌ��4��\u=�)�"rR1�3mW��)�z6�P�O��z&�����;^W�)N)�+��=�Ѫ���pJ[sGH���(��E��\u�}���^mρ�A��l�Y�)d8׺�v��
��>%�jh�1V�hS��+<y�zT9��K��z��=Hj��l!��$Ǝ�L��9��U���@Q.A[O���w`���)�K�g�!�s��	q�S����/v�K�
��'��14�ϡSA3!O�P�΋��=�9��7�ڗɔY�����D4d'�~�e����|D6�D�c[W�t����:9�2���݋��M����pO���9ƾLQ�H��B����1�4�F�}x[�n�`����r��w�������������/�M�����?���_��[���^|�D�wH���t�L��\���<y�>��do���'Ϟv�]�^���t����6e�j`�<S�z~f���^�?;aQ�ﱸX�S`�u,>�\�yN��u����?�\�T%`���ʖ���Iլe�n!v�2j���cGٹ��R6]��L7%��N���);�|o-i�^��B
��ul5�/]��@��p�TS�wT��6ň��$8�l?�x�]S�5��S��u.c)4ʯ˧�OW����]��n��S�IwC����z���XY�Ԛ�]ah\U��M:]1�y��s���{̐|4�dڗ�
߈U]i�{�1����voU�x�4���M�ڦX���K�n#쉵��P�0rZe���s�5Q�QW���)P*�5�^��֋��W��|b�f��Rc�m��B])�s�c�!��H4�{��K���a������_�����W\�<����?��͐���9"�~FF��ߕiR�R�İG)���"c�I�+ulw���<�x��p^�@0#�P�jU�K�Ԅ�Z��05�k6L�S����{½��jP䲚ᣢ�ƫ��,�2`|1t~BfX�k7^Z|�9�J��@�>�����(�ˤ��4>nXB$K�����w)��Y����=b��=v�e�<��E��R�6��y�}v����>�wμ����G��f�*LԐ��E
%� �;���s��<��_P-nB�<~
�L���0�C��#����xo3���������#�����"�k/���(�jw��a��<��4C�2�Y!&�3�ἴrR$n�xu�`>ߥ����7?�����ٟ��g���'M�ϤBw���3�}�_����ڷ�~auy��
�����I�6ZFy�Z�|2��������?��ppȎ�վ����[��@�x��Hld"M`�'R�n��#T`,�X�/,X3A���9�k�X+�bZ�<_=�1��U뾄��^�L��;�JƂ+nf�h���R��&���Jk¬��ӿJ)�6���,xq~d�6R+0tT>U���O JB[�����r�.9���%������ے=*��S�'#6�w)��E߉(�Y��@�MID�4eq�j,D	��R1��Qk��6v^����_���2��\u�qCK�r�8���keD�\ρ�Q�盲W��uu�E#/�<��B�q5��|`J��+��9�	U�������Q�rI��^}�؊:�%��eH�yx��|�O��΄�n����ʻRi�gn���C�?n�l�{{���u�X��C�
�(C���؞���Sd�����_�G�"5��8��ˆ$��*�k)�����-�0����3[��n5ȓ�������EM�2�m}��Xp�R)E��`��]�ެ(�w�OUb��g=tb����b��ϫ:��=P�|�]ɻ^c�ד�P�"Cn�ؚ��ir�D�%��t�����y(r���9F՜�ڤ��mKK���'��Zܪ2Dt?�F*�R���у��]��ɵ�a�X]�/������3�s�*Obp![Ӧ�BX���w�1bu9KrKn6���\����
�N�:*���8�����`�&+��)�G�/�ҒԘ��+z���p�.�JZ^M�5.Cp���N�G*sJ�� X2V�@�g}>��z�}��\���-r����������o��;��>��ϬB���mN��������o�������o�޳z�uy',�)p҄E��~����~3��>78J9����D��0-'�i<0nX�~�*P�y�z7>Y�6Lpsj�&~�g�����HK����K��9S���O(�fC��J�����7P�J���[���K���y�l��χ�R��ĵ4[,-�%��M/�\��p��UF����Wą��'D�Jǹd��ÿ���p�[Y�ޠD��ÐA�>0ay�)g��~�7ޫ|)i�V�<K!����	�z�Σ�0T@�1W1�(R���fKruu4c��d3F��~�1Ql�x�\d
k�{%�J�kjʱ��'�LH0���J��b�k���iPq���yc�,����Oa��.
��G�X����n�'֝��܄�
��\�5=�bCO����:")z���iD���U/A%\a���,�5��B�VI�\��篺�feP/A3�)��
���"��0b��{�]�Z%1����;c�Dٗq��ثFa[hFL5OuI�j��G�`�R��@����ÐZ�Mv�F���ȇ���yP��}��Z��R�Q��I��uiO�R�1�jXA��v˻�������wHm޲Hy4 ��qks�3���(T��%��w��Ȅ��'�M�H.��?F�lCn{�\{�pJ�s��#��^������Pm5�Z���l���N��%��p�:�>\bƬ1R���.��.�~fwF=��k�����F�#���~�q���wV���1�`��5�%�!�i�rd��k̲ن>�%��4s<����܀3R�Nh�3����j�;c>���!9ך���C�����X����W�����/��
w���~��*t��K?���?��o��?���W��;o�+��F9�g��	�bv<�G�k]���d��?��.��/o�?�����ދu�-��a�v�C�ɹ�Յr��˦�D�41�&�Ni6i0�t�tx�pfL�Z�Y�O}L�6�J~������,v���[��, �F)/_a��e��!W<R4>�����=�c�ߍ%��"�+��ckL��,���M
�R
����$� t�`L�Y!����E��ezK�*�^�꺊�Qǆ���*$3_�y���YG`ͦ�UӞ+��?c�ǝ�|($o�~��TA��@#"�)�[����뿦0��@�!�7��+������M�?�S�U7[����lMK��ص��S��L�ci:v��*MnJ�6�Wj/c�HR��1��e��Q�����{H�Έ��.�Q5��c���]���BA��u���yj
�+�>�� n���eg^Ub�g�p_y`_��\�=Y�Y�����(���3WX��b���'�
���,���
�����ݖ������D���'��
107;S-���d�t��(�\h�jặ��j(� �������grU4�c���Ɵ�-ϱU�UN�P��!/�K0�R�R�!g���L���ڕM@���o�򵻳�l����}�c���΀�-3� 0�mÖ^ը��w�n����j+��,s��	0>K\�Q���r��������Ǜ1CU��4"Mys���c��77q8@h��!RpA-�W�??������A༙:�K�����"���6/NP�����xl�a�~�5��)x�#�J����k�r����O�������g�;w�?�
����?�������7��� �}�A��aq�j
�.�]=1j���f �>z�=��ķ�O�X�v>۲�-��ܞҩS�݈B��%�7>&i���7�>�[��p;��MS�ف})Bc���'7ӃG��}���2�������	��*2����k�x��ƿ"%ܳQ,*MK̺g��[�"ȅ�ֺ���1�.�5<ShH�)ǰ?�f�Q�h8'Q��ؾ��*�$��Z��QQm�'� 
�R�T�n�sO�t�VS�Qx���HU�E�wJ��_S"z9��x1pbZ.�Y%������V<]��)���b;�"�҆�>�R+��z׫��T��	��/H;��w��ڎ�w�Q�x I�M��B��;*�/
ɦ�+��YOa����FS[>ޛ������U�xx�Le�#��5�Ь��w���#�J�&=������̡Uc��"\�9b���Y��ϥ���2�J��x�2���T�դ�.R��}nV���!%)�c<����R�S~Hćm��J�Z(�-�*����kdH��ma�;gؼ����5`�7��Ho�����6�K�6���h���N9����j�{>�J&�沈��?��q�k{�ĠI�ݠk�1��n��ۃCs��T�*\��\��k��$��3¦��q-��o	z�ƽ'�=�5R�O�B����>O|�C���V.H��i���"���/Q�����@��SN�8��&s
�jc�3<m��#�;ȹLk3�(���0�`n��~�2?��h^�w8(�	1)0�x�N���BUN��2�����d}�����?�ϴw��L+t�_��_��׾q�7��o��j��e�d$^�Y,W�Bk�����77f�\���;�o��a�^]��?�h� >����נ9��,Qc�VS'��{!	,���6�>��s\H�㯡)`���a��'0��߽b��T�mc	[���b��!|�&=9=7]3p>4����v%�.ʍL���Ee�
(BS��X�N�ޛ� ���J���eE@ JB���q�TUSa�����A��w��D��=V�[v�=k�4O���B�%a-�^�[���O���oy��L��&*+^���XK�([/�}��jӌʋ튩I�;�3�W��߭��:G�lءJ��]ޤ���_��B?�6�'rC���[�VQהEU���<��m��g ܙ@��ʣ��u7#�y�/����0���yx�>O��]|��Z���P�J������hVB��ޢ1m�W�hHKh��^k<磎ߛ��H5/�5C'����"<�iX���I��E��wތ�����b�俄�4��}�aUz"�#�6�X�¹U�a����w����
(<y�0<ښi�:'����f�֛�h���'R��4T���+�M\3�1_`�'$c:+���m��G��l!������=Fi��ȫQn�G�k��d,kݺS~V��B �@�]��#I(lX`�Z91���I���c�.��	uޝ��$Х���>�T�$Nλ�s��+���&�me�G�|�x�:��r�,�|�W~�?<&�	��q�s7Ɲ6���x"�0t�f��>zuF�9SS���I�2Ѭ�URҴK�UҦ���p�F\W����ۛ��/��O��_��Mk�}��y����]��g���_|����}9]������&z$�/kABX8l���>J�|��'����~��X��!i(��������o�nE�	��X�ю�|�dJ���,�ʵU����\������I=t���#\�h�/����X|B�cX��Z��L���t�:�����������1�TC�[f�),"�LL=z/���l���r_�i�Έ����#�+wJ�D8W�v�(����
�0����P^��*����O�f��Ҽ�6�~I��
6�:<�yI���}�y���614:Y�^�'(�~�HA���q�*\y�!���8�,��f�/�����b�ŵ����TGA�)%ۯ���!M�sm����=���YS*��?`���o:�����q���}���C�L�˲IU%�k�q����;�;���8u��w{�f��`�f��9���^vw�j��w�C2p}7�4�L3M�iN�^��_�������Ci�c�L�{��؟1 {[�)fƣlGWa$����Z#��%^J�u��x
��q7��#FQ�͛��1���V�	�qe<;��a�Z�]!Q��)��2��6sg��ƞ������pw�����jKRy��M�U�Q?U��D���^�k���Y�ʢ+kΓ�|�'�i���fk�ro��cB|[g@��ᴆC�'�c� ������U�4���in��}�Gչ+������������8Hۣ���-�#�_�'k��	���T���;V�s���$�Y8*[�n����e+�]#��u��6f7��㧾��������o�g��ϼBw�~�'����/����ߛ�1�ϙ����	���%�-��B�m�3���'�U�n�HK�r,������,�2º�"MM���T@Syǚ,��M�H�����&���V�\*��'���p)�o�#��� ��ѳW�;�-<͔�TĻ�X�n A�e��
�!���ƟjS\a��VQHa$'�ZB�e=���K��3��չ���/�9�i#�Ŷ�\i+y�?d�w��:��͵��Faȳ�KW���N�d�=��(��ܨ�!�s��BKk�k�~鏦a�.�.�{�1|��z/jS���W)�^N�'@�0Fb��Ko��'G���P(fļ.٩���_�ZνPt�OE�T�ݎ����*��N�ٹ77Eh�~��t��tdw�����2�^ؒ��zJ���K��3����np�W�	���.o�?�kS��a0��f��@���s��~�KI�� �q�r�~��0l�;��<������7e��ٱ���'`�"�������r�am�l�&ی��U�V�d�V�tIL�C� ����%�(R*���!��Q�sP]��z�@�I�4-,ʛP
]��=mÝ�LG�	oS��u�(!����d��N�z�k��`�e�I�Ĉ7���CSv\��l�2�ݫm�~:C�	����]�C����h3��3(O����:��pJ�U<q��6�x�f��C�ᱟUL���],��d?�Q��s��F8Ff?�����U~��&2~v|2k�U*��`-��"���%~���+��k*x1��{W>�oc:�tw�?�����/o�T��?~,��7�f�w?����?�W�����b���,qb5x�sj�P�iuj\xoe�q�O���wC2E�Mq�M2aŭW�D��Ps���餌�.�Z��6 i�/��ݬ�!T�,���0Flv��1i���m�zv�c��R�*��@X_�h�lz6�X�d�5N�����q����
7;�Lk=�gQ�CO��r����{A�-Fm�P%�2\5]DG�>޽��\Ĕ0AO��W$J(�(����U��Ň�l�5�T��p=�SR�w+�Q���p�Az�7/�*�����uo.�N�W��M�)8ԍ$շRb�O��k�r�]!�|�(�:�0F)�p�%��c��mc�$�܋����|t���,j��(aAJ�F3�Pa�a�u�T���E��)��)i��=ϳMU��wj����7����_���<~���Ю7�jJ�>�Qs�a�TA�,���~MuG[!��Y�	�?�}���=֗���fˇZUe���:��E��5�5S;�V�(r���䞈���R�N��s���T�z�;4^P�S�l6\��!&�,����h�䖶p��Wna[��y�9�^4�m�l*�u�c�p�v"�ƌW;g��<���tO&''��M��Q9���	���u�|3�F��T/�����6(H��*n�����Q�g��̼nd�1ƀc�[��R�܊:Ȇ
�������!��`vGۡZ��mhQ�c�'�]�ru�6xuDM�#*�AC;A]2>��&���I�?�pU�L��G�����AxD�����Xf�����s�Ӽ&Ͷ"�S�5�k�k�7����7�'��?�������c����ʣ���W�����'a�6l��h�"f�J;��Ж�#�&�w�~L�3j�c�q�U�s`����X�C�]�x��>�?��u3)8�n,�]S)|��]y!!Qi��A����Wݗ���[+[�Z��(��V5C�/�h*�u��C��c[�}�^O�O��l�'��M�@k3^�'Wy�k���Mw3�Hq��|z�=���pE�˼��Jfh�]ԱW�3Ԡga�C�mh� 2oZ܁��� �r~�|\M�f��d����_7%d��2�RȎ�	��6}������r������xh^�*ɵEW6O/���0n˭F�7C<:�%�n��w��Q��W�Δ����^�P�����N���ma�vA���~m�Q�(�Va�}�>��y�|�OyDT��S��v�d~��|�|wSٲ��u}տ����>ꥶ|�j*x��gokC4\B�\`���U8��.��Q�eQ+a�ܵ���Uy����{gX�OȤ�{E�sOg�.���s��U��Q N�{j��vV9�":+�U`�Wt�$o?zk���S�����n���D7�a�Oek?s�F3R�KU�Hp5e˚���8fA�n�	Ii�$��ؔ�-##��&�����ŘlO�o#ǭj|��tX~.���-䩰��X�ѓ%o~��"E��<��N(�4�m���6S����v�px�k){-Aq�ݼ������_��V)�o��ʵ�cI~�hŔ���Zd`JNC���'36ν���I��s�D�9)���(�z�|oc����/��wz�f"?&�������o����~�����ˋwnV�޹4f"lEMW���5��9i,TZ�=����>�������3.b=JI#Sr�oP�VW� ���h�RR��*1���)ao�v|k�#-,3dC��I� ��U�"m���{Bv��l��'�'&QN�v�vF���	�����+(t!���Ҳ�P�׼��z閙m�,Bu&Z��4�b���	C!�
���L �|�[%.�hL �{�H�$D�b6]�+�ḑ�U��|��L��c���Ӑ:���QNR�j�S^�pg�@��=��S:SAy�ӌ�;U����{Wn�W�E�n�/��a��wA�U������|�3SA4O4�?�q_i�{f,EdHq<ø�m���S�'�\�
�9�!�����j�j��i���߮r=n�v��^ܿ�����������6wQc�Z���ƺ������r����PQ���T���Xb��c�]�"�C���u"ڕt�듼��>��"���xˌ�N��аrᇹiViL�S��TMus��%���yy�r�LmQ�k��e(������L����g�Iں�֠VN�+_�ى�����]lzW0��~�W*ƹ�.V�-N�]#���{BBb����+Q_����J�w���Рv��(m���Bd>R"_4�X>к�a-�m����:}�Mb7�1ϭ�~|98>�P�s� I��+_ŹB��O�(��� o|J�΋���1�q�Y}�6�if�S��>y_*�e�Ȥ���W�H�}���ү>�;�{���O�9��wl���S?����������7>���p�-9G�\YL��E�˶9�o��ׁZ���{ 1������b2��(u������6,��u<bL�`P<���J�Ϧ��=8R�?����Uij�'UG�'�F��M|��HDk��+6�)�Ó�p��V!��>�����!y��؈��6���o:�I�G��B���G�a�*�J�uEg�j���Hǰ�:Sg%��\q���^_K�:�+����jA�MIb�I%�7ևW��_e~C�@�z�U��veo\Zih
�6Z�Ǩ��t��r��o�����y{�<���|��j�q�ϡ6}���-~=����J��yD�K^����g�F=�p;���^�C ���Q�����-B��=~���x��-b�������Q{\���RA���j�S�=�P�Rq��(�;��n��:�{4D&��{���E���^co�yc��ۛGo"�WcX���wR^�g�an�5���� &�N��E��ȅ�36լ�/!w֪1\�̈́t�9/��%���m�[��5�א_��E�S.���8S�ݕ�X���N��BM�")X#�Ex�bhF�8���L�d����9�Y�"
U�ڶ��r	� o8�>��N�^��F� ���:��Sw�Ea�@7����j즙Eb0|��vL5��3J�η��46b>7`��SCx��9X�	�YB�\�	����m7���Ջ�e�\�F)_: 䥱r� �>�NZ��ܽ�%/��v��`��N��������ڿ��?� ,��Ǐ�B��ݥ���w~�7���_�-_a�>a�-.��hU�#��P�x«+ہ��}答|��ǃ+��+���4��EuB��	����>��Ǵ2n�Nz���"�ASU;����7W
���(�V�#��Ek�dc[>C@⼒`V�L��8�,y�/[���TN�C_��"��/ƽϨ�d[�1�E�1�4bqi2�!1�K[R2S���~͘B���m�d�ϔ��8D�P�aӉ��卤C�<+0�ݮW�g�������"2��2�1���F��m�п^�FJ+ʾ��6��A�vϻ��?����Ymy��P�*��
��J��X!'���~�"���������f�FН���h
"P<F!�mp�TQ�2�j>+&}''�l���?�G)���S|输�	n���� o������Ow�$�ko���Y��z�5��H��}0��9�'^i�I���S��ܙ�]��|�
��:x)��̴�Ii�,�R��Ԑ+#O4)��)?�dp��FZJ��*�t�;��2υ�-��J�M�[�=$7{����[��BU����f�f��B�R!;o�MG﹗�[}��yja�DO8�O�J��o! F�.&1<��[e�,$�9O�cNf���d��{-^���=�
�s�#��Z�]a�m����1�?�����x������6A�����Y�m	#�qQ]S42E�<�iU�T�������vk���_���6L�"0�ϫ�	�_]i@�xV#�N�Q>��8qv�����|ez�{��+��ï~a�ٟ�!?�o�X)tg�g�����������W?�����fy}pF�5�/M�Xh�w0���7�V>��{H��1�����Kb,s;�A(�O.Z�� WW���,5*�Ĕ���M�)rQj��X�
s��ON��b��@�R�V�a���7E P�zG��������ḹ��ͦ���<��������4�[�t�5�`��E�b���� *X��iz�++��Oa��]#��][V.0w-v�I�p7�Q �M�oP�;���0|eiP�9���b�4�*�!$Lgz�,S��+~.Z���7^[��
b4���4ڐ�{F��� ]���Oᐊy��Є{�Kp(ŵ��� ��)��W���]�J�)�n==�p����P�J[���(�"��*.�Ɋ���}'43-r�Zp�ϼo�S޾-1������x�Hv��l������Z�9��P��))+�y�1H:���m���Oej6���R�S���~
ٺ���xs݈h��
MRTO���*t���Jq���"��RO�AI�����hH�
��r]�\��|�1u?��NSpJ��:^+Fy�ss~_����&��1�#޷�T詺f��gEĽ6tg���Ia!�{��kux,���=xj8{Iv�ӸV�9�9��P�+wJ��J�zm|�nƐ�I!,�(�L� _YUƪ5�S��t\f[cxLx᏷��w�l��FF2eLX���y�T)�ztD�s�
��6����/�+d"i$���ZO��p��u�ρ�/	[^�b�+�����O(�y��n���L!pf
]a��%X�d��2�Iӽ�z�q�o&Ͼ�;�[�+����i��c���S�?��;�}�������wz}����w,� [v�D�$EV6�����Qn�*�`�MQ؇��3-tJ���3Z��9���3;�q��;X�<`�����"U�l�u q���N��gU%!�V|��k"����ٔ
-O�e��.F��uJ;
���%���~�P0�[~v������%��;�7_T��ROF���bQdJ�+fk��D(+8h�g����Xn������r�x꺒C�zK
_OE)�a�٨��+���c�/���c3�U>�G ��:�î�S�3U^�z��8��>�M1���i�Yg��ʬ�Oԁy�����U0�4gS݃��S��������7�1���쏊�����'�D�_W�������D��f�E��f0�qs���Nbp�r���Za�׵�|�G��}bͼv.�Tm�<T^�1�s�Z��10�Sa�g���������o;�E��70�\3F<ZW��?݇�wH�'*c.�&Rڹ�|�	�����,TH�|��xi��Ę�hd���+�غ�>{L��^F���T�zm��Q`���t�S�>a�⪖���&�'�!H���1�^һ��J�hޔ�3*��T\���uPb�ϨH!�qm���kl'O��n�&'��F*�(�]b�v���[ �H��O@4��y�6�}|r�����0'nLv���
��P+I{�>���DV_�#}vFH��☸9�2�P�ƍ��%�%7��|�{AN�2�q��䬃ܐ�|5?[�>�����o�7~���Ol��?�����w6������o~���R�tw}�����*ȍ��&(����:�i���w�Y<���8�1�k��1���1�(
�z�vL�e99ۡSv\�Bte�I�X��3�dA|j���+6ℿ�c�h1�Ũ�h2,^����Q�66�8(����P��c�;� 7X�%�U����8c61}�o�
R0�bn�R5mJ�`���;Q��N�q%7����׶!Jܭ����� �Z�ij�=|��㗉�<�(x{k�[T2�B��:�x���+;���"7m�J��,S��J�@�zܤ���*z9�ou���Ek(XȢ�J�`�`|r/K`��"MY�Î���ޙ������ᗊ@d��oO����!bj܃�����?@gQg������' ���
2���� ����0_��;����e�յ�֐J$k�/�3���ۜ��5�T�7��(�.�L�1�հ�a�>���bmp���Ӯ!��l�4?iF���T5�+m�s�Jʯ"STl*�dHh4����E ��zo[�*�|ۗ�1�	/���Ǒ4�����<Uwf������iː�Y3Z*������Ag��ޙ�{f;�Lq?��͐ynQM��K�R���Q*=�y�$ܒu<ak�o���K~�mO����q1�S2d�/�r�B>%�F-�~��۶�9Wn��b
K�R�+���iۮڦ08kK0�� ����]?�<l!��K��5h���R�+���Z�x�t=��@�o&��ɇ[���ǯ��O�Gl����?�
��;˓����7>���8�<���l�+7XY�m�2'�s�t������`og���lJ�Ǉ�{�dZ��i�!�]��fJ����3X�~@U��ĮIc�3�RQ������]�9�`�W�u4'�Mk�57�$�Ma��hzT���@ïz���5뤑��b�Aj>���ƽ$���3,f~�J�_s�Y��4�0F�B`��y��f��斁�V5תBS���U}s�c�Tm��U��Ч�7O�R���l
��ǔq=E^�;����vr����� R8^RTBk$�?�!9�q�TJ���^��&�3�A	��|#���U�*9̀o
��^J��UX�6�M�M����s(��y��3<�xgAL��#DBR�K�#>�nI݇�]#����������3?L1���'���]��P����N���V��ߵ.��_Cn|�{D	��Z~��^�$����u�WTQ��}N{_f���q��\W�z�)J�.���АՈO�=F��q�io?�t�������K-z�cUS}���Qֻ[�x�R�}�>�i���>��!�\���?��H���]E4�"o|pl���/S��a��JԂМ����r�	ѱH� �[�z6x��l�`���D��	f��4x,��3���Z_��spJ�d˘�*?�0��:V2�����A,����	���T�*szC��_�ƋW�[+�(S�,i��_��W7��.2��|�jVNdV���l}�)߳{�i�f]��Z�<��׾���[�����;w��X*t��_}�ݟ����O�~�kĘ��X����
���0Ʋ;�+���z����	��_P�����W�ԗ�����)�Q)_�_=?om-���Ϯi2��;�����7JD(P6j��,��¨�&6�^���LA�:����ղ��3�{�σ$���D��19C��r��������Q�A2�v��K!aE)��]�I�l�M3.���i.�Z	��1�T�H��Q�vT�&���^R��sI�����tAa$���.�a�n(�����f��qHSO)!��(��]��-�������z�z�O�)�R�M���Ac�*�}y ��]�:�UrS��u�u]���aS@��u�!�t�ڍ��������:r�CodSwe��o�X���e�;�eT�/v�?�ր��!��ģ������]�u z*�����9#5r 0��DR$E*�{<���,'ٲl�
c��%[�$�([b� $�s����˩r�U��ϭW��@$�]�Qx�Uݺ��sv\{mU�z-���W9���v~t|�6�N��ۭL�k��z�=����ݼ8����R(!.5�����dz�T����:#S6�-�[�l���ƴ��(����q�Q,�h�<�&G���?]�ǹ���3�/�2;����{�`�1%�C��)+�1���A�=W�ogW1��h��i̗��r��HS`4V`����At=#hɮ�K8�@Ȳ/�cpQJ&8(n���1��i�^�)T�$ZO�s=	eN�ɺn��ٱ^8�0�(k#)� p%���/i�8d'�d�2�Nc�����B�58.����-����p�y�0�t}$�B0=#����5Z�͕S�#�SX�Z*��$��P�jF$�:�K�z#�o��w�uʏ���X���'�~o��������M��
�(e�X�����aFHw��J��(&N�l�7�<Βv���� �'�IL_t*�!�]/���pe���:u�J_36�9JpIɩ�}�sa��Wb�&vG��o��&�8O�� g�ޭ�J�z��Q��$����n���e#r���ਬ�c#Z7L"A�SPŚ����1$_�,� ,fZ�!�"9�5����ִ��U�8Ϋť��@�@)]C+C��$�ߜ	��H��ѳgͻ(E��j�]�z�1��=��*���!�D���g�P,u���ZJu$Gϼ-}{6��P�p����g�o�� @�
�S6v!kY��:�����g-�R-�]��S��y�ʅ�
����ȉ��+�i
^�m��~_H�x�ӽ�������{�Ro��
��>��� !*zX�9�v�6���z�z3�Q�����Ι�!��)�f��Z���~��9�2��P#c�	�͆���&H��.wV!{e�����!�����{2��r�3Z$r�����1���e9;o�{S���$�a��*�����4"i�*nDs`���_�F/1,�)lH�血s�J���Ajj�͕��s�֪l�B#�`T��Qikԏ�Wr����O'�P�h��j���H."�ux�g�tF�"5���%(t6R�.�#�E�,?Jf���$��3Cʱ�����eN�Y���������oב�CG'�j4���Ĉ�{$��(�k`��@�SY�ä�Y����7	j_���]
9���u�g޻9��;w{�*t�Ƶ����=�����n�A}984�[ܱ ���S�`���7C�	p3�S6s���Xw�u2�-«�_:b=�|a�`��k�s���}g�Ӆ�K-gkyx��GKeT%�۴���r }�نTX�$%I��a:��Exy��((��JS&5 �d"�q\2��[ '�e��^&=\�U����#��0z�8$ő�J\�3j�H�Dz��C2����Р!D���?(}��g#�s.~���4ol����F,B�ݠ��S�<�b�Ӣ<�'"����ē���B�iK�B(9�@o��U�:ah�ۂ�T!�KC�O�7 �W������$B4NW�EØ�m�_����|.�Z���!�r����_U�u
����g���T�޽y�K8�u����W��k��M��-��_%O`�7sWܑ�4����]Ne�D�V���w=�M��PR CQYy�p=z�vʞ��f�Bg-%�����!M�[�=���ie|�J��-��Z�#� �Ucp�r�S#"�i^�u��Kx�ǵ�(���¹�y\�11��b��*Pňh�UF�lچ����\e�KD@�:.�)��{`2n����8�z���@d��BM�s�ax��Rʽ"Z!ppy@ޤ�C������+��b�T��݋4��Tp숖�As��!#˨8*K��
'�!��|��U���T9i�Y!�}� �.X��NG��|�}�������|p�f\J�d>�T|9s�����u��� �B0�Q#i,��iG�g���ҙi����������n�z�E�����7GC�/=?�Ҿ�/?7_�n@����*B
��ǤJ��8q�n�Pk�w B	�ؠ�ٙ�P�w���F>(�7��;�Ʊ=���Kw<�|i2���^O�����%�� y��&,�&¯(�p<��S �T:�����[�@k[ĺ@1Ÿ��=Z��2����Hc������*�;i`�FU�B����!3vNcs��|$�!P��#k�sM������Z�XY�H�(A�E*r��HxV�	�Mi$a9� >�h^�OsujM�[���V�k3�7��dO*HH�w�O�(p�HQ�FO]%Ų�cH�:H��P�Op��#.��ܚ�^;�S�+�ͽ{�dO�{?�Lˈ �j�TD<i:C�E�
�w!	+����zo��V�Ö��ç�_�Wx�^���Es��Ȑ�/[L�v��U���'�D����E�F��ӎ�gU˟:61Ƙ �4��5� L=6C�K�(�����[2��h����qs�	�$�����b���e:�)!���`J�~ԆSO�k�
�^�jy�������IЫ�9x?T�b�Q*B�#�9ׇF�y��t	���E �V�{��l��s���89+�V�S�9�e��f�a 3������d���H����maȆ0@�-V�?�	Wt��J�o�����a�ɹp�*��^����X��PK^�1��`y0�rk�F �B�u��w��B�Jw ?r������y�s?q�}�]k��C{^��g5�]�U�٪�n ���
�R�O��Xtj�"�XJ�E�����G��[�Ń���lY�­�18�����9�W�MN�ZS�sǡ얹f�՚�C��!���M��2��-�CI�{���*��� �M��EΆ���Ζm�TĔ��X2�m�K{���
�������o����,F>[1�uy���0-�&2�A��b�#�-�>CbP�`;rx���qB��3%��*��КQ���Č!-.Z�ͱp�3�!@�J]�lxNe)u�����R�D�p����؏?�_�s�z�9��sR:�NˎqO��'!�Ζ˲�'��]f��M|�Ч-4#�UH�K�g=#~ȥ�vC"۝ �ԅ!9,J�H�9`p���Q	A�A4��t��eύ�S�NO�/m>C���[�N��ZE���

�zN���9=)-����L�$1),����,��oO#�u��7?TI�Ј��kD��	Aな:�x�5dU_H�ӑ2��ZS��N�Z�Rp�n퐼h1�q5�lhTp2fJвº�Ɓ���0������q��%��3���ˠC���9��z⡉�2��B�wm��Ծ j0x����}V�%OV5�H�J�9V�o��V����������Cl�O�x�*�(N� P�����S��2l,�D#�ah��	8�� ��|\O��x�tq�c��ZHpp]���R�S	b�:�Iߞ���� ��<G@�{�q��!�0���l��=dh�%!�z�8��ˮ��١M��܁E8=��!�^�G�:y�p���I1[��-º��ׁӕj�s��0��C��A�V\��T�D��� 
or�ٱj��7Y�[�1r�����j�-�Zs�x�MC���Oo:��'T�����}'G>�H�l��pR8�D�+[$�c��*HG�\��.� �D���r�E��`��T�{���+�N���~����W�[zB�o=u���Gw<h��Љg���Y�H0&u�-��J��B	�����z��vg	!��`�C�����������w����K��/W���C���Gѡ-���F�0J,�w�pV���(.s��o
����N
��͡I�
&��BP���ݡ�BHe���"
��i$J@t�91�S.e�5`pH��\@>�(h\?����� �V8�Ar6R)� �`�&��}�=�Tay�9;�	��F䔦L�ң���~_5�F�[������r�=B�K!�j��w葲���V�f�z$�w"���)��$�/�C�˰^��]�+��|�Q�ݘJ���*dBgE1R1�	��ޕ���;�!G�[Q�֋���ګ��	a�y[/=�a �UO��A����&z@�U���Ku�)�:��6�:n�_rj1��Q�s��ƹ�1=��n9<�l����-ߵ
������a���d(_ �*Z ˭Yc��[�K�̞���T<u��q�42$��L�K�����?�n�)Ɩ=7烔������Q
QV�0����Q���Y�DF"64,��e�,!db��\�\���&(�ŹcG��g�����l�J� �Lt$~�͑����z�(�+m�Q^�hFH��`��b��<�Tń��.H�I�<�� C�dH�7���c*ň��:���!S.������>�X#(5��C���$[5���ր!�8 ������;�[�?�������gW����:��W��f��׉d$MG�GB��|�&'�W�K��^C�/K� �Z��bǗ���k�����k{�ѹsO4��:o�c��N<vr_�:lp!��!l�Hm��;X�@�2Je�$�E��B?,�By�b"_�Nb.��j>�[�����[��?��/ʐ��?�Ǝ����|ta1[�蚞���t_��BO�~xְ�� ��Q���b�!z��k������JO�zE�f*m�s�����(�\���(2�����бB�g�8ٟ%!���	ǂ�Yω�+أ]����5�ȷW���P�<�7�� xER	EJ$Y'�W�Cz;����
���2amΰ�
]
5�����6(I���)�r�i���Щ�����R�G�"Ο�uQ@�#�t���C���g��U�\������	=H��������RˋiU q���}ϳ���r��Q�vt@F[/D�f�;z�+��؋.b�B��� �JL��r0�"�1����|=���B!��sk�P{,�ꑊ�5�k�sZ�YQ��f@#��ِk�Ѹ�T4hu��%�yd?z��(�<{�_�]74����#�O�؇Ƿ�_~0]��x.�ǰ;�-�����U��8S]�\ȖU����*:�������F-��{C�B-Zϝ����7"�q��L'�T�ħ�p%~F�"������]���c�SC�vzD��a�$j��@�#o-%g���J�bp^�N3�HJ�
@nY�7���s״���Xꆨ#$k�lH��!�^)�������P���y4�b��bOd���z�%���p���/tF}��8��ӡލ�%�L#N;Pr��۵$�z�-x�~V�Hd�p?���.A������/}��ν�wN(�M}��W��޳��O�U8��q����Z�+�EYB�<��-�ILj�����CӀ�Delސ	��&�6�$�W0�����̉O��7~����+���W�q��ꉅ��S?��E�������IP��䂜��`!��E�p�F���V �)J�G��lz椤l��DB�4�U���=�&Y��S64֮[@=�(�U!�HA_j�E(�[�xC0��2��$B@���o^=As8vH��U��
$���R��OYx�%�%sTd|y�m.�{`<����4V,�������
����H��$�ݡyD����yMf�Е��
n
Q��9�bT�:���
-����|"DBK>]�ja=�'�Y&0����t���eOP:e4k�����Yc��P���,��{UE��{J]����y��:��"�{i�FS��5l�Ⓗ���1���`ʥ}DU��@�g�&��F��+1'zM� �5p\������ẽ�2x���1�
W��4ݱl0YQ�fb�x-�^1ږ��N��;����z����3��<�@!N-�SI!���֒U���r�Kĸx�����b��jO8f������la)�#p��i�Pf`�"H72z����m��0�%�#mkP�Vl�,�2mMEΨA�NA���y���]�5���gK7(K��*���Xhw9��a�@kE����@LcZK!7�R"��O~l��~����f�}Or����W��k��N*�29=���ι�	�F���b,Y� `M���k�F^� J��;_tG��ڡg�_.wN�w���B�غ�o�ͣ�=�R�f��F�����-c2\�G�'d^��;�gb f`�.�J�I�<'�B~�
�t_l|ӳ/N��K��9��_���}��+�����◿����R*��ڊ?����h8����"�O�ii�ȅ�MH����a7�lx=\����@-�1���<�?�s�B�/� �M%lÖa���k�K3�.@>���g@�u ��ȿ�Im�\��2�Ϙ�� ,��I�͂z�l�BR�G8�v{��9�xA"\�,�G���X+��a
���ٰD���&.��tUJjn�����pL�M���7��T���J}AL{'ޞ��x@riˠ� ����(1����BȆ�=�"�����󵚠��<5$��b��y�O�� Za�P��Qf��*�<�z��'�ENW���[�E�
�����'K�Y�²���ݷ��5\�q������q��<`b�x�BXd��w)^��f�W޻Z/\.��f�v��Ўn�@P] I���ry��S9���7r��z��OxN�5��3��dJ�J`'���|T�0�C�
�S����F)��i.��- u��� ����©�My�<�A�G�����U)Aõ�y���	�e�7��u�5��+��2�_FE��K$�b�����]��B���R�HI�����=�I��Ĝ�Oß؈�h�Xc����L��?��k��K?��D�L��w��x|��9��mU�4�7$��.U*b�(��V2�(��6�J���~+����V�u|u�����E�2����w���B�t$�޾�xp׾g�,�r���ں���t Z�?�D�a�_�Di9�\z/����B�',qRI���@�WJ_�����������ك�����o�f��ރՇ��?����3�O��C��=i'��z�Y$�y�|j	�P��D(�.W�[:�1�Ć/S��&�E%��Z9Kd��hM*�7��%��������r]�̍GXg���I	DQ-+ʧ��{%O�K�h
�1g/��D޳0#�p:Q`���P�0\OEG��I�Kx^�mH�a4����ߞ�M�x���	��D!�7Z˭t#x�㣎��Ɨ=DC�m�_v�9$$��l�R�jh�^w�1��t�`���̊l�ϼ�*>��5���i]�|�w��۵��Lm�%#�iO�J��#���7m�r[��s�����Q�獍�;�zSQr�Lt�I���>;M	�&�ݿ�
��X�WǍ�6�6�p^l1{(�Rt+]yM)�vgְQ#N��B�e�ɵ����N��5jBr"16T׋�]�ư�f�%������h\�m�������Au�4�4�����~�R����4d���j M4-� ��ZǡX��0�(K������;�R)�3��p�2�F��(�_q��yؙ�v̪[RF��)qu997�#G�T��J���y����Vr�әa��U@
���&�",	\Fh�H�p�.]���|��ݷݼR�����������@ꂫ��ty}�7d9��yn�|���?w�s% �ݜ8O�K��4C��0Nŗs�g.�ֳ�}3�ş3�9���D6���l[���K/�]�9�u��t�dD�rd��&�>w��E�&
��~X} l�0u1QMk�eV~d�����<�S����y����V䶍a@)�K�������r���_4��e`=�H��!K�E͠$���
�3�y�&�#��a�2��wqnkgW �0YY�!qU���C_T��T�����BIE�PY�e����F".l�Ce��G�%/"�xE�
���+F��J�ކ"������ils�hPG�z�T��L�=LH� }rG��Ø�
��O�1��Guj&�Qu��_������s/��:��@�,�M���<�;u'����0.�.ay��3.��K�h�K�1���<U�D�fs������(E˳�d�UT��3B��t��j�TQ� ������/���UǸJʅ���E	d��=h�H��ͮ
U��Dy��K�����b�NH�t���^�������i��;����3T���HZ �	J\�V�O�f� m��(<��gC���#��v�"O:(����rF�7���eSqvF�h<v-A���f�I1`�I!�19;�qM�W�$5�N��b�Q�����C��`#Ԭ@�k�k�-E��d8[!���[th�L�Ie�*`-K�$(s�yr���"u�J>ȇ
�y�"e`��a�D�2���A{�����W���ٗ3�����¯}���ۺ*�[���<�g.��~��N,�?o�@!aW��ֲ�x_;�%�.�(Dg��<4zl	`,̜=*v&7}������.\�<���9��/�����=��ٿ�Zl(d�aIZ�l?H�g���2��� ����֟�!G�3Ӌ ����`Ҡ���&�^�W�)�r�w�>v����}��}+P�7]2p��c��7��������9򮦛ZW*�`8���D˞��
�K�@�P&� >@�1|�B3��u�da�aԑ���6�V-S.\*�׶
O5�����D%L6(��E��Vk���c�;��}z���i�C���B��c� ��f���h=��E&�0��N_�2(����#\[�� � HTr23$��]�W�N��D��;�|��yߪ�Ux[/�z���T���?�PQ�����E�[e��*W	�z��J�n�y�_=��\�M	��Ǳ��N�O�.<���U��
#�Cڈ2a�ԖJd�ޞ�n����/��!}�m0X#��±Ɓ�ջ.��E�|���g�tF��,�xMa-	��uK,#�vh��T}��j��y��6�z�r�㤵6T��ʝb�c�s	G����Q���5�t��A���q��,�iz���Ʋ��k��Ǖ�<0�s�r�%}���:�Ԗ�1�1�"��4:	ph,�xV,ہ2��A�G�$@��:����!�v�9a�e�tN��I~DU"+밭-F� 2k�zF��o��(�����D�{/�#e$�c�DU4�H<�T�U�(�]�u��D:ӥ܄�Ë���\�0�o=�4g"����zvfߪ��?������l��DT�L��֞��O�>I��oE2�&���^^ 
͒��0$�#�?ud�.@���Aa�`���W���[����o��K9��sJ���\��ojt0���|��pp`���.;qaF��/��%L<��*C�1(�r�=`��I��u����D�Y�9������>��o}��8���g��k"�'f�ϯ�����]�����d�dY:�� �P.�ϮFu֍�c����yc��BX��ZU	B��.�UI5f�J<+���rm��R)����p�UQ��Uqn�����r�֔(p�S4����{g5�^�8�)��땺Q.)X�.s���Zk(c	�ū�?
)��!�����'eql�"�s�&|���\}��׾�M>/�H�n8k�%e�2�nX�%{E��t��;<8Q�֣~�6�� ޙ

J�v��S��RX�Đ��/�޾ �E��(t�_w^�VǱ�Ǳ^�}����w:v=���&I��m�˯�z�S18:t�������k��j�G�5Z���x�v�8u���/���ʟ��i�.�(�+��W�δ��h�]�N{�����F���x�z���Eɜ��zu�gF�سA��^��iՀ*n�.F*Rg��P�nlR_N%�}�#��;y�-�ř#�	{-��:��!�')��{렴L�>f��0�'�X'N�ϐ�5.X�����p�a��1�?���FM�t����p�$��'Y��.lP�ܟ�(5�#<�6Kt	��	0%@���#F��5�h��ϝ4�#�_�}�o?��v����+���sy�ᙞ_��o������2Ԟ �+��`����M�H��/�>c�K��i��y���p(�`�l�TOz��k�^��g�{��v�)��Fõ?������L���"�#�����r�K���9��x	a�0¾,I!G3��bEh�H�*�-� �]e��R�h������-߽��oY���ͪ�0��{�~���׿�ء�/�\40x}<:�&_-���vOE����&��j��%(E���EZ ���%T�u�!)$Y�����X,M��r.t��lF�:K� (�D�Y���cN�sC=Cn^�XC�fq�2H+e]:4��:�X<C|�XS$F���3��"dXA>���ؾ�E/��*7�F�k ҽf7'�W��F�}�+�.X�袚:��'l����f��1j���i��K��"�&�S�@����ˆj帞2�.2��+�֢���IoM���ݫBױ�T��j��(���HI t�W� 8����p+�����I�۱uz�b��Ih��%���9f�r���}$,�:��r��z�
d��^��_q��pO߬!�Յ�c���3Ǜ���TH���@z��{���j~.,bċ�A�kKG��92�%��Փ��*o"�9�|~(�� &<���HSN\���hz�%���y�or��X7���0�!�@6�)a�k�ƹ^����"��K#em�^
 U�<�_q#�'`u��i�A N�|N�;���*`�a^��
�bm�};аt<���ټ��ŵ1
��Q��ś�F���@h��w߼�k���_�!��ʇ������\,����ɔ�L<SqT�|F"�<�&�ᚓgd+���T
5v��,:��s�����F�*=�sN��	]�}h�':2[�Ɖ6�X�$�
��*K ��Y#�2�"9ɑc�B���hP4yx�U�=C��{Q���������ũ|���ĩ^3�+Ǧ�?z*���L���Ա����NߖZ�I7`0�(H�bm$I^У�C��X�nj ���6���2�E�KF
'w�^����!�X�L�Q`j��#6���cڢ`ӞǺ0إ���<�Nx,rz�샱�C	v��I�XK��G�YzI�:B��Y�u�B�]a����!D��P�=&Y��(L������^�� �q�JɥHt�ǅ���'���''�
�c�fJb;�+9
��5+��9!YOP�L�*:�2�K4�
epw�;��-�������������I��� ��hV_KB���՛3������<r��m��F^q��s���i!L4�"lZ��OX(��������ջ���}T\	������2�?��L�/eC���@�.��p`�v]���Va�X h�*g���*����yl��H�U��F1�)0�_��cgڍ
X�&�'̷1zes�:e�(�(���用0�*�E�V�'�C���ih�.gjV�0�Ra�\�[MLpmI�Lj��ޕ�=x�'vh#'�+�U��Տ��*��`� %���F�40��kFLo,�
�r3������~����.8�q(���;�����囪���f8�i2��u��8�L�1�B0�[��5A�.��j:�R�q��G[:��W���u�Z���9��o^�W����1���su�4�E�Ɓ���1$,JLN�+@=�o��@�jL���|o�5�h�Y Yr!�*v��ε�<S��o���C��_�<���8�Zsವc�w��o�������x��\TE��D�T\���ǒ`���U�*��Hw5,(��j`bbm=�����3��g+�R�Ed�,z�[n{T*̴��N{z^�Wq5����m.|�lw�8�lX�"����)��向ґиz�T6�Ìo��t�4��L�i��i`���C�3` �d�މ�g(��rvE�ܹ*\v�R�	/��
Ԣ��n�M+R>(wO#�Cjs_�(�(�h H�As���q��u��
_�E@\Njب�(E��g�1SD-��j`����uoO�������:@n+��#�Q�2�^ߊд���c{�E{o�޴�� ������U�i�����h�i�@��x�|f��݃^��I�s���R�Lf�����K�V�yQ�rǬ��2��4��W +?؃��㌈��&�U=yQ�H!�^8&��N�W�gڌ�S�8���I�$=h����vq�����(�HQ�ޙr��τ4�+��Ri�0�Ζ���ŐժBB��`�2�;#gڹ�����4$���0���p�ʙk��>K�SV��m'`_�&�g�o���%��=֬N<�}k����{?y���?�X��:������������G����D�7̚a��7Oɱ#�Mo]�V���1��f0DPFR�����S}h���'>{��9Sw~���
�7y����;^�������dfd`�R�E�c�X;&�O�`-�3ǂȚ�X�1��7j�*,��/!���I�1�~z�&f>�;w<��Dyq�*t2x��~rՑ���~`ߞg_<��s��`zpc�X�%}@�b��Z�` �s5@xS�eZ�Sԭ��� A�O(X?���� ��µL�,&<�_<t;-~]͟ʣN2OP�r�2e��&Bg�p�mi�Z�"�	�ḑ"����	�:�v�p��\}<&+�1R��"2�� ��Y� �1tX��Dѳ$��9s�xZ���­� ��=�`aG@{��0�/m3)���Q�nw<8΃g(^�(~
F�b�Chl78� ��4��4VCI�W�OToU�y�5��G��GVy#�(��7��JS�O똶Ba��t��j�tL:����/��&i�q�]c{w|Q|?	A+>C��6;/ŋl���\�>�N��\��$���k�gV��[+I��-��A���%�N�0��{f8�ר��G��O�k?��L���Y�u{�V���,A�a�y�ia�za��� �OL
�4ѭ5�J��aY_���f�8��%`�1n�v�+����tՓ(���uI���6?.�Lux�b����iL���	�M}�`��?���{4b|- �Z���]���#R���DF�[����҈��>�������z:�,���7���'?p�ɫ�E-��kO§^<5��s�>�k�]�O��dDE���s�+�똈u5~��@/�Ɵ���!Q?��4X�4�l�ƙ�]���Y�~������/�sף���F��!�Na�#���.A@Z�")����"�#�/�q����02G�k��3R"�dO�inx��ß~���1&�<x���ٗO��<���w�:9U6Fz6�*�H���U�����˛� ����} ��Հ��B�HC�������k�	 �G��$l��H�rOG�ҩ��P�-������䭇�ܜt�B%h����:��B� ��H];N%�y��X�FB	���%7;� 6H&@8�0�x6�oe<��f��C�A����gj�Hi�`� ��b��F���=p� ���<��$���~:�=���*����)e��]�bi.��Ԝ�����2{��r��$İ<��K]�&;������F{E�AO������E�tl"�� >�AC��q%�W�9�)t$Y����"��Ǒ�;T��a�̂���ii	�:nu�#�̲1������ ���p�Đ�y�
�s�
���b����~Yv�u-�8T�bS(�<��t=(m�4���3�dC�>�֗�,&(���{�y�?�o1��%�a�q��M��G.����F$�n)^gY-�n���q��/qX�r86�Ñ�����E����4Έ��Uc� .
~��a�������#�@\)?atp�*D��r��|1)sL�����/�'�~��߿q����S�5���w<1��H���a��i�������-ܔ�f�I��/�?�����K4�s!��^3z�sW���޹��3�w�^�m���}����ͱ̚�r�����n���\��B
/^[L	ַ  ��{B�Y�����0�+�Q�N��P��^�7~�B�nC�ܘ_�k�W����O�.5>>Wv��wb�>���Q��ʢS��UX�MP��&�6�,4�Dd�
��B�A�N���,CS���̷��E<T��p.�[m~��'Ka�u�� zC�"��P���;)yѸy�O;��!��m
���T�d�����
4S�c����\��H3Ҫ���ɜ�
�/ޣ X�l�'�=�va�� f)���������
W�i
�P�R�ƀ�].m%O�L�f1{�<���D%�Q��B[��$�i�|�+\��u���i,?����:�/�I����N���%a�e�L����}5�t�19<����8�0X>�g(,�����x����_zÜ�L},J�w�Q�0Z#^���\�T{7Ѿ*�c\4:9��rIy
�^��Veܰ?���#p'^��(8j�	J�G)���oV|	�q�(�.d�D�=z���hJ�"d/�9gI���r�?0�ZV'���m�R�'
\##^����.�Á=���J[��t8WBV���7� ��Z����rHy����W؇�Ҡg��焔%B�M�0�<�T��%�V��^H8��@�m�h�_�����5s�;);>�����w�vS+�~�J�aC҉�a�y~	<��9'�m�:C��+)��9]�Z�۫U�'�Pw~ӕ[O��3��w�~�B��D��_{��#�;|o"�f|r���w��L��M<Z�L�*V��j����dH�H)�&1� :?�TY�Q]!�vp�Gncp��O��?��Ǐ��_�~�L��g߿e⎇����]{��>�=4_n�Zm9�N����&`��L��˾�H^�2$��2ó�l��BNu�<a&lOvr���\�o<���^����$c���	v�=J�CCv�l�D�Gü7�)It�,ōx1�-��xdP49[:2JB"
�O�뱱i9���K8�s^��Ue�V�	�SP�h� )���B��z�u3)8
q��&���V�����*Q�PY�d=`	�C�@Щ!��ן�%G/�I�
Z�����iz5t�j���$�-{�*��d�P�Bn��kǧs>Jx�c�X{
޶�~|�͹{��4 D�zF��$�W���Iu s�|���T9��?U�2�����g��CCD��PcR=T��5El�8���]AE2@�I����Hm���x)(�	o�%�i�"m���9D)�9�ES��`����6�W:o^���s��ԂB�k��9�����kA�r\c�!c����E��L���\�;A
�����̹��|�8>�&�U�BX�Ne��
�\��-x�1�у�"�x͜���E�)a���e�F�2�dOăŇS��7o�u����k��~��WL���7�ڽ��t��N�@�  �M ,����^4�J �Z�#MYD����8�8D��~@f\���e��}U��_�~ �s{;�:ݿ��'?��w=x";}cu��;q'�v�:P�T|e�9B�冀�� �����N%&�����U �b�"Z��]\���� �����{��������o����weqy/|��/�����'&f��t+�kB��X��$]9)�f��!s[D8���@��#���ހRg��CtQ?NEͰ<-�:�.P�9�;!#���i�j���	�.
��TYQ�S�H��z
��	b\%��ñ�� U��|��'�E��Hx/�м�ق2�s,�(�ąׅg�9zM��%�Ǔ�X+��S������'!���ar�Yj{YE׫a�EϟT� �w2Y�=�Z��!��3V�q񪸭w@����*V"x�^O�.ЎxT�6nng)�m���_���̄p|��=�����(GE���P�;� k�(uU�N��\��[|_��Uxj��Ί6'�m�x� ��.�ؚR���9�-{�K��=�Q���7M���gkN/�ԇ�sKUC�4�0��g����� ��|U����v:�ށ�ѤŦ�	Q���U ��|�X7�����g��u�Q0�ȩ�%*��NcyZ�P��K�D�?��\W��u�{��S������g�ӄ�F�$j`�7$������}������+����F�X�!l�,O�3'��,`#B�Z�x�H��Ő�v�Z�~2-�~������ɟ���P�����zy�_��]�$.�\�2&�(�Dצ��R�
�KDƎ/Q�?���X�L�.�pʻ�|�˘�޽}`�Ѕ����
���V�=����C��8*I��ӗu�T;���K���6E"k�7횩y(���|�&�zh������'O|����<�{�s�_~n��w�=����{��xn��{+<pQ���r��% ��`Y��k&��"���5� j �H��S�A=]X�P<��#��k}ZB�8�w*u
 �%���=6�N�]��z(֣�F"�8|�R<R6C��9O`�OO@--<�n�'���9�(����2��'��.1($O��0�r� ֎p��������`8nj\ا#7�2���A/`$�'���|�=���A?hl�1B�SD�xH��e�U�|�y^��T)k�M�����W��zf�M���E�/�@�A|T�wRY�����������mOQ=�=��zO �����'4J`����Z��Ox�{��b�A����|P�!�n5��ys�ƛ��|��i��t�%q�ծl��P9<prH����H�3�jU��)K�[��f&8�*D�97�J�[�4�4��a���f\�x��{�a��g�
Q�� @￁+����H�s�=	yt�C�s٪Q�jPH��n:�ը�G%
&+V�`��놬���f؟�W��<��-���99|B0Px�e^��fI���4:�ֵ���,G}�lܩ��(�ު����u����ˊپ�7�˽X5���K�9�����W����Y�+1R�����j�1������
������7D}�Ao����{��}^(���f>���~��������o�N?-S���`�P% ���TaZz���(]�~�
t��D
5.�&I��U߾{���/N_�9~�^�7W>|�Z� ̮?�ꁹo��Ҟb���Fh�]�T4�/�3�/3���ړ��C`}*���<�;���h"�|��I
�t(�Q� >�.�d��4z`!� �z;4m��16*�K��YI�9�^���r%���)�O<2��*�U��#���ֵ6V��y��Wv*���1��?�����J�/��(Ę�QTxK�����(؈֕zhF�74.���)���J�)-(�1�o
��8��U����q*���`f8)n��ᬎX[�� �Kٔ��;7��Ԯ֋�R�s7�%�m/M�qQ�+%� yDQ����L�%)}F^uQ���%�W*t�FC��P������ ;�q_r
�'[�����0jۆ�r�'� �l�-{�!�#�"F�TB�Y�H�LJ��^�s)#߂���0.�,>Z��C@Z�N ��u�j�G���6s���hp1tN�����k��Q�u��W�[C�ҚW�F�WM������F��<��^��85�,��N\�<&��j��F�Q�4�����FX�hܠ���V�H-jG,4��.������'��:���W�;>����w>ӌ��7��`
s!�h-�J$���3Y<�ͥa�x/|�U-�V�L
�����ށx��k/^N#�;W�y��y�W\0�����'[����#/]E.�B�#�[�#����l���	c�ǣh,��<�h
%X�(�P��E
�fՏ��5;��}�&��ᕢ����G��4uϳs�������<��ܒyw:���?1V*�M��BE�� ���������Ћ��GM���51�L�˱ �X#�baKW
U�."Q�|Ȗ�PxI>�BQ����0�)�ܢ���h�m�&��z�T0��U��b��6����d�qG�X1�&�X��&�Wj�3�u�=2�YC�~;��kM���=��A�.SB�b�ˑ!����U+��b��P�aw��r�k���Y��)�s�Hg�/��H���y�6*�}Dx{�y�b�/ڈ����n�/��_�;��-���
���~����x�?�g�)�uKN\�_��9#��T�֝�Ϲ?UޱF]�C���h�Q����  �:IDATx�k�Pk�~��c(ċh��snj1m��c�k%1�g���DL��ٴ�ËHy
]@k��4&�N܂���Y3/*VC���sjh��I��t�A��������!k�{:'�`�ۂzgn[���#4f�lq�Zk��F��Ƌsӑ����Ay*�9�r��FspP�U�������^��F�vP��:K�b%_�9�o�t��W/ݞz���������������vǽ�7N.�?l2�}�~!�E��p-_�L��C�A6��^R~��8y����Z���_�϶�G�����]�����v�v�}�(����e�?�n�qp~��hj�(j8{�0tU��+�pKx�!db����iW#�&<t60�Aq�3��C�t��z��zφ�����=ٿ���t����>���~jۃ����x���<s��я�|C�I�2k��j_�(��u
hT��z)a�#mm�X��9siw*9r+��0�l�����(CA�@�uR�B��|�T^�,�fZ?̺oI�z�H**���D�r󔗠�%���Da���=-�JM���ֶxJOI~�l��`��ǆb�@聟�P?=x*~����)��(���
<�Wrᱧ���yR���b'�	j<?���:|J����1�UD��h�M9��l�����U@<���t`���3�	.�+�X� �N�Pq���䞖����yt�Ġ�8�*�e����WV\hX\�UV�?�'�jzT>��%�4�����,N��2)E���8���FL4M�)"k4
���\��0�i�Gj�E�[c`��<�����h@(�E3X%�S/�C_��:7�a��z�0�z�K��[:��x���h�rn0"�s��W����T���#��y�
�B�q��c�߁wz�avd�Q.X�	ƣ�:�V"���� -�Zd��F\M�;V��&��qǭ֛��	S�F��c#��7]���o�����ṫ7��W�?>�p�ϛ膁f$*/�VZ� U����S��e�!�~�m2�2��!��4h@�[q��������|t�?��|~�Q�|6�]������}��V/�<���bD`WY����bRTD0�R�O&�f d3�j7���Yj�iC�=y5É��~��<���M+to��>�i~ǡ�߽s��'wL><�����snt���-�u�q� ������R�BjV'%x�%��(��N����*y|�h�� �@9k�0$/%p4��\��6�3(#�����NI��Xe˝��K��X�p�wO˂LI_�z�N����QHσmE>	�L����-�!Ɓ�����.�����P<Ao+��VE���0t)�żn������9{w��x]�(��O�r[@��Z���F!�T��|�ۓ�����S�hN>�����;��� z�޵y�;M��\��=O��٬<�=N��+O�â�Xʻ�CnG�~�+@:S��Ѓ������ j��:�2Ϭ.x�m/��qS*a�(���D�8G�%�Z�d�yn��G� �B#Q�x�CR1��Q��Gq	�ktEJ�$��νǫJZ=����O��ʑUÂ����X��\% %������=x�1j��ox�7K�\��k�*�*xF��֚7�\n�V�h�Q�gH!�q�*�;�T�=���Y���i5g��ߵ}�Љ��ڕKw��D��L�{ܵfvɹ��L��_� ����u�t�B'�+	�X�OD\}&�%��O҄��u�k��CZŷ�
ת>pن�}�d�i+��f����y�������|�x�8
�G� Rڂ ���.c�1�*PZE,Nv&^z��虞��l-d�J��Hj�2�
Aj�L,44z��|���s~������&Wl�s2������;�=����,���>l��-�({���U�3�[g=�
�B?�1�DG�G�N ��Q��P'/3�=���C�`���B�Np����m&	��nh���LQ���6dܩ,�=QYq��(0=.��˃[='
X�}���w�x�g#�8z T��^���D����^j�Yc����2� �0�-��#��-�C��ʄ� (�%�茀��;�@"
�43";j S@�L����[�"�~�q�h@�+ Q5�}�|Nb�X]�	[Q�D:�]<��9�$:��zʄ�]F���QkE��\w�N�,�������}ԭ�c�W?��8i�Ĭ�AO�r�ԫ,������8��������4{�Ng��5���8=_�TԨbT��6�)�* `�:᜔���}bl�b����Wb��N�~%T��ʟ򷎡Г�ow�������7�`��60i[bǥɾ�|�x�)Jɬ�"�8׭�)�b�k�0_kX��1�9�f)��>�^gC^�\7�
�2�]�L,�+�pb~aӦ�s_��[g��Lo��_t�п���?��.N��x�$U,��F��i��,r��C��t 3({�F�Ă�p����,V��ٱT�k/[}NvT{��?�:�]W����=��p͟L��L@P�TRe(��2H2�)���JB���U9@���s9�2�& d�JmU>��W���>����`��!n�t�a�_�{��߷�����P�7�~'���E�˽Z���w ���g2���Jޔay�A�XȂv��[\s*��w��Ħ.Bln3/��c�)H�a�{�-(�X"��f��x��S�@,��M�h۾zT�hT!#�YQ�*%E�YO��3'�)����@<^+�'����Ņ�hs�>z�<Ckx��>zҢ$47��A���l��.dV1��]:��o�3k�7�ߔ}���(o���:�ne5�zh��5t�c�1`�9��T�j^FK���a˝��@���4�}W���_��6�/�bU�ZMf�wfyO��r~�"�!`�x`�Q54�CED�}��yC�$��\B��W=i�{[o�s�Y@k6��ʝ���M�����$áA�]��P�)�SGɋT�Z��|"�$�Ռ�l���lc�4�ƞz�	���і�lA9��È���b !�z��y�L�=�J���0�Ay:W9^�a�֑�� � &D4��%`J(W��� TvcCfʤz�� ��^\G�AGtD���@�i6g��������lJ�x�uWO}�=�:����wO_4]���r	�Cu�iT���W��L�`>�:FZ�a}6ʘoN�E�T��(D<_7�����t��s�o�m��;-���������_���B����5�Ayw��],���$M�N �h��R)!)�Ë�_,�ɩ3�-����O�D���[�9�'/��5���o��o>t���b!��w������%/<tc0��тM�P�p�D,!�zz�n� b�M�Ŀ
���<	nn�}) Pؠ�����p��6�l x�<:��Ǔ��O����P	Y���0s�PR%䁺< �Ѷ~�^�6��*B�mΖn
֬�kS Z� 
]&yp���r��U�^�r���ʅ�{�1�\L9��C�
�S�{]�N�˕(a=�W*z�S�*\
|��'��T�mK��r?*��)��uU�`�{���{ц"�R7\#y�����w*o܎��u�>���vzل�=<��r}!�.��ip�Л�>cD�֪��{�r�,���:OqM��|G�7o��'z$�Yc5�2��amǗF�V;,�*{�w�@��&�A�y��l5�1F2V�In�
��B�DaQy��Z����ԙז�~jWC�'Q596SJ��v�4��:a􄤂B�8�D��?Av��!�/Y�}x=ǫ0؉�)#��>~�k�&E���P�#2'u�/�Ɋ�ߪ���=���)��������t���>:�\��bL����>69�O��]<�57���a'�N2���Ni?%��v�LO�]�O~�{�/�e�M,�yg�&��d�(�Z�ݛ���~��G��J�yG8�<t>�뮼h�����l�I�]�ɃNk��(��^C}�<�a�PrP��r��p�O� aJ/�F\"F-x�N �s����7���n d�-�~�#�'..M�~y|磏O~�]�gˁ�[��&8���h!�ғ�r�(Q����BoVLJ��)���u��N�ȧE��'M�W��ts���z6�	b���aC���Ȉ2�ǡ�k��m���#w>>��zX�O�?��Բ�ygC���U�H�@zyg=�0eт���x=e꽯2Z�a����}yd:�1���~Yڣ׮�=���dm�m�A�������՘X�;����E][���ed9�[�zv��B{�f����
}�:We�Ut�W�����|R������q�w��ׂ����ed��><WU֪�靪�� �QI�����G:�֕�:�4���-yo��MӴ������;�X:n�*QcA�	�^o�ȍFE�'cb��2,�NU�Z��}��D9���eH�@�h�Y!�!(TX4j�ݸ��X��秒�!�Ůf5���֜tzk ��b
/�>�<!�&�@����c�N/<�:r���W[nu)�������/_���W\�7�+��V�v�r�?��׷Nͅ/
����(L����Q��r:���az�A$e�����H�L&;c�kr-�O�S߻��u��u����y�����\<�����>X��U�����&'����M�(�Y�La����4:<�,������"y�Z��G�z��?��/��'ގ鳱'C�D�ɧ��ǿ���=���|���pr�ߟj4��9�4�B��'N�=׃5�l�P���x�`[yQ�̷'q3�q��b���sXC��������%<-�������$D͒ ��׺a�WF�$O�����E��E�
�S>©��Z�����B�FT�y��M�+�েm+�DHo�$����Z�Is��r��a��]�)^Y�Z���R$},��9�U۪��!�a�S*��7��〷�u�-w�R:ލYﺭ�T�z^���(� �L܋��8�b�[�CP�d^�N�o?�����E��~e������ۗh�[��T����S�;dg�"Ȁ�w������+��{rNz��jnkL��EN�_犀�T���Ҳ�JX˩��@��,��<"�u�ܐ�A��t� ?�=��P���YbV�#�?�E���Fz��A�
��]�\x�T�Me�DY�*e���B���M}�o\�q��7�μ���[�x�rs��/�}��τ���5()�k�M`�ϝ�T�XЎ���(�~�NAU?�D#M�$������ܑg�lJ��+?�j���}>�w^*t>�K/;zx��csKŋ�N�s�;��>��n�z�����'a��� ´7�%֥��ʔ0�v��n4�9x�3��ԕ����-Ϟ�|��qĆ���m��#����.�x��}��+�<=W�������5|�H��H�∷P���s�� 4�@g�/�1 |�@�dV�M��5(�a��$�߃��;�	�-z&4��z5�[$L�rv%Io��Uy�Y�����ɘ��T=��2FQ��(���VyMB�|F6�j��8��5+䩤xn(:���Y���6�9tjE��^e�-}�"k`<D�P�Qd�"��\�F<���^V���YĚ���t�{��g���v�~�ն�ѲR��Э��ʃ�w���r)�]X�?� ԆW��~�Fm��}E��i�����,_���=`�W� ?=���^ZB��=���������=�nfv�$�nC�z�6�Qk�';�1W�'w����u�e=x��T��� ��@�RFd���M"��&��$5Sb��ٙ��.�0UD���YCB��Tq��.��Y5��w��_w���/�����O����Õ�?���������
��� �ɣ���б��Y˼G`%�U���D�����$�C5[٩�h�+.Z}��}k/�u��V���k�~�O�xba6wk8��ݴB�fҢ-C�E�XZ̼��ȟ��N%M��`�B�� ��eI@�$B����N���}�z3���=+��	�e4����?����=��]��� �����"�������J*����B��W��d��A��q��(��gs��e7"J�'OT=��(A6���6Q��Z���YA*4��-�k��D�LB����%�ks��/��¤���xA"�+O��Q)���,^=��m�UJ�p� ��|Q))�z[�]˛;ߑ�����at���:�"���s�&mj��u��&�;ɺ+p�3�g�Z�B"	��M!�y퍂�s���ۓ����_+����n�q_>[���/��L0RӼ|�b(خum����knJW�)s�mΧ�s�*���4���ư|G�D���o@�4�bǃ�;���(��'��4��4'�]f�OFbhD�������1`[���b`���B�WJUX��J�U&R���"��'�P3��F^�
d�#N�k�YF:͊��u�BĢ��V�@���7�Ӽ��Wn8|�ţs7m�
������9V��fb�x36x�ސ�:�DT��H�#Q�bf����0]���L#� ��$���)Ͽp�O��6�7�p����[���ؾm����KOW��j������<�;1gU��ʮ`�z*JCE�$r�yt�����M�2#.�=�k�D��Hm���/\�����7��6����c7�ƛ�{o���;�����9��>��o����@ G�b�#]rJDЬ�V/8DA��e���U�/C�T˨("��C�,���a_�F�A.m9��!iIi=W	m�K�F�����a%oJ��YC�%��r�
?IE!|o�7Ξ�mp�*Ƀ�7�����(���:�=AQ�iM�ܐ
r1����Z|�w9�+s����>��ۋY������rV+P�����_]F3ѹyuUD�/x�FJ��T���<����ӴѱZ��=L k�n�S��0|X^~ކə}=Ղ��%n�|<DG��3�V\���e�WNK/����԰�c�z�J�<�����S��|��!����WI�~�R'�����r5����/�ʼ
�����?��X'�c���z)�R��!���P�1��D��jyޭ�|�]�@uǚu����z��_��y�d�(��_.'����{Zё5�Vb@�����cT�V=�Բ���2M�X2	�c	�<�1!��}��KD�m[��Gqo?N�<�����y��G_88C��w�5D�W�m�*�u'IK��R��"��=a5��b���0`Z+��w�^�X��:L����v����mɥ��dz߶�<>��d��ޗf�z���c�w{O�-_�mB��� ʉW�)tB�)��XB�+
%MaMo-
��aꮉ�s,��c|�4�,�S`
=�P`�G
Z�����XjE��5�
�ao�����r%��t�~�AF@X�%,�)-]�V�
��<�N�^�6MQa��(8�RV�-s���a3�x�<-��镶��#�^���\��M{�C=H޸ ��k��Z!���B��(��ƎT���읛p�X���)�W�w�P;-ބG���:��Sr�v/Tm�
g�n�S|6="-�^������� ٱ�I��f�aޓ��".z}�7��O����D�K���}
� O\�9�ˀOߡ!�O����z���:y�ÅN�l2D�]B���cdޓ2K|�.X;���3"�P��0��wȯ����
�R@t����OI9�Vei���=h,>?>}��-�;��q�����u�������C�V�?�𱲓�%b�&��4n���Bǐ�[�ȑg����вD�������[�B���w��̣m����ُ��k��}0�~�������L�ѳ.��X��Dؿ���VE.��w ��3��ؑ(B�	,�L��j���Q9+�U�� `*�T|��z�������nY�������]�Ipۙ�|�q߾c�}��=S�M��\�s����h�5I�
��8��<腜cCD(�P���0�
�9�碀!��o�Z3y��h��w�l�E˲?�b�ޛD!R�C�qT�z���R#�J��*k*�؄C��ee�]�0����m�LU	���H`4,��kM0��[	���eC�<5�J��H���T5�Ge��i*F�)�Ty'��YW(�J���J_k�U��}��T9iY�j6���ŋ\�tt�B���e�{��A짗��y��a���r-�$	�Ҫ|��]�{�wٶ�C)����C�[��v�$ё��A%d�q`�G��-��������侁������.k��mH]�Sٮ��G|�������[�u��֍@W��358%�3�ǣ�H�K�6v4#x��w�£X+�A{��ug�� �q�\�HB���eT��[���O7ܙ������o	>r�Ʊ�Wo�8�������R�7���۪f��x&݊��}l����ƨ���J�c��$���f�\�}ҁUB45�R�H#7�-�{նmG�%'�����
���gnY}��ở=0wU��@�\O1a�<�d��eWl�Ҁ�p�� r�(�T$-E �Q�&����:�Nԡ�H�ޗ���O�}���{�Oe�ޛ��3�c�<��g^��tzi�*�y]
b������ 9�#�:�����N��P (w"�U��
�kly
ˀ@z��N�5r����?�㲟;�R0>ax$f�R'�[T�I_W�^��m~��UBߪdX��M޶Lv������v�Ҿ�����O�{�/
�o�}�W�E8�����O%���XEJ��ؤ���(t����A��5<�SCz�����o��;�������ϫ�lK�p��l}��;mf�N����qk�ƈ|�����0����&U����ʔƢ*��B��Q|�r���E�� 
����G�w� �ȅY�d
F(�L��E���O �Fypx�K()cx\���Qiɚ@N<�p<���/m�Yo��ah*3֨7`%H.��V�V�\��mL��7�����nX{��.Y����ūֆ����yvhϾ�ۂ��JxxD��y�c-	IapӠJ]p2����C��àc�Z�m�^Z�*��/�6�h�y���
�3��7�;���K�"ľ��
�������))&�5,&Z�5xo\0�������@6�˙QCv�(	6�H08��������+to���~_x�x���&�x�ك�;|Y���6��Zł����%����A��ޱ�jL+07*F��k�T�lUU����@'8�vei�w�IlSf�)����'3=�#
;	yR@�r�b� #��J|끋�Ge)�.�J@Nr�P�a;}*��B�c��^����R+t�i
=�"��¿�+ �'����%��z�
�{�M����ʸ�U��kd���;�����ʃ�W�^~��X:ޝ6���_�D6V��yƒ���ۿO�6�~e�����(m{-�2i#D�۔�hg-�~�sk�'l���<�m $ώ9^pܑ3س�DNo���
�;Ցg�*J@+�fȖ��}J�r"�IH��^�/AD'�q�E�KJ�a}�HFI-�F��[-GC�R�Y��U���c��/�Pd�Ʊcl[��ޫ~<���g�Ӈ�����{/�5�@"�@>�H3� F#v|N4�8�8��x����U14pB,i�1�"-l�4�I��b����^Y��']���y}|j˺̽/)\�HdVe�y4&��:iS�d'8#Z!4�>��&@�3��ρ��,�` Oe_k ��֬`dk5���]w���'�Ͽ���?������.[aXN��=7�����z�?��|�����j�`�oC���=h���5D�P+ЇyEv���bT�"��k(c�Lhb)o��ɬ�<"�0
@�a�x�;1,X.\z>�	х�%�H�j��k�����l�X�~�ӝ�Y{ay���
��z�
*D���*j/W�����v�s���g+�eo\`����G����kkl�����]���J�ke��S���ӧ�!=��<|�J��&���cp�ɓ��r��ep����N�ڮ��O>$.�<݊��YD�e���M�-k��<P�����k��&�BLBցK�t�?9�@P��@zы�0(�m��*�:_�(9p�	鎆e�)EGD$�P1Y�PB���P%����% �'�OG�9{=�4$A�u��\@mlq!���r;z⭧�o������һڿnס�O��G�`����A%���z\�^�
��"m�PL�P��L�V���/����[֞������U��K�{������'O<3_���D�k���yv.o񨔥@��sQ�;�#��i�6�6��i4kA�"BlM�k��0�7Ra_k��;�ٵ����7��}[٘ެ�p��}���➩���/�|��2;_��p6�>_K^�$�1_4*�������!Հ���d�=�Q�]���ȝ#=!`8�IHy�2��H�%����F��pu_i�MR�l	#�y|AS�J���5���ݨǥ�9��=A�y�XK�5���Ϣ�R�a�!��U�* G��(G�Y��a|�`��eؐ�d�W�۹�^�aە���X��47�^N�1�ӏ���ڗ}ڹ�6���B��wy�VB�\:|� �g$�n�G:S�v���<'ߓ8�^�����5� ��g�Y�o;j òl��/z�<�`)��D��}3�˖�<f�s�A+D� H���C�G,	�%���}���V�C�`�#)�s�C���.b�[�r���@1��i6jy�F������ԎP��{�?����ٛ��`�'����U̬�po���f��;�xo�]�w�i�A-��>�Ą(���HF���a����eˀI@<�th�y�Ba6�?x�E��{d{�c�*t;o��8>y����ˣ�Ѿ��J�#���ڈB�;�Wd�^.Z������'��G.�TE�U�٫%6|�� �a{@7���ƎL.~�;�>�N�c=	/NQ�mi���.߱g��ώN�-m+T��A5yQ0����6��$"�
<w.N��g�\�2zd�C���c�8&ГYB��9'�V�x:�E�Y��HE9rmp�� �V<%���A"�!ݶ�w�N%4�'+���-�*
U^�D�kHVC{��7��}�)�%xW�F]�١$��W�������&_["�
�0:=�^��y׶|����_��^�B�Q�yM��Z�I�֝��ʿ v:`P�Q^���^>C����E�RY�0x�bdX�l-�e� ^O�}X� �)��(H8]������h8"�T���a6��+emA,���2f�׵U�G"��7�tbd *�#N���p՘2ү�eV�o�C�?F�HT��q�@��(�E_�t����r��ݣ}���gf�m]��o�h:c�I����������ޡ (�+ ��Q41�t�ikg]?��S�|Zx�ƞ�}�r��fu��͛2������^{U��t�}��G���������w=_*$���x�r#
��lU(�,�&$	hj���[Z�y&��ux�9(��j��]�`�Cq���3�\%~���ھc�0q�:����^�ː<_�_zt�ޝ{[=����'O�n+�[}��K�Nz����� �T�;��˱O&u��g@�O���P+��� �G�]7�wH��An}��	a`"<&"��I�2���lˇ�V���̻y���1i;��G�{�6аr�d9V��+B�������!�5��X�2j�!_*s��T��^��G~�9%:
��V��md@��՞���1�טh4rT��xP/-!�̶ܩ�� 8�c_�_>��q��
�����xQɗڰ3*����jQ��g�@��]��(S}��s�-��9�C�:.Rh11l\�z%�X�������6�`�ۢL[h�5��k=NC��wI�������m_�{�{�ϡ� l����z����U>�o����l�p��o�ꞓ[7������}[&�N���T���~�[���V_$�i!� Q�V�yII� B���3kH��� J*eD��<�<;ٟ�~�6;��x�B�xj�\4<�q��^8���狮F�&0q"W���GIæU(�:<���'3CA�X�$�-#��r6�-	
cf �M�>9y��N>�Ӿ�j&?{��硞�/�=u蹗&�w$�jzq�|�yI0]
E�6�V�$<�(�޸h�"v^�%7���Cb� kl�^�AJ<(�p�>$�0�1L�񯠧3ڿj�v��șNh��ї�*Y�8�u{yTz�m���$oI�A�̖N��ɢ�= � ��$-k��-�<Yދ։k��C�s�)�[w悅����[2WC�a�����Ew�v���b?z�/�l5��LV;����v�x��K:�U��>g*��;�1a7�+>?���MmHDBC�,qT������8�� 8���D�j5�T����!��Ta`-�b�&�(�8�	�R�5B��ۆ1':Ej<�a�m�)0}"
]qaO��4*���b�h�UN����s��x W�`�FB�ÑP녁�ȋ���O��/��Oo��(5;[e�k��^>��P|[��1��D=0����&8��A�'QI�^��l�Ƶ�f=�ܖm����g{�����
��^=m���_>tr��e7��Z���=�PO�V�vd0�\�@j��T��@8�V{�!��P�u�C�}/ v��57�_-��'��|'*������3�׉��3������=:��p�b��ñ������éTQ�����S�E.w
V:
Qv�r��bP9�xM�L+�nL1�C�)3�U��ꇰ�=�8�pt��5�J*e�, GOA���Er����k]#L��4w�p-��F6��lQ�ֳ��P����ڄCL���f2Jx[�'}���"
�>Ñ6��NPYP��i��(߷:N<X{lmB�RT5%X��Wx�TfڒS�O�W�w�<:]�6�k���N=��!�z��陽{��p�[�/?����&��:>�����a!���܈�G��I|��KǄږk��~ �<%�>�<��yF��hO�/v8�8T��pU��l�D��Xy\�����Q~���qXgJ
0���S�;N��(fMmi��^��m�OZ3��Y��/���pN(�� �����`���!=ړAPSb@A(tvF�bH�c| \�t�����$���T� b�Q*�@>$Vk��;�;n�x��w�����@W��6�64�f������ǇЍ	YazZ����`�lP̘t��Y�~�(Y��dL�j�Jޔ p��SD<�D(�O���.��7����+S�	�o?}�H7���7�س��t����Gg/���]R��6����`#Г�H�B)��3"�&�;V=Q�to�c���r#U$�i"!޾4G��"'- iX��8yb8�����j�y*�$���%����8U��`CQ���i���6TGp�vUb�ͪ��,��ۊ�RE�?��~��^"�����ѣ��S�m�goz��wݼ�f^_顯 ���Z��)tkٯ�S65щ����^��d/��A:�Q���`��w�5Dt<��������:�~J�sq�	�d��bH�w��H�7��V�(��ј �#q��Ib����v����Ap�;>v�S~JۅѰ�[�f��o��h�H�O�=�U?��6^u�n\�vnˆ��/ܺ��S��߿�8����z�ċ�zu�0�1�P���(s�i	�����D\HV��Uu1��|��^��r�z��M�{���+ǲ�x��6�@W��6��E�qϑ��&�=R1�1�M�����+� θ�!_b:@4�{
QL�B�lRR*��ւ�^C��H�����*wK���B���͝O���<�uut�׌�3����i��O����їL?���\��\~��lᢚ�\�$VC$����(�ıx9x��s��: �؃�B4��'�86i��He�|;���&��;<U��+���/�UA9 &J��d)\�����2�Z��xW�ц�=��`����.�@|�#l�aZ��9���l�X�b�@��R̩�ao�jF	�'���^�-ۏ�hXaPQvnL󔞧�=�F�^��yN#�%4.:ٟ���f����Ǭn`:�X�L��$�I�$�(�U CF�^�g��dR6���G�ڎ�T[~�����2��
Z�^u򽘎Ճ���8��22T�4 a �`\�i4"�	�+`.+Vj�b,l�����J9=��v���7��_�i��ɫb��A�m�?�C�=�8r�Do38����/�������w��Xf�>d���a=>�/1�H��t�x��Mr8����(8��ɸ����_0��~X7�;�i��w�տM���t%�����q���Nz�{��$C����5��#&�$�����&@��e��\�#,_G>7[B�ݗ4�z��K({�U�m��R9g�#G����P����.\?|�ƫ���r��JI�6����w���O�'��u�������s����3�נe�����������E�p�/�����$��K�>���$�h!o�+B�9�&�<x��D_v(wU0Z���x�;*��zp��CTY�(Щ��q=2K*jn[x�!�07Sd�B���z`=������d3�����{�����ָ{�m����0�k������ČR�`T��4��[���sO�mc�m��'�nrM�mc�mNz��d�μ�sο���>{������O�Z�2_.My�Xyd�p�H�R�2��[�9��{Әy�o_���qeze��#xh_��qoDpuU��
�>Q�3��S`����`j��aGa�,�|Q!�I�z���l�*�鐫��i4xwͯ#�^=�WI������zM�u�ç`�ԗ�|l�y����k­Q��=�w7Q�$��O�M%�l?��������U9^�vKH���'�(���D��"�Aڲx3�HRR�i*�k�����If1���5H��ށ7�t������6�r�F���yc����Ϗ���V���X�똕���3U�V�|pZ��x��rrY7��0�r(yxJڍ��d��Ϙqj0���U8�d�@Ǎg����R�5����b(x��n^��B��#���:�f���!�w�qh�6����O����pf+�G�5�<���
�EA�-6�(��4r<U�x�Z&+i�S�]�r(.�Zʅ��n�)�&9�B}��N��ֽgD~Y�^.���#2$ٸ����I��YҧH��2��I<1ׁ���OਥFˀZ��^�]֒F�o�w�n=��ܫ�J�r�t�����E[Ǚlv�w���j�j6}t�v$�x�H1GmXHYr��H"I��g}��U�%���&U�6���}�R�-�u\��v=�B�>^�KϋV]�d{��q�pC"�,0NU�:a�Y��*��w�ѣ�:���|Z�LDqY�RE�S���^�E�s�V	Tc�v�C�o��,� �����-�]���h	[��f�z�YFn_�p-�u�@i�$D^A�=�UZ"��IYU'b�q˹q�1)���L�е¾��9�����s���������ڶ������4(�}[���֑�����4e\�M��?��B��'�%:���\L� �|����n״� s�O��92X�`��8������M1o�h��im΅����}�C��w��1:����p��s�s~2�q�%7�<��T���ˢ����NdL_�=�i�H�ۺ@��2ay Xq�"^8$�\4"���/��k��Z��em�/`�������
�
E���~4Nq����E���g�1l�ކ7���N��>_��7>�*�?؟��e�˸���(�L��Bg{���c������~��-�?ߴ���d�Q1V��lZ�D�ί��=���w������d���#2:��³@��K�IN�^4�<q܊1��8�u
��#����끆R���j1X���j:�@�I�
��%��D�$_��OZ�K�]��x��n�3p���8���䣚e+�t�b�����ZR��l���#?�~ ����y!9C��O��8&I0���ɧ�j�	��t�ܙ��:D.= �t:�m�"�Cqa-��i�����~�����ۣ}���,v-us�(�yna�zb�M�bХ&-�j��L�I,�\A��@\<� ��xx�%3/�3|��2��me�Q+Q�J���1�pj[���	E�h�Ɓ���}҈�B�9���`�\�}�q?��v�~�>�߸\�4<��(K���D_�z	5���%f�6�{�Ҵ��~��0�E�5�oY�z��v�_|���5H'���@Z��9O��o�J{���<�����ؤ�v�#�v���)�N=���o��������,˝���&�B�3��$����`ˉ�]��S��/Z��[�{9�	�g��c�M��1���q~,���������/+���΄���vի�S}�ڃ�/�A&ێ�*�������O���mtXo_���6�ڋjn�`>��۸������2��שr���!��y Ђ�������Q�j�ފ\���a�8𮏸�e8��f`��.��J��Ξ@9v�'�R�0*�|� 58�/x3����n:- �BF�Ƀ�*��6�s2����[1"%R�̐��^k9�v�q����wN�M������������"?�+F��ðP5A3� ]���&Y�`%Q7LZH���x/�+���W͒ݪ�yc��6��:�fs�!�Y�����	c7T�?2Y��J��3yO�����Y��h���*�*�$�	Ȱ��d,��T=1�Ze<���}��
�خ���% 	���`�˳T!
��B�!	��շ��D�?�r	��6Iw����U�&��k.��b���21�k}ys��%e�?��縄�����/F���l5X����uR;���B����ك}1ũ3`ٌy|���[�:�n�X�oh�on�nA�%�l�'�d;K��U�>���w���?�z�zxz6�6����X������Ao�P�9a�ٻV"(XK���c��^�$�z:����?a@��E��ժn���юs���^��e�M+���Ow��p2��ӪJCW>Z��j!� Y+�Ʋ�s}�G}�go��0�J��u�|��c���kZ��#�Aɀ���(�<�ܑ�a�,12;�h��:GE7��O�jrњ����:�ET�{1���II���Ͽo��^���?!��v�=�"�z���W?�\X���qJp)���23u9�]
|����<l�-� x��U�|�P�p�n�{"w���2l[��,�C��1[ �/ʫ�ڳ��z+�����~����^�}m�24fcs.ė��59��yvs~"Ҩ��7�gsre�l�±�q�5�,�4������.�:�!끺J����>�H�$(�,�N�K���yѠ��s�_�� ?����A��ޚ��7�	��K���N��K��Z`+�\���g�^��#cR:�ɭU<ˠ�;'�{��kpP��n��r)-���$B/B����}��4�H����4���W1�`�/䥀/���U�n֩�C�S[���vQ��h�P\���t���p�2t̼���xE֬�=��8�̋x~�ɏl
��ʼ���
��'���;'D�R�O��W//VAN��l�o���B<�۬��,�������҃��?�$k�,i�qs5]M2���R0���Y3x�5�`��<�8�q"ɐ���+���~tإXU�WBF�=C6#s0�!Չ͂�Nm,���g?��L���>�c�ϕ_��_
�l�o��)�Q���
u�dz"b���^�[2���2!'6����ҾA�6�B�� n6�s2s��ԭ3�l�]T�(,��u��Ex���X��(1��o���a��8Nb��'m�o=L���}U�Y\��<�p��-T��u�t�Ӊ��31VfE����cЛ��1]'�-��E�^l(��v+�~AZϴ����T�@&Dhޓ�DBl��L�^�[f�稶��DJ젍K��B��Z�\|R�R}5���m�����f��������G�O-�6�����T�n�	�g�ݰ.�ǽfˈ6.@�(T���Ĺ�xh&B�\�u�g�v�����vL���~l�Ƥ�q�¼�� Y�2Ğ�s�|�j� �Mr��	��>U;����8�@��5�Q�yU�N���w��V�Q�JEg�խX� �&��q�d��b"�sǭ��F��aL.=��=������>���$ͷǙ jB|C��vrw	LYw��Z Ι��
%jTa)�gY��l6� ~�0��9u&b�Hu&�1f�w��^�62)9���P�B����QBFF�2v|l}��)��o�����9��zٖ��R�?\��=��mf�^f��]S������u�,E�T�V��3�=3Ly{� �T�P�}�4m��g`𮅬�{T[���wEu=��;���*�XS��������F"�//3��4�~��u��k����d�o/hp�m��Y��
	4'�¯��vrv�y��p~0�A��/2�DF�T֣�x#�P��
/h�������O����K~:X,ˇ�يE��{T��{�/�n��])eL�b��NQ�Y�kc���j&z�R9D�[z�"N4街]��C^��@^��j!��3�g�Rs[R�c���Z�������}8���vK*"t>���u��ñ� ~�!�ԟ́vc6J&yQ�хgư��R���}_Ȥ�_I���!�m\�G��pW��M�����H���B��t?k�6p.X�ǁYO�>�'�Lo$�u�c��a��}3?��%0`-R�����֩ٍ��^_FԹ��I��:VF��<�L�2Zs��y6J���~�r��4�@0�i5�*L wJ.���[�-9?���<�O�z��>���ǟ%�_��y���k,B�U>�e 2=b
����:&����.o\#o��J�NS M����
&Z�� CR6�aX�w)/�=Iګ�{q#(R(�� &/WE�50C�����.�G�%�G�'�1���1��Wu�7���O�N7�v�3��VC'�9�JT1)���u��P�2m�c+��� �T�N=��ACzm_[Vbx��#.q�FS��%�`n?sv��rN( �ݤ��La�̔���1��+��?CTa�}D��7*�x4Nwm$SY\>D`�������QwF{]"z#l���ʯ��u6}����/ي��(sX����n'��稤�����8�PqK���ư��;k:g�Q%�(�z��a<D%���\� ��=��09�KQ�7�^�h�;��3�����ZH�	(O��?���բhS�A��z�(��������?*�l���a�B�얩J��1q�d _G�!x��C��ԃ�4�&N.�j����j�fn�����_��ʩ��jm@��.F���6d�p]f�u������l��~U��0���El����]8�q���?�y2�V��1hā��!t��
΅��)�:�xxD�g\�Y7�JPh�U����RA%Ry�ps����4=����aا��R���)\S;Qvo��}���_d�S�^/MU'����E�v,� ~OZ���̰X@Ҕ��IS��0�u�A�%ϥ�6u�W�m+V*t�Â:
�#��cL�4���!�"�ߣp�����1u�*/��0`����@RH�L�b~y��\Z�	:
J�ɟh`?;YQ�%V�jش��̯BH̙8�O��׌�mM@N��D�t>��û�h�F�ѥ�n�&��`LH'�
��������7���å��B�������g�XhJ,d]F�~T��J#��#:<���=z�!�L�T�L	�k�Z�:|�)>��8�%e�h�7�d���+�O���Z��P�yms[4�p�Va�cpY|	�_$ش������I
E4��\�|����#�"��@��p�dZ��,u������Z���o\��P8ڏ�n�W�KnX�xCj�����~��5�
�?�OnZ�S�OEW�g���+��u��,�� @I�ҍu��P�~�� �9�O�ߘ,��fUk�)�$T�Qk���
n����� ��2+���rf����\�P���[jis�n��?��ο�
4�u�Ԇ5u�5h�B��q6$�@��D77�$(�I�3��������9U=QU�f	����*A�B1���,����J��',SW~�f�`�*��9S������8������{$�͇"!|�o�@N�:��)U0�/=/=;�0lk5օ8�k��kq��OP�c��Z�@X]��]��T�aPQ}�}"��>���_tdCYJ��}�e2�谜���y3z�jT�)Y������x����b��}���#q�?;��O�vG��>��u�O\l��)���7ܾ�
��C��FfD�� ���� ��X9��hI���8m�����1E�v��PЉH���9B��D?J���ƛ�S�7
�D����V�bƘ��|�P-��?��D�CO�����c��WvR8P�Ӎ'���#"���@�d�z���d�gTn���d�C��������io"��%ѭmnG�|#|�=Z�5��X�w��o~r
n�e�{98�aތ)�1l��<��o�Um��+����?Yt�P�pX��UhT�:U.FkW�x�F/����)��9t�ѕW��uk>񫀐C�ǿ�#B�;�4�;7��sP����D���'�v��6|��G�#ɥ�r_��WGJ�|g�=�+
�+���5304�8���
���Qʅ���HQʦ/Tw�����t��$���P��^����������ڨ~ѓ;W�{��1'���m�D�Xrpx.P�CY��Ë8y�P�k��7k�=b��P��KTQG5��ַ���Ů;	�y������t��־C��0}�"S7�ff>.
(o2�_Fd�������<�b������c�U��(�ⷊ��V�!1I �|1�l��^+��n�m���B��:�$o�S���6ϩ�;�=�S�mB�(����Dɥ�Ի�:#Q���Rz�����*�0��<f�P@��&�e���0���g:������|�������%�X�F%7>�7Qk�G�P�-f�L���jc�	h�6�jIF� :�n�����y��?d7����>����	��r�z��}�` .�٘M�5;�=wh<�)��x��/RJ�
!���'��4�ٞ��J���̵��bk�r�D,��BV$����(��&>xU���f��&:��͕�g!7�h]ďG�aE�0#�$���ʉ ��`�[s �ؕu(PKSE�PN�Ѻ��C�?�u����BU��p�BvvL���gǎ|ɫ�v(����.)W�zܨ���r�9\�2��V�,{ �0�P�xǜ>�=��W9ˏn>j���CU���|�D��o*�d�j	Hd��6�p��RC�g��_�BmW����R9u�0s��S���#�6�;ѽ�k�^3��q�ϕ�!*�����%�:�.����PT����j����q�R�1&�F02I�A~g�P���?9h-�.4G�������8ن���q\E��ӯ���ܢd���L�w���)���q�1�[��u��]>���x��7[��d���woh��iG���uF��M�P;�y����������Q�W"��;���Vl���?�%�������v�'M	[éјw��y�Y��UB�5*�v�M>���6�8o�ς�r�.���F��p�������Zek��ܐ-�"���c�X��Qi	q��Jy�?�=��6�i�Ih���]]���.�_��� V(��b�k���G��\�����Lt1n돣)�x�+(A�k���׵><OPqٜ�ߓ\S�G�2�V��Y�+�b�1�5?���QQ^�ǧL7�����L(h{���jEr"������8u03�����T�_�a�җ��t�I�h.҆ ip�D}X㟁<�Q�%aă��<�x�'7�O�w�u��]�K�/yO�.
�c���d��K���OPR��}L��M�����\����:B����9�����!��Ǫ ��Pz�C���7(a^v�-��<ch��
<غ
`�1P��ߪ����j�z����E=|�,��R�����G���{����ۗ(>9 ����F0BNvV>0yv��}�d��P0`�A��o�Fޙ��ے6�o����*�ǋ��CC�F90
2\hZU)�� �ٖ�q?���f|Ղ��z�K�������~�QD�,��.�Rv��m�.�y�`v��r����󹾖�������2����y>���ģ*oA�.Nv�*�R��Чhw|b9��|�U�q.�4��\��gɭ�d����Ra6��R4�!e,,��Ki��l��:�@-�y����lC�L��������H0>0-�0K����0� 
��e������x��0���o�,���!N��~5�ᚮ�]��+b��_�(�(��H��l=��S�uK�t���c��DF�YJ`���X]?�Z_4!�u�)"o^)���8��1��q�?䔯��v�Y'���*ş�~���}C���\)��I9C�C�8N��Rɫ/�8�k�L5=��֔����釳[_HA��S����#�vuң���~�Ϲ!��֬�R�$����OeȈ�R>����i�۬�~��m݈�v�L~X�i�d���JE��~/��inv���x�P�-�d��z`^=���Tl�L���4G7v_ݖ����I1��>Ԡ��r����7���+����(��RL�Բ�G���]%�c���{��]���o�����2�%�6�I|�YB3����n�sݼ�M%�ć&L
�?� 73�Q�L4 ;�-�tkt��U��d�f��
��R�F��YP06&��JL�eךٰ	:���-�?<R,�r�d���_=����;�����X�3���_ �G�+u���b����yn��9!V����v��a��q�`�-r���w`tJ�Ƞ�?����y W��vO��^�3�1_:��v�~m�}bfk���A�AS�nTC��:�F��1�+?#/p�]�Pn��+��yI�$�b������9ɸ�*������DI)�G.b0Rز�u��8�!V��W�s��m��_/�^[�,Vۯ��� MTL���	7�q����l���}�rC��/�~�B}��уp����#���܁Ë��W�����Z�v+�4c$�+����}8G�XacDa%�0"��x�T�c����6m�Y+��?�9�ʸ��66�2C�X��9��d�E�aQ��vO&5���g�Bi��}�Q�e�@�z,�1P�b�\��|A������9���i��'��?T��[��������� GZ]�`Z�Y"��Gy�8�Y�*V�&�f�, �#ݪ�7�km���u�'~��U��f��W�H/�$ck>�<W�j9[H�Ej����>D�K��()��k��^��Kp��C��߆�MHz�H�g���{��o�OH�vqe�[�F��2�4���]{�bI/0Β���I�+�op9sn�l[KE` �q�{���|���E���c���h�)0�LU��?J�%���D��S,�R�����1h�Շ>�f`8v߆�����u�B�O/��/n�&# �t�O�������,<��=��M�3�-7�O�r���	(Qū~T���)�Gn�KB�1�Hقͥ�A߂���	���Lp4���2����'�x���Rr���[dʹ)��O��^�8V�J�7'm�}�oӳ��M+6b"��~��o�ӹ��.�����k���du揁���[���7i���u8�F�Mn'(d����������FJ��SO��Z���f7�&o�1 �}����sH��֔Q^��^���!r�d��ܕT��hc;&��#�~���� ���{#I�{00J�W����#-µ!k���Bp���ơ2:��"+ɿ��IbƦ�Iy��b\�p��a)�p�/*�b�U�]�
�)�O�|�!�qB���[�F��un��k�G��R9٩f�X�7�������q
��ga�O��Xd��KU�a����5��#Zܺ�%���9v�dԠ��Y$T�k���A��+bm����}��o���k���B]���~ϖt:=ы8�q�r�N*E�ULv��%���
��P	�0~�d���Z�'��S�;�۞U_rhг���`�����r�=��[�>Q���ʎg�w~��Bx��z�y�|��/��,���A"Yo)�U� g��ӇẴ^��͞<0un"�@�@vT�:4���$�����f����q���:¦aL�vwA#�o��?z˻�vR�NkA��Ï�4���ݲ˞��az��?6�� 4�_d�r��$�n]�g���Y����r�:�p[���̞��� G��{����Yz���ll�����������������Ҹċ�Ѻ�����I/�� �*�:�ް[4/`��11H@I|5�R�a�1�(/
h����\)��ԕw4��:��������i����!i��K�ާÉ���)�]�*�P��8аg��������,"n��K�Y�J�~�L��Ln��S��I���K_������<���/�2+x�嚌!�(C���;�J�+Gi.�� �F�9��h����R\��M�����p�y�C1�ԋ�i���F�;�I��������Ogoo-R��fks����4���rP�l;5��14��g`�L��H��`k;��+���%�n]8���\�X�X�
���ĆQ-��T��	s�׮󅄸*�N�'��v�I�e�kE��)�VIRJ�;��	KƜzF6Ŵ���/�����%n�:��3Y��yRBv5󎅔o'-j/D��v�-@��	����$D�/��%�׉b��"b�]tJ��R����`d=8�]�i�?qV��M!YM;5�0�A���c�U@�-��R�So������^�N�=(���F_��/�$L ��a?N��?ã���|6j� ����!q��i���s"�޺q���^j�� 7S��)Rp��Q�۵��M�p��^�;\ ^A���I����M�Ab��I��,�$튠��C���%�9���s"��;KUJ��4�i��s�~C�X���ޔt�^�ɳ���6�}x��_��7h�v��u�&���0��G�\|V�<�v�T��@S����{�ϛ�� ;6&���m��
�&�Q��Co�b��@]�B>��A6��a��l毻��-PY#j:[6�)�8�#dA�'�O/B���;�W����M�d$t���ބ�so���1��FP�jL�>Ю�@u}�g�3*2*��x��>���F��+%��^���C5���z ���v8�tΠ��S?�7�����H��T}d��}D�up��Z��#Tp!B?�|[�I�@��$�^8�i�i��<b@�V�#�&7S�d_���K�M��L����a ���� f��͓6�x:�L�t�-.&4!��5؄pC�ӾQ��g{��Z��2Qչ_�v�:|�v�����1O���d8�W,�s�|k�6���,&ᣜd�'��������R���z�������)d�6�DsnP�`��h]@bJ7ߗ�V70��@�k���]ҴaXQ�R~z9gM�IO����Z1��YCC�����z�"�DY�R�DC�_�N<Jέ�vl��a����_��� >�Bdi���*M��6�;�I�y!>��JZy��!GΎ�H�ŝ�y�y7������-�@��>�p_�A���07v��d'�,�؉V���*[)x�/�a����wĂhυ�m�#(�8D�X�.k7�e����V���2t��k���hx�4	n@GD(wFUXmW\�7�����;�4J�p
G%!���߄�n3��l�FWH� ��.�e=�T��M�a�w+��e>ծ������땀���nꝆ�w�U���蟲��l���6>&�J��An�v+>����\<�ܦ�tsޘ�Av�~W!u�'g�D(_���X���jTV�\I�b��!4�x5��A�R�ni?% ��wB�p�M�k�Q�ك�h��܅b�P?M\�t����5C#ծn����齸^�evu�����4�p4Sr��I[��$/�����\WJ�!��)���Jb`ҡ'�
f�M����l�n����J�L�2�d^;J)�����.��M<��qTl��/��j�Cw4{��6dƗ�5.N
I	��B�d��!��,�N�Q�i�Ifp$Ӕ.g�W��mr��Z}w\'��%X�9RA�C��Dp�U;�!|~#�3��y�O�����N�p8Q~v���ԛ�/���u�b���% �_��5��#�;�A���T� ��
�6K�� �,\��b	&�G�0VI�,�����A6Lc�&�
�����cE@�)ؘa<h"���i�Je-�oֳ��^��z�'�� 7��}����#!ݰ^�30��ݤA��c��#�u,-T���\���[���Ǣi���L����V�c
�7�3Q)��k9��z"Kr���H��sx� �d����Q� ���S�S�qbR{�d(�����B���!jm��M���^���)��ǉ�s�~N��B��YTv�4���+��O�Κ�*��1BG����`��_�
��a���-ߖ���ļ��84�Ѷ�ү�������:��:%-����!S���A�n���1['�A3�����^S���Ű�,R�M�dX�6a�n����2��C`&�H,:3e���B@'f�쒜Z
τ[��ݚVUK��èJ��7�S����	�Ӏ��N)�dq����q,��vyB���㮔mh�Ra	;<*�� �dE���ҥ첝'�;�q��&D�xh����Dc�%I4G�uH&;L�N:�kb'��b�\9�����}�Q4��'���6=�D=��;���@VsP�J�0j�>Y�	e2���G�?V��ri}�0����a�_	I���O��n�1C�����Z�F=S�}/ݧ$���v��פר����b"[82z�ɕp�G��0\�Ee!�{���zʸS�q6�b���G����Wk�g�t��ɇ=7<qǱbx,����ƽ_LR��IY��J]�#=�5��gmKÙD��Hoɑ��9��ȭo�F[wb�'O}^�ʊ,��N=�˿�ש������#��i��@���o{�K��5���I�� �>�z���Q��~�/&�|=.�Fb�拤yQ�7z o��K ���8�����hX-;�eG�-)F���v/W2m��込�x��;v���y���z�s��+K�@���?��s����{U:^�$����v�o&h:!�>h��UV�b1��q����FIN�)~?v8m0�-I׭����Yx��-J��,�"RS�/ ��1Z�K�!�#�|7<;Y�	BS�8\8)���` �.X3�fX�3�6�<x#1��ƿ��8=��_M��y�y��|2K=Uo�y���b̀p�z��{q��P'aCeL!ǖ*R�.!��T�#��l#������U�ǩ�VOq��R�A;'�"/d�{��7$�*�*����/xⓉ����kt*M���������
Q�S�Kl�͕���SgB|�Nc�I�9�@F��Zn#�����`~��M���D�]©��|�����S�U�3����,@��Bt�;��DW�f�#6<xDi�LY�G�|EHI� �S�j1�	;�u����blg%�5��tA���:v���xu��J�S}Zu�Os���b��F�����h#$�/$>��g���9&3:�nF����xB��,E�d���!�#��V�;y��p�?"]?��oR-���X0��@����F�����Z�3��hdf�C���G��D0�ZI^��=��S��mr��(n,���I�'��X�XZmjQ64�{�`�����7���yâ�[�i4�5�z��ȃ!�3�Q��s��}�~v?(t8=םN��8�^�=����pw?f�tA��+����Ra_"�&�Nx,�6����T��S2ǮG#2��@��%�2��Ou�ʚ�-�m�\=dpvﭔ<����b��~����p�>�٭C�B��(&�vK�����v����p2p�|b�2Hhf0&C�,D_�K��)�̈́y�k�Ko�^P��3��$���d�8�8��0}]�Ӫ��O�4�O�����u]�[w����蹩�(�с[��EM�<�E��:;w���e�p������6�'��a���V��Q��W����PV��D��B�=�0��D� \<�h�k1N�����8����N{�G&⪻K��>-A ���)-��Lȱ(���B�2i�z�����M!�73{4�|���8�:�o�~�|i~<�Lj��͐9��q{e=��ѣ�%�/b�H�=��k��d�[���#R���Yg�שS#�\TԀ����:�WC\���D�Rx�DlB����?���z����/�X��v_���@x^�/�)���k�Ha�T�Ȧ\�4ӾE�
_J��KY��4�Qϯ*�0?Ɛo��d�Îch�5ȕ�*'R�'�
�0ށ��P�4����	�<���������S�����P����q�X7�j��G&��B3��|��@��
���аE����Px3%ɕ�g��G~��H3a?�MHx�����i�5VR�El7+�=x���-6�n�z�>}��N��������q���þ��~���3�\����C���H|���vj�R��Y�9�C������4M�*��ȳ(M��4�vk�^�n�b:'ٸBNq��+b��"�>�G~=}}�oC.�~�+d޿g�#�t����R�X�2l�v.
��d�!�q��cjߌ����\L���-����"���\T*�)`22��*�F�C������G)��i��C���:Um�z̔9����
4���8�9���2�/av�i!%/�(�Τs�T� �����O����!T�4��P@� ATi��g1I�G]zh��[N?���U�9��-��hF���$_|b<����#���GBk=����n�3�!���u�<7��,�0���_������v��� τ5��:��=E4��#
���4��!��[~�i��t[ϕu��酪��HI�[�H:[�AT3;�%�;��ƱF^W�c\��.V�����g���R(�o���X�%z�p��~$%G��qM�N:�YkE��HE��*8�Թs���F���x�#�9��8�@�\5���eB;hۮ������'2�i"�7���OO�xky��I{�uG���	�V�L(�N����p����4���t|C�3�,Ay�N;����p~�X;q��/JpG^I�'I�Y���`�{3Rh�J���p�/-��x3b�v�y����WĘ��3��-$օ$F�kti�t� �D����mvZ���b��e`+����vc�� �h���H�|����Kk�i�M���z�`>��&8�P��a���_F�Jp2��u>l����|���b.�)��O�Y(����먃�_�h��HgEO������K��lǽ1/����Cm?#kϠj�� �܉�uG��z���:S�f}V?E7�Q]���#d�H�^���6A��7����]�	�S�!Jg
�IN�p�F����f��9���*��D�_ `���z�����r�e,���F�/dr�v��Q���$����Lz��8�h<QL%x�l<kfB!�~�>�R���}��u)���o4=)zi�� ��Rw�?NY�	���ro���b����0����7�z7�;'VDZ7\TQZ'?FF$�&6-��>Hy%>�IZfx���N�ħ
����⽽y�ɥOB�'����/I���>i��o������_�O�}�s���L<� �x�m� nEf����몡	*�2��HN�-�#�ĸ��9b�	L��eFz:���r��1G��8�x8MI���pG8��x�8�'�i���$Ǆ���1(	Ԋ�(~����B+|�!��X}#����
u\��4j��">��J�:��(����S��Eq?0�k�d�oɕ�e����]��)�����������uR�4 ���{"J�Y�+�cQ\tC�ˑY	�Otb���O��ig��a��3*��~�J��:@�{r��d��r" ��N��[�,�UF�����Y��1�b@��'��@J�2�9��<{^z?��u�n�ֻ�����C8�����}��8��Ӎ	��hk��|�zC�rX8G��)�~.{Z�ӱl��. 7��yQ�9<��&yx0����n�|�� �W�|ݬ\Η�$2�՚f|�_|?��ت��CTe�NCUY��������wմ7�4M�2f�)�|e�d}P�!o��օ0���8��N�v��N�����"B�Y���R��0-|5G0r��`���F]��l��&��������v\��I�vc�&�MO�r��04����PxP)�Ѕ�
�Atb��v��Hr�֨x�;�&�B��ˁ^u�����k�j���J%� |*H:v�=tu���!�����Ye���F�}-����+�4'���^����c����"�)�]��I!���~��VT�H&�C{��H��Jz�r�#��&�"��Z�����Xlۑ�6�`��Ӣk�[D�5J&>Cr���[d$;H�P����1>&��b�|b[���J�a��ЊB����� A���ݙS�U>���4����<���'�-���ڰm�,4�|�w�jR�B3�`]��0�L�	|:�#%[������).�i���{�*i�H�%���͞8o9�����I�p{އSv����pX����C�;0g�v]��m[۶m۶�c��m�vǶ�t4���L�?�u��ԹG=������e��zR)KE"W#�~��8��hR�e�$*
<�}��*��~N��w�o���XW�?ӱ��m�]�X�]��,Ă6ؙ<Aj�#5�� �/�f�g�n4{7kC����M �E�kGJw#�*�-j]2��lmǻ.F����j"�{J��ҩ�i7�D,����.�8^��=l�����a��� ���/�� �)*6��L� n%�0������e��q@�Vz����	'Xh���@�0������L��:�(1�+IHE�ӌ>��F��gbeXbH��Z^��a��\�����N�0(�(�*%&V�riK��8�UF�O"��I3�i���\&�c��� hn	�K4Aa��6���äO�J���7}�q�[���|�>o�����Ϧ�V����"PG)r��ٙ�.��&Y�q�u�]*���en���x�"�ê){Xݔ�8l�H�"���SVXvʪ����"���<��x޻�:���� �ѩ<d1?|���|� ����l����7��Ct��<7��W�8\ڶtKj]���'�/Ѫ�Pz]���2O	j8uh� [/d왙c(8�w��$���6N ���TgA�,l���K��E�`r>�w8��1G�����*2�_B���g��$��h/v������)5��lY�&?�>�s�~�*�����.Ϗ�@D���&ʼ�!x���ڨ��K�����/,��!Lw��|i(�?��账̇'v��$��e�9"�Y4�ah��_E�"Ē�TVY���7Ձ-S͟]1����Pi���R$Q=�Ttj��!�y��B��lp�E���Wp�
���A�V�ի��Y���� �@ʺ�!�R!h�B����T%��`�t-w�%��+X2����\�4��s�ڜ��C����*Ø�P	� SX�&c��8�.�4hl}o�*�F�]�!?B��!e>��:��v�]�ԋ�0�´�gs�Y�zD������y�ߎu�Qy5�����w3����H�n���Tn_��#�!C�rӵ����.��䖂����6�Wb�����g��'��p���5�`^�bJ�J?!m\u���	^wL��Il�m�,N\���뽈����]����W��¸��@�����[��@`}�ʸ"��g�Ng�����8�$-i�o��[(��H{jrW{Ћ�c�o�Y۝N�"�&���y�ʪ�������	42���*4�h,�a��K�� �5�#�Yw���Dl]��I>�6�?�I1��b�7�e�6Z��Wj}5�-zh��N=B�9+	\&��\�+B{��n�e`���7l�8�oش.F0!�\���c:�EG�p�� ��GZ��4L0;��\^~�M���73�Ϊ�9���ȿ��'������:v~>e��i�T��Y�?UN2��a�s��;�̝��\L�[;'�O$<�h��,�G�o�>x�׭ֽ'�m�pD�DB��ՙ���!k�a�{�l�a�5��	n����<q�)�sQN*^� �`�j�I�^�E�c
x{ͤ��k[�����*�p�+Nl	f�+`�����f���Q@@0�|�
=�|6G��Ҝk6�jE��1�8%��N�t?�0�]�S��_µH��7�uD�DVF�S�Xz��	�6��I-'�X74(p? A��P�8��u!:Heٙ��_�a�\ s��1�ge�:U�����KW�*����C��as��� �w�b�1Ņ*4�c�^-VFf��;����7�!���>靄Q���ҍ�̆��FĿ+(�f�8�N�G��ag�G���%~��X��!��>���:�D�kh��=�iB�]��wD�Q��ǥ�Џl/%�ǹ��?�F�B��G/����4KD=��Ӗ#Ua:�0:V�
#��K~S���6�j��֠XO.��6D��| ���ɬ�^�ufJ*�ɂ A.2�H������Ii�M<5�$�n� �0Vzм+��&ѝsFII��b��.��ߨ6Hex\�1��Ϣ�~^�uTq_y�:�=W��\G���T�m��朴�g~a��jЮh��R��v���H`�u�=��3�{�<�]��L^/�.x6E��6l-t+���ʔ�+�T5v�s�<��R\�E�)	�
Ov}e���8���J��+�<
�;D�6�|n �lfQZpD\��K̖����.3IW��	w�-`��/��n�v:�����͜9er�3�+�C�v�3jɡ�T��㟅y ���ZJ��	X/8/(U�4���G��2y�ɥ4q�=p,��`��}MW���Gp{T|���X�:}mz���h
s2����Dwc���+�B'I��Ppl��AȚ#s:
������Z��fH�R8d�~���S�j��2N�6��"���D��%6t���a����	M���(�I��x�UU�Q1#A@4��ם�
Uf��&�Yz���?Z`w�'LAG
b$'���i��/���mʱ���X�drtτ}?���R�ո$���ὭP��dL�bm[C�4[Q���&<�Z�0zt�����c>��a���?[�!w��ਫt��J�b��¨=�e�l�E���1�0��N@"Q�j�iG:U�h2ĜW
���֊�4ݶ���4�b�-{���|˴Ż��Y��+� 9�Q�>�����C淏]3#E陽w�F)�cH]%�����&R1���U�F�`�.n�!�1f�$�D[��i?g���k���J�5\'���X?@P�<�vP��fܑ�,����,(Nln^y��?��Θ!����J�G��h;:���M�l.|�\���-�cBpl��^}^��5�847	�����0B���7�VTC��G
�5��%��^�������Խ����Y�(#�^��DEdU0�Դ����PK��"��0[�\��d���$�� ���L&Z<��IA�&6e��4bP����W��/*����V���g��"��sx"��-��c����j��q�,DL�`�'�k���[O�#��jf����ǣ9 t֖*�-��䴕�H���L�o5�N����.�X��f�	�#��E�Y�r�^ɭ�����|�9�TB���~`z���=	̅(�_,�<�Z��؃3w$�,���l�����>SZSBj��2#B���*��h�k6)`[R��,?;d��`���2V���%&Y1�y��pAp�����H\���M��)������֌$�PϤ��o�Z�{]\Om�|���HJ�X<����٭��������"��>5ST��V��Q\����L�!j��Ʉ�Y�O�Rb�˗:<�9���c����~��h��ȋS���.C�[	B��
1�]%Fhe�k�H�
ۛV	�-Z��C�y�
JV�~_�k~���[߁ɧ�`RN�T�rÙ�y��;y��,vz9��������k;I�3�x!~��d���V�6��Nˠ��|�c���V��
IuƔ��e���k5& �%��M"rC$���yA�G���t�������Q/>�l���C�'��L�GR��r�c-A(��>��	l�?UkvwcU|���":%��%���{�*E��^�5jGJD��C���4|�;�Y.��H�ԛ��9}�3QxP0mQ�P�`��1^����z����&�C���P��b��\0$����-.쨁x�5�sE�ҐXh4��flm�Yd�s-��g7�~D� �F�2G�W�8�(��D�B��I�"i)\7Y� g;���-5Z��?�����@()���'}�q�"�����2u�l	�8-�~�������5�Ә��/B�l�LN`���e��1����|޵�S[� xH(P���յDn�F�d��BYBv-*�Sj�o���^���fs��@Kq2��H��b���I9�}� �����@�b�$D��$������mM�A�L���P HkX�̕r�z]��0�h�
*#�ʔ�霞��%�4�Gմ2�� k�_C7�nB��)�J������@J�^�l�C�c�hoGFa<OW�N�ǀ�S^� �:�P�%n!/��iep#L�E�V;�#�b6���ǥG��	���$�+aq&$G��e����!\��u{�A��Z�1/����r���R�o���\��o��,
��.�~n{�f�|����uRZ ���=�;0܃H�SQD��S�wMR���>0�wL*k�봚E9+��"���2:��g'2	�h��>ݺ^=��N��W���ȿ]ƫ����+�x�[�a�.���v�V��v��3��R�W��d��꜔���nI��#��9I{�>B������]��º�G%��U��e@:$y5jrk3R5\]H]AKlki��?)�Z��rS١ĕ �7j���$Z�tm;Xcx���z����Vo�B	G��>I�A\�^c���꒝�'G��H�NxN�OUڜ^o���Y�46p����)񲽚S�=E[L�Ӊ�{�t4�
[P3	.u�دO��W�C)멳E{e3�����������^$��
��q*V���UB?��%�tVw�t��"q���NK�V�U��l�Q��;�:���#M�Yn��K��Y�vŗk�� ��)����d(����X��6��Q���u6?���,�h�+g�٢FȔn�!41�T��YW�v����)Mz�^͂7��wl���t���>��պ�4�Xn�"ٯ�p�U��C\&�ZU=���]�^�ިF7{�r:-��Mvk�S>��aR튰V���s�V�ӄ�*�/=6��]�OԢ��O63�]���K�Mg�<� �%�ы�Wj��o�(h\��U�2T���'�(�������pΊ��)�R|��9�:Ḧ�g������:��;�{�����A���L�-i����q�ElZy6T!l���{�W2ѧ;܌��;�d�r�E��Vq���;�
�P=�^B}2�����x�n��U�N �M��n��o��񥜈Ȋ\i��J���4K�P�(�,�)k�ZB�Uq�K/ ����>�o!��5��\_D㲍OH�G���ξ�c!�o�QO�+s� ����h�w��j39;��װ�Ųgש��*7�o��y(���g�������f.o�7������B��~7�(˻�o+�$������������3ES$�ER����mQ�SPȯjQ;_�J��Q������B� ��DAsq�v���T��%�a����Ɋ�O?<���N�U�&�V�_
��tu�P��V+�>����U��[I�8~ �T���n0�-��EQNN�FS�\�����
�
�]���)O��E�t���v�͙t	�~]ȻB����bі��#Y3&�O��|��ʾ��'w)[5YKu�w��Le�Z����E���f���L2̸їҦV����T�,���CO~�����YDد�ݜ�2�5@(��ګU,�R�M>5�����%�������E�(���A`�����}�D�m�����;E���<��j{l\N���)y�N�Ν��Xu���n�8s�]W�ԥ͉5���0��-y�!���у�x�=�.yZa��pzfdx?Ty�9ZcB`��Hw� `Pf���E���ܚl,`�3��&G��$��I�ʔ/u\9JUWdj�a�~*�`a�;|�D �5�?� 
mJΧg%R�<�[�l.`f���G3�KF헺�r�*����_�ey�/8;g<6��c;0� "��C�9�n��D�H�eA*'�O�.FU�
9�ӢƖ�N�P�j�FE���!�����["qC�3j�����ӇC^6���jW��қ����g@�Y�]w����_P����o�`ˆ?�2�0�������^5R
�O�|��@�����t���2����G����*C���Bw�A^gp���b���
\h��e�H;1|��j�2r��豘?:5ա�oޕ#JlC�D�_Žu�����k<��q��k���U�3Љ�x�	>���5�*9�P󾅜�cVq�+E��l��2�{e�ZUb�ϳ2ٗ�9�M-z*�JG'qh\�v�5�B�-xc�'Ч3Vf���fm��O�{���f��mp��aQ��ԏl-�$������w|:�V��9�����ի)����	��|�>�Y�-4�EQ��F���)�i��#� ��ip� ���qBu ��55���&�FM�I����"�f>���, H�L�O\��fz�՞ӗIEǭ��wu �dj�Tv,�,�j^׶Z�
�"j���T�hg�R�R�W�N!T&�b��!�/�24��@D��~^��('B���i��6�wH�z������z:K�	��=�^Ō����n��泏q
�-EC,4����`˚`5zu�+���/x�����3-��`��->� d�����[�{t+�]�8W��9
 lT��nSǘ1�p��N��;XM��!6F�����+����aSJ9���n�cY�܆ˊX/�Ɩ����۳.g3q*���gA>lq��͑�.ven)]D��ײ���-[|�8�Nn�C�gM��+6�9�>ҭ�,��V�ʹܯ�Yy=�˱�.<�Cޟ݄���]��LS�W[ZM�N��n���c�,��p-kH'�U �	PX��Ď�r�"��-���6T���
b�L�Y�c���u�F%��vҜ�C��R|��0���	�X~��ޠ�0�����rj#�!��,[q��D�=��+GN�����M`�l6U2+�b�27'��	1j�v���8]�i@�>��y�� H$�/$n��zd˔�D烈��k�r0�Μ� x&j�[HH�Y���V��פ�C�;��Y>���Iy
t2�sS������������6�M�gy���@8�G���?d����* ƾQj8~y�����7bE}��:�U�>Q���B�a��ן�:���;��-
� �&L�O��(/��z]5|�]�g�D��U"�5�vǿ���HǊ=���
>Gy@���o���������к^Im6�hw�kg�.|����������w
]OOT[��`�-q��W�n6��!�v��Ќ�� d9Q2�k8@���lC�H(�>c�N!��᠉:ZS����u���?eq;Ϥ�B`��߼�/`�VoI�x����RpkL����.�'?т[�G��F;��s)X[}˙jˬ0�ԯ�|(^g���f[���$^Q�K���x�KV�̓/N���ᩊ1�<z�h�j�"��F!�<x�R�):�}4;���w,i}�=�S�u����}?�ckٷN��eYH����'Id�ˌD|3|�48�����z��K��u(�����|R���R'��D��]fl-�`l)��|L�I�:���\�g�ɳ9L����zJJ��!AqG$ܤ��ޛH:�Bգ��o��:_U�G�r��0���a��&G��$��f�\A��z�L��VE��e(�V:ZDʸUCՕ�y a�i�)Œ"�C��*����1�5V��~��i_�C/��:�x���P+y��ҢT{�9�RA�g��]X�`�F��dg_����B{���aϚ=Q�d��o���bH&��/rkh�X#	f֦�N��6[����ݓ9���<[Z㾌��y�u�T�؟��;Q�F�.�gBo0�W�܌�c��lhqv��[؄�'�	G����emW{�Q�q�R	�W�>W���\�<�3ҩ �@������s�0q�"m�SV�N����Q��a�������FL-7��t�9��U!�Y|Cm�����x�t��.���t��B���9�=/�K�JR�d�(��[��G;�0�ͪ�Uܮ܎��%�s��Exi�1�@]��[����/Hs@F�b.*R���*�k׷���ǂ�:''�r1-�i��?�翎ܥ�l�%׈E�l��+6]ݧ��Ɨ��U�*�0�������p����$��yV'�������>��>�ZT���P�ƍ*.����T�ښz��L:���O^C���x�_e~R�F�4v)'I�@��D�d0ӳXZ��Rj*�����f6ڲ�RE,�^�&�����)��+���)�]-pUYe����rӤ�f-���>�Z���5�2j7��SE,���'��E���(Dc^n���m�3ў�SI���^�Q_�g<M<f��t�&w�g��&5�C�#ʭ�-me#�OlV�=��3��T��Q0�r�6�57�7�M~d��50��Q�_��ŘUӱ�]��U��E���v���o�d�b��h`\������VX��M��M%���_^��KXG$〻��5H��-���;m����k��MT<�8�:��e�[2�?� �_\}�ڭ�،�>����P��j�c�o:u2��t�vd�AF�<��B5�C�DB�z�9��-|�����Fu����E����EO�^?����q2�B�eč���M�j�|j�	�.&��|�E�ɇ��a���i�����>�/wS��Ԭ�>6ipzgJ?�O���ܣ��I9�[��c�&ƪ�C���7�������ԕ�U�q��=��l`w�oj�K[ ӊq�F>j��d��E|>w �j�3]�O�Q������<�eW��e����f]�C͑��f����'��g���"5_I|5�)7�H�,��r��=��/�c�vS�ٹ?�¶��`�'z�b@_]�sR�FK�JgR��+r�9-�搾�K����0a��Y۠	�[N*�?�m����_si6�]����/:MVj�hD��+{�g����Di m��f��������u���F�Iӆ�������䉅}@�W�"�UX0��Ƨ��ގ;���ףF_&}��5||��Nc�N�B��*�dk+�q����4a$O̪�7o���Jaq�����ä|���KvZTXb'���Cj <>�rM9����D�!`xd�K�����(�Rɳ8H�H� �2�����V(�}¦4��G�@���6s�ϥ(I%��&�f)��)B��%�Zq������6�'�|#�G�#k��pGa�2i���c4���_Jl���M�h:��p�xmnَ��3�*T%�e'��µ_�4r�<�Ci���^v �Ơ��O�*	$��z���'��V��[�ϯ�h}U�~L�����<�{��^�y=��� t�D��s���~�+a�3�W��A�m(���T�N������UM{:3Sr7� \D
��e�1��@�ѽ�Ǻ����o\M��71����ք�gϥ��g�ҵ�Ճs�s	�N�5��'��vwݯ�AJ���L89�˔F�S�m5�Q|�5�Tk9�Ät�c�ΐ߽�u-j�+RYpr4�d�V���F�E��>L��h�#[��!�ڒ�;vl�s�I3�t�f��g�����c� ��؃+�����[~*'�""!W�MrF�E�\mtO&��J%��@�g*/��F�0�S�]�
t惋i��QTH�]O��b��o��f�07�G����M�����A�Qto�L�h��nkӪ� 2r�����?�u�!O�9�w��2�A��(2Yw���K'p���#7֜��
k{-��#V3�:B)�T�jr�9����LUF�n}�����̠	U����o �£2�D���/}�1g���	�2$�4��c��+1R�*�)O�~⥆�#JvF��亸Y�m�����j����>�.�Wn�}���+p��@l\�	f�L����C�}����X����~J=A�E~nʏ�U�O���.�/-�}2�D1p��R/^���J)\+qT�0f�5���'6De^��^f�H��~�C&Q_���Ԥ�2��t��Wú��.i¡�z�0��Vc�s���)A����|P��\V��%�R�R&IPW�B{��%U��I�m5������l^V�)��u�H�y�||؟������\ۺ:H��yBI�WBS{�L�u���֗$7�|'*���\�x��٭Q�jp>1�E�م�X�U��E�@bIe��e ۟m����研h��,cƩ�(�zey���?e�G�C(��3z�ҵ��]���x�[�+���ֈs�zR�Ƚ�*��Y'0W��|뇠^f�t�{p<8���J�\����>^P�@��d�?�� �l�.=�o��|촄7�S�1	��ש��e�D=�'�)r�m�m��輊B^{�Q銲y��[���ɸS��@XY�(��� LEؠꄝإ�J&H��4u���(u� c��θ�&ä�\ɖ_��H	lAV�f;"�����<Nz^q�LP�����7GLc����Ky��g�f��^��������֪3�f+�q\Y��y-|(--�K�lUix�����Z5��+���D��_V`�EAIc�{g�k��}bu�{^���e�ª۩���yt�͒��w�,�9T�f�zJ�0@[VQ�&4ns��kӐD�.2b�
A��*=h�n�YFL܈Q,��7�>v.�rS򑵊z��(ܒW�{�j�2��Z�����o�(��t�!����^+�MgԢӭqM��v��gm��6���JS%�F3�R	����H{�;���6���J�'3~���j����I�����#C��+@�'p�j�������oE5�`^���~>�Q;\-��	�`F����|�(��N�aN[I�
��a�y4�[t�[�����+P6�&f�';��j8��aJ�T���N;�0e����XE������^تe��,���dȅ��0�d淞s�q��<�o�hU#�٘�O�(X}܏7���:=�4�+oR�J�E@u��MG]���ߕ�'1]�^�o���x���	�0nx{өk���RHL��	}�#���vZAB?�����z�!��ٵiV0R�,'A}�S�nY(~���6P�"5�F��؁��p��Z���;횺�7`	*�w��Aπ��-'Z������\�x�k���Bm��W�� �����ۼ�x 5T��Լ�^����I}F��*�qn�tA���Wڗ;������v��m[�|"��fP�R\?t(�G���G,6�PD<����|=����I��g���4�l�pY�p�-Ѥ	��\���x�<�Yv�0ܤz����7�Oo�	�bp�^R�D�s:�[�O�h^ˌ>���[���d�	�c�8�o�7�>yi��/�M|x8�%u������ٴ4=��3��P��q
�pP=�Y����܉��)rqFK�,�E�hh2'{�	V�%�p.��.4���a��Hț�6���������j�.�ln �"��oxg�����I����z���r�Y��/����`� �Nن���zu3%	Jt����rg�F���F��`�g�觑)l�8r�='�'Lک��.� ��Rj����un8�-�sU<>�O�G����݈kЭvj׆��4����i)�M0�]��P������v"]4|W)������j]�ة�A�[r��8� �OTfq�����-��[E�����ܠ�
�h��]���~Rl`�����[�M�oje�����<����|ZX����%)G�����z�YXHd~�w{���_�)����d1�С%�Ծ����Q5�̪��u� I�������琎&*pXf��Rr�0�8�wF>y�h?�x�9^�`@��K&Y���,=�%�;��_ϛ4�
S�	�[ˉ3��r0�����`
Гۧ�<�ڍ�ݢ�Av4)-�.����ζT�����ɋ�_�݁C"A[[9�C�~��U��/֐�h�*�ST��r�E�f��P�OQR^7OB%���i32�J vq-���7�'�l�l�,��������Af���'C{F��*G����..;��u�c���=�5f�fMt�b��g��=�Q��Yw�S�Î��uӊ���Nar��&�-�V	3�<� �����;5�̈���^�'�Ϊ�=k$ʻ*͉�w�B�?��G.g��w������{	ab���Q��D/�8�{��t;�9_Ҫ�L�z\q�0>0(�y��QX��0�E��Լ���}����2^� ���hՁ�H]���9� fK�o�2T��o$����(�Õ#:�9�,��k�8�뎕�/��Tvs���g�C�VZY�0
�6� �t���SR���,��o��/?��Y6�p.�u�$�R��	)f��	��V0	> ����b�� �Â���>���/�"������8��LƜ�s��ڊorR��l&(r'�64YU�c��0c�93QV�m�xi���46�nk�U'r!��|x"L������7x�ލbw%iL���Ő�8��ɀ�rr�ۅZ^l^�+�D�xp��ct�DC������
�C�t��Cf:�%	J�)9�43&�l�����ܽW�Z���(��J*$$ �����ŨG*EǊ�%��:�c�z��wZȮD<w�#|]I�/_�:�ͪ��0݆K��X��ߟ��s����d�5�M�]5K�̺ΌET��(��]���a��6�|��0n��S��+j�����{s�Ю�f�qm%��%}��Pf)��zP���ԁ�1ȱ�-@
�cN�i�o <�ZoL#�p��\��R�>]fb�S��c� muzˌ�l��t�M���]�Y-i-w��9�;�Oo�Y���J �6@�s�۹�c�k��?��5��E��"W�t�+k��?_�wh9������0��w�������fT�C�c`%�?���M�oH� F�u;;�M�Xj#,f��o1w-F�k$��h�o�͒��a�ɯ�\Ą{�B��i��6�`��{��}0�cCn��]��7�OȎNn}?.�'*Z��¯Ĵm{vrLM=���e�ޏ�2۷�3�T���U��n�X�#FM�x�uSb�(͊4�b�7u֤ h�]rc�s�K4X?X����?	�Y��yÝ꼶�����i��FS���E��0���=�5��;�Ho%�@�R�?��~br�[&�v*�ʸ�m3�]�ۆ���R�Lk��OOt�%�I[<6r9��"j����،�!�:��i�����j�TX�3�p�����.s���������Eo#%<��Vs�N�R�c%��>��.�՛k'�_2�`�|����d#̅�[�xWK�rf�q�����`��3�MLG�;�ɔ��<3��� ȗ�P����?���{L5Q ��AS!>)��h�^�*���J�@KiK���D����o� ��4*�4(��Z$LIR���n/���VJx���U��G>mI�T�<<4��Uᐛ�<��&����b̓�Tv��$'5��^���u���5D�iO(�뀜b��$����Mx<�����tq+���Z���Hd�ܤ�A4!�����*I��n����X|�e��;�.M��|0ΩZ���u{�_iX8��Xu���ko���[mnǰ��`	r��O�+�-5b��Ǧ�z$b���J��YI����,Z.�Û��i�����@͆4r��_�q�������I�+V��ړ���V#�녇(Y�D��Z���{E M�o^D���\B+�6���!�5:1�OYD��b���B�>ȪFG4�ѽI�U���ݹ���H���.F܀�	XXo�o�] 7@�x����o�#d�|>�_����M"����� �j�Ҏ���Ó���S����8>�a��n-~�T3%����=<�7�Cƺ'KY�y!�W
��2���d���]N�Q���f���E1���T%��O�~V ����S�4�
�Tu9�h��&�M��%��Z3�Y�����-_�g5�!�L���ƙ� �X|mH�l�l����ݟ'_)����^����<p�;������[
�����q{������ϓI���1du���,�E2��Do����u��L���ime�5fc!�F����!.���؇U�>�0ԻM����v�5�u��:~�9|�qR��5՞��PBi�O�	�]��`6�ߒ�8���B��)z<U.��К�5Ԛ8�]����N͌�IU��ń�},�P�����z;��h������ZNL�9w+����q�vc��m�VEb	:��c�����}]���v"�p!�P&��S��L�n��WydŎc�=+z�Dщ	!�C�h�V�����1�4i��M�q�ߌ�.q�[-�#��w>j��,��M���Չp�*pP�!�*V�H�rҦn�Kլ �Ǌ�J�x��'�-zpp�%;���{{���V�+�8��$�J�ޞ3�A��Ζ��߮0�0��2q>"dtVi~CQ���(�kںvΨX5��
�I��ڡ��d��*t�(^��wt���)��~��?� �m?�?���Sj�M���t�����l���%�	�'�@6����c�M�81���鮁�a��t4�U=! :U��FEy��$�0@��n��K�ϣ�H��#��	\�N����||�g�t*��V�*b�C7��2�S٩¨��|�(6⨋��qKj�B��39�؎q�KV�(,���a1c��Tm��^PW�H+_�"�g�5*�/ɨg�C�bo����	�ɥt�����ŕ��������'Զ���.=YW��Dx�ވ��x ����W�hX $o���.�p��9�m�$Ԫ8a�h*%9KmuQ��&���aP�ש���s�&����87������W?.�i����r��{YL��o���`�q1���3m٫��
�\r�dJ��i)��xȀ�K�'O�!�ި��|�qG;5���Gk"�q+e�!��AɈ���X�W�b����Gg�ґA/�nO}vv3T��)\�^�"��KѮm)U�-���;X� �:�9��>c6�'��~��W�OA��@��%�#���_���W��W2$��Y��4?���/fk��SX{��X����%���ө���e6@�N���j���F�,s��h}D�:z0�
��Y��%l��;nd:md�RS�.9���v��P�2�r���4V��R��)�x�?Oy�y��b,"B^��وEr8���0j]t���'�YޫT2�^9pÄH�dxپ�o�W�"�j��e�ƿq���Q���x��f����I�g��NXNf1��Ⲵ�%Q�˕b�3�CR%! ��2}��ｆ��*�Y #�j�y��HT�ב�$�n)��������hԏl���l�Y�dF����x��.Z��=D)\tuC�t�z�R��bPP�u=��	����_79L�.�-t|��j��l"y�)O�5��[yV�[�s��e�z�`;c�S�K�H���+��D�ll��^����AV����5(���,Z`�j�uۼ1W��t�<k�K�@��@�(���yɉљa�nǇ=
���ԌTqS�$��֙�d]�~������똂�!]p\G�b�%�4b��|x9kz;�	�&���R�R<㘔i��$�p;���	��gx�~��<���0E��
f��=�bn~�nHs�	:+���$�'Ėk�����;.îy5���ݭ�,�o9�%�XGl�rk�x�%�)K(�}�R��G ��.��;WਭS����>����jz1]��K"���HS�9�<����W�*k��-hj���z�m�i��	�e~&4��^���,JQU>P��Kc]����X����LpzT����fMi���������W��� ג�m�tc��K�T�AҰj�`��չn�S� �����󫥦��6-������ݤ�7ğD�����{�1��3�{�V�;���T5�I~�h��8�k{��A%����%��t��+�t_��B_w����zl��=i����}���h��w�ǋ�#�%k�o�0O�scН2č�yb$�"��Qz��,�����9iW{��x,�K�h��>"+����64�(��ɪ��5i���S�!�+����[f��f�K�7l�S�̷�X��P�D"X�Y�y ��ؼ؟�����Ѳ�����(�s�s͆D.�L�`��M}u�*2,%�.��5W��� �f�q�%�n�]A��4f����|gL<�'��|�ꂿ�������Ű�ؤݢKwoۢG-��C����ڠ��SaDJ�N�����`
]��>�Fӄ�*��%��7�Q�<�vk7�'��.4��r���@0R�W�x5}6I�#fO��Ќ����oz�$��^��^���}S./$��Q>ٳ\�2�N´��{|U�;zzm�l	�)�u�O�<i6���RM�(T�3^/�e�1)�
 �/�W�}��/�	����<?u9tg���v�H�G��vI���xAx�@�x�e�|�0P�d}�M{�Êk���B�)��A�����^D��E����O����7�W�5�ƙxb۶5I&�ضm�ض����ضm��y�;�\����f=O���nq�����vES�C����j��>z���62�a�>������)��c�nO�-;9f.�x��Fv�J���Ɂ���$.���,��/�P�!'d���(Y�iܗ�P�g2�7�?�l�cVRd�.oѮ�c_�A/�.��C��ɛ��:���F�u���6�?���o���}�	�']����F��=��σ]��,0�_��p�r�R����P�k��?r�=����������qY{��)nv��.|��(��u�:���I��~�k����:�;��%&8�5�4�|�t��!�b趸I�Yz�ui"]>_�8ķ\ h�L �uر�l�t����io���=_ڒ�.x��ŕ�lqM�'{��)ɿrl�b�{aX��	�|z�p�x�꘷)����E�V��a���d%)Ӝ\7g���+�G<KR}c���b��7F�v��E���NU�6��p��������v�"q�{�#�/sP��u��'�v��5bI�pAkUS'}�RY�j=��''��#q�x��]�#�� Ӵ�HB�0���Lw���yÇ���h;.�=�����/�$v�i\�ě;b��
m-��x�cxՑ���x/nz�v���O�Vmrx�@}�B�rth��̦j	aQobQt?'L5n�Ck:���i��XS�S�4�_F� ����a���I�A'�����l�^�Lq�./HD���v�&=�?�*x����b�^���	]c�jԿ_�J�j�h3Z�٣Z����~t:�b�G::,C:&_3�@�P�-�v35�U�4�����lp������F��������#uu�h%�DK������M�=v�!��E9f���ɍ��ܺ���~�������]έ=J6F�����F���;<�[w#o�~�_6�w��458�S�$:����R�r�������vX�"�U�p����6<�?�顈1�!���&��'�EZ2h��30�~]q�4�UC���86VE�ʺd�B)&垦�[� ���$;�
i|8ěMC\{�&I;2ց��v~ hl�Hm�BmdD�3�K��֑�Dյ�HcZ�male:�='��Q��4�^����__T6�z@+1���걓�� �}>;�ܽSG!��<"�~�з�Ň��x��%��z�9��%��T�����n��[w�]u<�<�C�,�<>Dk��h缢E,oB��Bm�g��Y���`��_,!��^?��~�3[��d��PYMI>�H�����^���w����
� ċC���|�d��)�#6Du�aJ���1,ְ:�y�@���y�`ZstD���E�'a_R6��R,(7JF��f�����s��hG��H_a\O�j�#C��0F���v�L,�"��қ�s���Xu�D��Վ�0�;�io�|�ޤ|�G$����婯�����*����$
�$�ʢ0	�>@�gQm����?�Y��*���~ĂZ��Ÿ�^�k!0��2t�tM�
��A��W�䏚~UӁ�6�.Et�?+d�m�l�����@C�J��{>hP�Ύ�`�P�0W$"��Nf��Y���Ubq3F{?��x�-�8�v���nu���,��埾��?���E\h�Xz��r
p�Z�m����t	����x�f�^5.ni[hw(|�?&/lض�T�R�����(�^��.z�1�nz�����Bd1|��qBt[c��=���\�

ؓ��|[�	�����e��5s	��ԇ�����!:���+x�㨷�m��>̛���(<[͹��N��&�X�Dj#{�E���=�Q���퉓���h��Zw3�|J�@�D�)0ӏ��<���O����>��)�g̮<J�����L�tnFe����W�.�F��.��}M�M�K��Ԟ"sO�jAn��y�R�i�G�4�e(��a\+���(I2X ��NIF���&?M�PC��vC��9� ���G��g�2)�,l6j0y61�1�K�k{12eqb��$R9�u�Z��C��g\tLz ����N�:s�ϙ��I���,4���3�iW&��z��P�|detV<T�C<0.�#����K�L~�р�ʻ�͍����t�&�pB��'�;Z�Q���v#��o�{kh3�I�%X�+�Ķ�$����V����y���Ռ`��8�M���#^��L=��[n�c(��{��W���ܺ2�j3/&x��sӆl\�l��:@��"$����Qs&~�,.�mD%޺.g'�G�������B'���d������b +������O�(�b�ó������Iu�2�4S�.�J<i��Ur:��N�2d����\��ui��c,���+�C2�Cic����\G���;I���ØS/�#�J��Ty��L3��� ݪEQ��ע�}�[TV˂���(�� �;�_���w6�"I��4Q�uz7�x���h�`>ev��M�1�u�,T��w�S�v�0�vj2STZ+��V9gHҴ���ȕ��G�$�,��Ҍ�
]�0Pj;����h�(�S��53�ҥ�Ng>3r�F�m^_�KJ4f]�\+��O'�H����h]���R������ԭ�(�H��=n��L�2׍nB=��ʐ�P���O���'&��D =�CTZ��8�����X�pnr�3�߃���_@�
IT}��?�wn'��-�>�շN���y���ez|�[ <�˒S���,dOan҈!�i�d�V�Ѡ(QT/�M�8CQN�^O)9=o�:�{Z���ߏ��1J���P��L4\DEH��<�� ���<��!=�X=:��M�[u�j�QV
���F|ꇋzح�;q�a�uu���R:�?	�[3Ki�JM�^�*	j'N�A1{>�:0����F?����[��: H)���d3�<M{�2��M:ɔ;_ɐ&�|� u��{�Gү��D�O� ������1�C�2�%Z�����H,�Z���ݧ��P����d������m� G��_!��f�N�VUl|��-�Ll�o=��5����%��i�'��	�����n/�w�EI��A��>�i�a�!+�נQ�1a⧴�Y��##q� �6���1C3��I~��V��ĕ���[��(�ɍ����r<���_0W�ҿ&5Σ����|2b��"��t$��ڎ�(\f��Z̉�����x�\}IG�j�s��r��ӯc�v?_r���ĕ�	2ZY�a�W������VV#�����ױ��p��ϥ�wn#��B���M�0�X��������H/��Lc�[�P���铺3��iO�p82��v��N"���]���Fo�x��:�ٷ���O�.����{��h��ƍ��r{���w��$�U�v>uO�Fq�A�ɸ�x��ѓ�@�yVs;B����r;/��!�.�-<%�$|��CfË�n�3&�+b� 6�o��f\���|`��u�趽)��E$�(����Y���nO�q|@u���}����	����rr�N꺫��*�zZ�A�p��@N�dG��,p}vi�Ô�?A"*R� ���H���B�C�9 T�.�l����v:�5�=���l�8r��+��Q��h��J��S�$��$�Q�4��%޲^�x~��W���:(�o�[V��H��˾X�w�b`8�T��-���MnY����غT)[f�{��-*���T�B�B��&��Wo�K�!���I�=yޛ��,�=�&  �?J50����fb��0�M�
���}�����N���.m�ͣ=���2�#;�A�$/*G;�i����ł��5�^�J�<�=2��*�)w@�i��Rܠ�����Wqb�#�OKn�x>��}�˒%�lӀ6���&oB ����!����uL=�
M��������A{ݢi9����o�6�k)X�d��Չ�>�V���&��)���=�DͽG3_�OJ����/��K���� ���xA�5��s�J��x�A2���=�&I�~�6��PE�ƈ�|�	mS"c��ܡ!�|, �y5B���ۮ�;������ib�u�s������1�̋�ZB\��)�e�^ڦp^�'?��
H����|��O�U��1�&���U"�Lz	�����I����w����qŒ�g�r�)�CB0��T�8��Kp��h�BK�f���J����m�7d���g닸�n�K�- a4q=�*�
���� �-	���������J�9����V~�A���P�]
�IeS�ɱ�m�������>ǡf;K%�c��5/q;[�'�<�:n �Pc6���F���I�����uT>p]*l��ʢ�[�3;��I9x�PTBZS'_ýy��`3� ����ĸh�E���j`�e������3�U7i
��a����G�v	|�#¯�/�a��Z�U:kN���^��������O|O��[1�l�iGo����y������u~A��{��п���i���󜮩Rͥ�>��uAv�N��m�$�E���Ua�ϐ�l��)?�Ux�@ǁ�U�L����^����0������H��U�r�33�6�ZpÍx8٪K�N�_�64��	q��ɓ�K�W�p������n���d�Q���j�ef3v|�ܲm� zf_��K������������]�:��h]Wޓ��Y5iT���Q�l�g�,1���8�����H���`Y\��B�γCƦd��FG�h/���讑:���E�ʧr����EG�qA;/Ff����L5�+h�O�8K9%���������ש5����Η�3L@�D�w��i��z�����=.�0�C d)��E�o�ֿSh_)�-��������×?t�c�Hd������~;�-0�p�-^V�q�S�9Ce<6�o�,a�i&(;��EܗZ�c�p��S���� �w �jK�{|g��:nJx�="9�~*�7%:��̯�J��LN�9�@3Ƣ�pd?�.�B�:�BN�S3��=���uWsK���,�S�]��'F�;Ŭ#���B��ڻX�@{e'n~C�B3a����xpq�\M����ˠ`��a��7�@�����4���AY��]��%R�q�F�kv+�ä���s����\5��~gȯ��7`UY�������%fJ�!z�L�5�G�s��/ȃ���j4	 �B�.�Zc �xy�ZL�YxX�ш�`1�c<�r�m�8���1m�(�<j�/��x�|��KLu�5ֆ�<7��.L��ު��!&��s}���i��&�!���ʺ8-h�K�Q��ū���I�/��D�f��=R��a�kfb'vu�����e�D��>Z�����y�7��04<>~�9�m'�g���ڕ��w��>�sy�A!ٵK,w���MB����<���_��٤F7V�	�jl��}�q��|�+���l�(�Ʃ���=^Z��DI7&��<���Ȇ'�����%���$���K�h�͉�V��1���bY{��;�-81��
oQbE�Ld��z� 1VN�^BW��1�l{m�n�?�P��܅���c��F潲��$��Y��[汴lqp-���'>��FN!��* m.�a�)ֿw'���lN�.^\Х&�x�)Ѥ��p7��'i�khC���J୩���-�����Y�Z� \;����؀��\4��P�h5���1qL?�����,60����4��Ù��������}qZA��k�qt@ϒ�h�K@!>�:����l�5���(}uy��C-�L>"f��ŊS}��;P��+p~X܎���M��J�}a�e����m�2�e�6�8�Hd��ʭ�[�.j(�WJ����V�H�YѾBGuem�r7J����,v=k�:��I���@UYn����ZZZ��."?�Afg--Tq�o�Re"���N)[��D�lc)�ůMǜCZ��_{���l�CX�@O�"�U�M�s0�� V-�n����$~&^Vz*.�����A|B�L��,#+��.�!*qg��!H|��#LEa�e����լ�Ƒ��������5�}ě+�nd�:�,�#ZI�}��� 3I#J��x�Pr-e�~
��l�?�b���.s�p�z���HL�Z�N�~�����yZv+��%��ei� 	W�c%�@�R�� ~�]���eaS�;LH��HRI�ԴߨZ��=ٔ���L�d 2-@Ň[t�>V�⫃��_�64��!x������Ts��(�&U^�����a5�s��46�'jV�`>�ݽ�ū�N:�_�]����Bk:�Cc��^������Dv�QB�޾o���h�{eg���.b�����(�P"JF��ֹ�0;�-�i/z����]������2�W�Y��'c4"^�y/m~�I��
�A�N�d���B'�oW���D��2
z}��'��-"�q�<Aۍ�Hk/����#uS���ӳ��lOA�����q�M�i���ԅ�ܹ��
~�r�ˮYڄ��E�����_H�ߠ �g��9����ٌۈ�;M`v�̙��B#x�m.z{�k��ʨġT�,'Ȣ!9�ҳ� ~o�:q;�څ��k?e�M�<:�����IR��i[�?.h��g./g�|h����Oc	O��)̅TH�����}Jp��֠�J#@cG��N���خ@���!���3�T�{ƶѢ�e��*��A0�tf�W��;��iwޮ�i9?e������!:����c��V������A}��w?1+�/����,z׋��dq��h�~��NX4��?����n��پ��saqn��m����(@I��_ҥ��-ݙS��a�w(u���C(h 90�"�K�ѣ3��{ZI \�tal}A
7�]�JZǪ��s�ҡC���߃��|,�V�\��s��7��S����Ն�C�v�了���D"[�L񊛩v��P�P3�8TkE�Zߣ��^^E: ��<ȯG$p����:c}$P�[���UeKk!�U)HI�Ӆq.���"-�9�$`�\���8��z�o��m�͢�F��gj��n�4%iJ���ʲ�d�f΃�`ֻ��B?���L�rJ������"h�+��#��3;�?��Ef]�jY�b�o�d$��[��)���l1�w +%RL��Qϋ9Ďt�����_������z�(}��R����M��_�f⦠61���l�}�e�V@�YͪY���v^]��|�U��^�a�*������{�u�s
�&2�_��uڛ��@]�@Jڨ����t��5�y�A`8#�Ӱ^�n�f9YA��G�CUs�����!z����z���x�e���(���>�R�ɔ� ��ӛW�B�I˪=�����ؑ�(�:�h�ᜦ��������]b���z]0�h
�����T�.�����!��.(7L��~J�=Ziq�ơ�n8��YQ�~MM�y��}gIlJ��6���w�U�,cU��IO���+�����P
�+�~'|�e���Qr=���QVc���1��]��z�R�e�5z��(���ғ�d����dO�>��yk�i+�J��^O4��]pǣ��^�̀�%�#!cS/��C�_Sxn�N��N�#�+�>�u0T���%�Ѧ�+"�Q�']@K�qk�9��j��ޓ8�0Ft(٪z�<V;O�-gܮ��?����eކ��`�� �U����-����s�� ��X��?�ҳ~�/n��k�I�w�]i 0��Q�uλt^�f�EÔ?��{�Cv�"��y��t]ضf�4]4��,�a�$��*�z3�JU���ߞ��n|0���*)v�F(�BN���Ê�{ϓ��-���^���~s/�?���"�G���M�����_�DT�(!
hL�4���GS���O���k2Q�d/z�4��7x�eR�J�ƈ�����G	��[Cc+jÎ�&hW�)��"·I��da���J��8�3ǋ��"H�q���A��%SsUتb�R����te7��������sGd�R�P��\��j'0szPp~�<˟E\�'\w�!d�D�yF�������7�G�є��1�*����Ր&W>�m���!�0�|��ݫ>z��?��135V�p+1�[UG}��d��^f5e����?`�P��]^�[���(6~�}M��[b����Wsi��tL�Rͮ�(�)���� ��2��y��t���h=�|��$���<���Oq���l����P��YB-��`�;�T|�EW}��4V�7���d��b��,��	�2�B����ؖLңu�N����)l�WN�&U�H�U�^���ǻ�&��j7�R��zo�,�l���䄁��X�8|���hDķ¾��'c��=�و�x7�ݬ��]��>��JU���G��5�C��fc���e[���ܘ*���K{�d�>]W$��L�Q��H���KKZB3��&֊���
9afɹلVfJ�Ken
��&	U�"��F� ë�;���؃M�O��gn?c�[�:��B��b H�L��	\4�.���֥C�;Yˊ�(W4��d�m��H��{�-v-��]�bct�OO+�k����7`=�5�[V�]5�V�4�)��}�L1��O����o����o=��pY�I(1��B���W����J]Qz���h�W�h��|t(po?W���ӵM��Eb����2c��ѷ�X��ق	c�g�x��RX��%�������isQυ�;��2xI�("`�l�R�>K��'Iq)�鵻A��#}h�J��Sw[��=�)}ETժ����"܎�2�ee@�l�뿙��6]Z��I��Y�RE��8�h�'�8�����_¹"6���r{})�����5�!|��ɯ��w�ɰo��0r��dx���21�B�A�wn[�uc�[�<ʝT���mJ}W�Ovd���N����q6�	����m`\�5�����3����S'[B��
��.����'���퓬Z��)�z���(ӄ����l��p��A`��Js�0Z��������l���Q��=�E��dVN\|��_h����6u���� ow�sw>@-rr/u�M�����%�]�_xuR���0XU3����;�*17�N]k�R���mC���'�)�D ��jk5�$sׄ�� gK�0~ּ����HL=n����k	?.8{a���u�u6h���6��A��~.�\"�v��S	ht7j7���ECZ��"���o������'Y�y�ʅ'��.~ \ U5 1${�i薦���tدEy�<����^C!��b�)j(����"���ŗ�d�l��{ ��/��!����@H�\IS�Js��Q��3x�3��GG�+.�j�y{�Ȇ��?&��v�R�"N�f���⻄�q���Da�P(�D��Ŵ�����` �@�aX>B�a}-��� p� ��a�Z䲄�� ��O���+�5����Æ�m�K���n���>��9���a��I9���f�3>��"vZ�$-fgk���l{뗀#ɯ��SSvc���)�xð�Ҥ���KYM)3^J8ok�s6@��33f:o��T��Q6��x��x܌�����4��� v�0G�����֌��>}ч�#�p�\b��s�
�+]E�3
�B���4�3/Am)΂Ge���m�U^�>-�
:�_�&j��jC8����m.2��њ6|v�f���!�NG��Ҹ�
���?Hms1��!d���i����(8dU��$��k���MOb���K��'1��Qy2vKY)�fS#��2?����0����͇��5���Xqp��]DO�u�t�[��i�MFe�tP��9�A����Y��s>�`D�x���2Wꟽ1��w|�+Ֆ����n���o4�=��7�C��Eo�#�b�����#����%�)�";����Pa���c�$�!�&�!Æ#��ϑ�����DF�����l�u�5�����3��9%�н��b�#InTA�]�T@�(5|\޺������dn\˸�%c�]&uܟO����Q
+�&8�5�	��k��*q�=�k�^p�-pVG�խ�]�;��B%�J��۹<���i�&&|>�2k��n�n쾯8�w!�+�~�ԑA4�z��WrZ�N��OI�b[��p��k�H0�Ձ�{�̡?$}�"^����i��&99��uQ5�`�KE+���O��Ԙ���磐��,wݟq��A/jS�~$CI�M��AGD͏DC!�ˈ���i���t?$�N��3%��n�7��'�$}�&�OBݬ)*&����5F�]�M/Y 1���`�I��Bd���P�YOB8F��G�F��L���%���x�?N�B-�� o.\��-� ��.�z�< �OUG�j���)���R}KAC�$n�Y��M��~:���4N���P���W�^t@aԄ�vk�.i~+K�G���2�q���hX����کi�#����/%|�~ʾN���bb�.]�V��{�������m�sQU!��uge��6o��_�ףi�~��2I���H#�ȋ��>�3Oom�51=~_ﱼ�f�.�b諰$����Tc�Q����%���s��E��JO����bsq�q#���B=,"��uw
}����r���}4S\6�4��ٛ�Ѯ���Ğ�\�O�����4_�}]#a�D�}����|إ��r�ֵsdz��,���>6"�*�aEZ`'"��O����I��?e�k+�_S5cEJ\�uz������!x9�FV�B��D%����;�*W`���jy��/9�Y�8��v�1^�ɱ&4{���<�C{N��EQ0��S��������D��ĳ~9�E��#��5����0\$���b1x�n�i;9�B�c�E�	�
���t�~C�R\)�eԧ�ۗ�6|��׭�k>������
�&A�nnu�C7�{dIX�COc��)?�8�����N�3F������{����	7� $'������"��:�@�8���+]�g���V=��g0����H�`-���%����	� g7�zwm�٬��06��򛟟�T�n*���V�un�9�d�n�Y0�ۋ��R.;�΋���!�N�d�����?(oi�|�%��8w)���G��� w�-��"�o��f<����������yM��2����l����xP�ZӇ���%~O������t�tp��B�蒄�Ε=f����JS�0
��=��	3�d�C�O_6>}�:*��@�JR�!��KCE���[��Cl K����v����'�q^`�o�g��3.i����$EU�sȶ���I��v�]�5R���\�@�c|�4&�'b��]��/4f2.m�jn�M�ٺ�貜#�-�>�^GE��k�j���e7u��U�������z]y�W�v�L��$Op�Yd]!y����i� �� *ð5󶾲����r���s���	a5�Y� ��w���d3�p,�����/Y���۞��T,k1n�6�Jk��V¯�e$*�&޳���Z�Pz@�ۙ�`���H���'U}�Z����z�|�(�(3u�:�<"�b3�w�5@�<ٔ
�f�U6�AGܤ�r80!+7J�F�v=���	^��E��1�%��E���-w ��ٖ�i�'&������%/��������Y,/��s}��O(������J���0�\��������V�X��ݍ����5r/ �h7V��M6e~	���W��P;������}��p���������1�x����o�gA_a��a���c��Tz�<٪�Y�.�d��6��+�M�Q��wC��x}:�����N9XMc���B��E�������
x?�yX�w���Ӡ��!߷1��	�����8L�ލ�b�g��Rcu��I�Q�B�wDK�9	x��J�H%m)�L%�/*9��Z�y��v�1�\�݂��X]�x��ͨ�k^<@�5��BʻrWV3�\��2g-�>���n�@HKT=J��Ujn��3�8-��H��5C�9e�*K��dG
�� _Z D)�mV�TƊm��@��'���6��u=��d��WD��r�~��hU����mp��OcX#1��s"O�ҡ��O� 2�>o��m���޻�A��ӈ�|����ˢ�u=,���D��LS0ϐ����1ib�
b�s?�uO>tm���8�5,�<�](��Ep��~-���.ǀqk����2��<ٽyU��;���o@Cp
ɡ'�}{Ӫ��P#��c�J��%�d*W��?��m�z=���n��� �+�E�i��`�n:�3�u}�Z<�s|O�8���k��+�0$�R�64���&�cs`	������W~�W���Fcΰo!q}W$\���)?n>-g�!���フ�nX�]�
�*j�.]kn�Ac|��Kg�hڋ�^�\,��d����Xa��_rT��Q�1f�7�&�>J��>ڣ/%��m��F`E�?��Oƫ�����O�N�@���}��C�qG������IJ����8Ϛŉ˕�<1AP���v�6�vh�(��O|�b��h[Y/�$�]�ڶ��pW�h���tR3���Zr�=�˃������sYW6J$�X����A�"��K��O��w]>l�j��V�h������zE{=}Ȣ��z7g��Z�L������aYߙ��c���
?~�JЅI�"��*E�n���4�ĕ���������k��'�_�Nw*��D9�BBf�y��*���y%|�M72�^�$�1g��J��5Qᇵ�?m2dgk��ܗ��g�5@���z��ü��;������W ��g�xG��/�V���@����m�uue�*��<4�c�͜�O�|EL#��#wy���b��e�e�Ǳ�©�k��O�rsЛ���&3�>!	�=�N�+0b���cj���9���''/.�hV���i��B�&����~�K�r���G� 	ktF!��ͣ��}��LA�"�nvz��\�W1�Iˑ��ޒ�����c]�E!�n��y��q������񽅎����7��U����-��`���M~��aw���f-����Êm���j5���J-��X�o��
6�`�NP.�J���Lbx_�W����c錄Ua;�3u��o1��w��òi�/i�徱qm�tޱ�To���ks�ٺ�Y9iɈ��������q��#����y��!�֗�plʄ�E�n+x�H�ψ���@���k�@� ,Ѧ�x�*�{�:�j�W�/�W=��Ó2��(n���r�0����*�y6���П�z�F1�^��!kv���"�ba�Am#Z{��Ch�Y�j �ߡE���V�V K�#����
CgRC��-}eSʒ�K5��e[���V��M髽]����!��4�`z�0�!2+Χ_;z)v�����z	��t/b��\Y/=������_�}Ii�֪V��xot�R������k��Vd�:0�ݸe���X��6�}T#{�p�ӥttn�,�mµ5E�A�����s��V�ws�F��@�	Q�O}!�y���"
q�����-����*�ڳ��)z̓d�2����"���r�[��P�{�����f(�4��f`�
�8���`���Vd��G2W�Ԕ0�9�'�{�G�DDj�@��g�u�N�KJ������H�����*r�v]ϻ� �����1W����F��%M�׊u���g����=���U����"�i3�tO��:V������192��#q<�L�N�n���$7�+�f)��gL�������SY�6��c�C�Hqql>h����c4`5�� ݙZ ���ߛ��sO��s��g�
��2���d`�⺲�4B��v�,@B�����#��������n�ǻ�t`..Lծ�t�/u�;�W��i�%����Fvj���a\5��	!Jh��ihR��u�vx:�f��3����=�wE$Ȓdo�C����w_�Y� �驒r��RdWM�����{;|�_�{��ύ'��.���g��Ḥ&��ĭJ�ρ����3'�N��~�}�yuʇ�{���ߦ��1��G?��gʦ�^ ,!s����f�R$tIsiُ�&e��`.0��,�k<v;�Z���.����C+��僅]���Z�Ŭ��}-�����Œ)<w��ɫ����)w��bԷ��Kp_��EmӇOY�,�g�Q���b:)�W��Rq�.\�4V�FZ'����K�	hn�R���c:ē�8׽���Ӛ�3 �s<�[K��	���&����헷����9�Fz���a���,�=i�)��9	n��MKU�=c�g2z<`<`��`�T��4��ظ}ܫ쮴�2#S�=�yXّ��?6{�6����Q�_ڳU�-Ϧ[�M��h�×r����@Z	�hz���%F֬e*S�/���/D����fhqnΩ��_�A�-��0�L���
�!G*﷞�߆�ɞ���I)/d�柰@Q�i�5S�dzp�9�4L�ژדK�h"'��a�\�8V�T�Γ�
z`����_,�F������pB=�6��d3���c��<Ym$_���e���7P��3�wi'�W�,W/�#6����D�@«��&}Z�K�bv##;GOtau�3yrSu�5���f�J�����x�/�`���L��x�R>��k���9���8pT2�'Pg���?9`�������8x#��b	�OD������\�7���d!:�@e�ڏB	ʇP�}�'ԉ����O���7��&򎜾KY.���z�GM�N���hܻ@�V¶���_��[��y�k��-�9[S`?�3C�z�`#ܺ����٫�T���o�vS_W[GΌ/��~w�>(����.�1Fy��g�����3W%��ҋ�l���rW���:�a�BU���� ߙ� �*iJ4�����N/5��i�!ɺPi�cN�nh�1S�,�l�ES
�G���-ni��7>�8t����~�Z��5���i�r�����48)CFRA�	��*H=���֨h\�X�����N�F^^����<�	/^ՙ�_���K7�+��Z]4�!;l�n�:�?������ֿ�d�q��V7���"��tY��y*�$<)���g���E��4|��Ftls�����w&[���a+�c ���Iأ8��O+���3�_������,���^b������t����ѳ:0�l��'��fL�C��՘px�4W�[�+��q��m��y�ԩa{���cg3��^v���Յ����,�\�D��� v��C^��sv=\�*m���7��7bW���^7����q�ċ�"��P�M�/���f.���]l�6M�+f/�i���c�v�ՠ�q����b��]R�}p'�aL~VKV��][�:l*�Ĝ"��B�a�]Z�\Z��M����i��^��vG&�\�άp_�����|Ȑѿe]�L�֑R�&��̑VA�'C���	���v�`K@OuδI�N�o�^��X������u�3�姳���gq�?��h.g�f9iz�gy�9�{�<�Y6�i�	����w�W�hzu0P�i���s������9{��ma��t׵ڵv���i�A�ӻ)�G��}���L�}�)�(�1㆞��w���G���>*iS���7,�;�Mũ�п���y[g��U���-����w�:��]/�G����2���Z�Y1~�?��?��m2�o�YN@�y[;�GRT�w��~��PK   �cW���/�� Z� /   images/d3087b83-655e-4811-b17d-9d66f7a3b2a5.png��US� ��%�[pw� �5�;��ap� �	n��;���������}����˩���>�j*��(�(   ]^N�  �  �#!�'bh� �T�JI��KIQ��9[�:X �9i�jz�K�ct�B9�nyg`q�,�"	2�Rp����+p9$�)�-��_b)���k=�zCéy��0U�����M>���ô�Æ���;9 �I�Z>�`�^��\i�s`���1 ��Y�"��ҥ�[��#w�U׺�o�11�S� )����G.�+�9R�Z'v��.�@+�R52���x��t4N�X�i�1`{\$����S���4.G��?�b,Wg6������"�c����Y5�G���Ǝ�g�8��1�����̖�?G��kk*�K+��T~M�N�U�7�'�5.�<��>0^d�tx�V�J#��C��}�2��s��I�a}�o~1>sǞV��(~1IUQ������	j���c�����4�|}�t��v��t�X��`�p���r��{A=�%9���A�������k�
;����մ�����gH����*3�9fL�1@D�K9 N�s`)c?�9,�Q�	��l�cU.��!�/�<t	
_��va8�x"qBTֹ�h�3�䮛X]) S�������T�h��oO\�Ŏ��9�H?�d�a�L�&�xu��}dް�Xp�_>G��)��h�o�Mu�c$W�ZB���C`�9P��]�a���]D��f1�C̮��$��B����n)-�>5D�&��#�K쨑� �J��!�F.I��i"�������,�oF�~9B�%����8�C�Yu� Ef��`��-⹠�#9��.ow֑"' b��nյ�cBQ���}[P�D�$�
��h�%�֪u�C[Z��;s��Y�AQ�,��ٴ#�#:�g�Ѹ��B�&�tB~4�X��\�ߜ͙8�������~,�}Y�Fu�+L "���c=�|0a�E@9�v� fo���k�y�T[c�A[���rmd����޵�?��4+!ULA��<�/��EBWaEbE�;��-�L4���/DΔLC�jJ>,�O�[)r�aS�m���k%%$�����UZ�rE�����_���l����1��:+��F6�}�m��|*��h��eB��ͨ��˸�ͷDI�Oۚ�]sZ�MG��_�'J� KMP�ܓ�9�7�7Q藤F��ָ�^���ߘ��Z9�ѕ���j��'��b�1�r{��M�MM�M�B�N
�s�%���*�uY�YE�Mk�������b����He�6�fN�N<}�}C�Y�0��y�xÈi�㉽x��x�x�y�m��Ŗ$���O-�W7+��Z�E{F{ z%��N��.@�7�i�>�
0�ա����ht2��&�l���{A��E4+�,O�9��M��K��s�ڴ�;�������V�N]	�
1:9�'t���u����8kV�J~_S%k�2Bg��wSs�OKū����<3M��d���	��ꑳ���<���Rx��dsu+��O--�zMgY�?��4D�D��֙�+���Yfd�F��o�G��֩ʑS����-���!g(g�������K5�W2m�&�.P��Ѕۙ�/�)����������ƶȑ�~�v��_��i�#�p�s�M�����*��y��Ʌ����f�W.mN��v~d0�Eb�F�����u������k��#�+��iv��j�J��C@����ˆ ����z���'7�2P=0-P��5���-6&>u�	�ktq�_���eFޗ�������eT�TsIK�Wg��6�Y"�"e��anR��b��(/�l ��������H/�Yj���q��8�T��~��`�d���0��$��l ��V>�Y�w�w�Ֆ�m�����:&��cpx7�e���|B�
aY��칺�������'dNdD��+Iޮdi�݄!3�����o۬+Ԅ��Ha����V�3��)�����%?�Т~)�9]�[8Y��-�}����#�"B&����q�+u:H�d�.)���q�X��eAO_��ZEm0p;���0��{���}�� ����v�BQ3=*��Į���X"/:31;�8��~�n����7��6�{(ͱ
Mr2�9&^��&�x��o�4Tm˺�8�~�B��L]Bm����¾*H��Ṿq�����ӗ��o�s���OO!�ê��K^N.�:{P���]�2�o���~?��@7���K,':kb[��Xj�2t�t�H�W������Ӽ��+���_2@���Lk���ĕ���U����8ue#ť�� ���˯����v�vUK��i�u�S��'��'b3�Sy��]h�E��ʃ�b��`����1��4h��׃]l�Y��v}MF��^!���Dyp�q�_z[:$�����������sY�JU.�%»�jre������a�4}��������Y����0;�I����\8htu�<C�ȵ��ө��r.$�q�'w:W��Щiã{u���t���������w��)���Q��w1�K�}+қ�q��X�yCaF�&R*������f���������|����K�'�{
�g�|��4�#��֠@�٠��X�g�����	:ֵ	ߖ�vVvޗ�-����;?r�:[���/����O�O�}�Ke	3���2A��v��wW��D��~��A)H�����? ������ge�pY����W���yX6��<XJ.
��3���.��u:�IF�����^��w]P�CjAg� ū�����2�=u�~�^��?����  �����m|���v���q�?~��������������c\8�@���W��Tfz���I��>f���tn�X�7�sO����훠�e���APn�u��[�sT\3�s��e��s��R����o>x����?��?��?���A-��uz�I-8V�����M��U�*��/!�7/��?�B����Bsڇ*kB��S�����Bwo	�gG���6�R������C0L����/����8?��v����2��fjU�s���b���}YU�������_��3��I��`�0����fnE�,C���M�{Y�<#RSM~�����B�|��O�m�������bu����c;���x���>�[N�V���׃G볯���榰ѳOUsZ�>+���i����zn�4��F���fͮ��U��c�[7����S���y����M���RGQH���d�̱,�Ie�������ᶵ����szm������������%�����������c���A����}O���ŏ�KϚƫ��'����Z�U�p��j�P[c{s��1�y37U
>�G0Q^P�^�?�>X�(�>��V�֕h��*��!�&폹����O��ſ�K�k��tT��|����;��Ck��e<�Ҵu�A�SlF���-�����'�d$/�l���=�Z���ׁ�p�/Ϫ��ju���(jۯ/���έ��0(p� ���@��$!;�P"����^G�#w@I:gV?6!��"���_0rBFKK�`�R�e��h��+����O�p���D6$J���*�Yb�.L�vq���@X9��U��)h(bo��&�7�.���h���o��g'I �����W~�	���p������n�^�ˎ����xȅ�o;�GO��8�k��8�u"B�rC��]�o��t�A^�ܓ���e==�sXD̦�˭�G�q�o��Y`�����(��an�JiBi�~�n���-l�J1Z��'��шp�t;�@��m �R-E~Ҋ@������I]1��{2�Ñg���pB�(ٿa�+u����\�G�������_]�z*j�.ʙ�//����id|,~��X�/9�v*.����G��xױ�tC:��Qj��C���v��`Hq�Tc���8 �)�g�����X;��)9��������YzRl4N�֜&���x�t���_'���X1�!�ϟ�5gn�io�,�M�c[&b2�O W�ݬ_4��k��7�';f�s}���a�o�>�b��l�dnAW��WW�||��n7֢W��&Y�7[D�\t,�lf����ڻߺUI�H_��	M����k��͍�M;�R'��x� eV<�S1�V�׺����amE��tc[=o3&�OMIA-�s�$��,�W���?�$B^��o�5�*XH������ ��3��w�C-2
j��r#]��s�0�W�m hX�	F�'�}�]�M��U$0`+�
���l`Ϧ�W؃�	�#r�&k��En����_5�yfr�xx��Y��n����Luq5Zol,-�L� ��m����)m%�KuH��6*[_U^�F�Ñ�c�ֈ����r��E�s��s�R`�緍<w_@��ًd08�5��sp�@�V�� �8@)5����m0&�wJ6��{#��\�o�/}����9�ڝ;��n�{o���U]���(��)�d_[�&�҂��/�o�a	�m�0<�8�#��z�Y&���xW�{�ޒ�k��A����ԑ���d���R�=�����/p!v0Z�`�`�AGH-_"��H\F�pF��3��Q��d��}�ë���E�3�z�����̉�i���O�����A7� qVT��*���h�;���71�a��u����.ͽ9]'X7.Ҩ�,�sԱ!�]b�f���`v՝��Y�;~����xK��;2�@Dݠ��"�ډ'�[�Gdg�9�5#�QwZ:����#	g@���S0c=p��ƥ =�/��0�I�]]�@�/l�5-�~-,������%=aD���>3}*�#&�YYp��������X��GA�š,�1<r��K�n~a_Ȧhk�q}P���a	�^|��,�;����	j4+6z�r�~:��FG����>����}����yI'�Ŭ����}�[�rJ��4�Z���$�%.7*��P�H(T�r9	�Y�-���p����L;�&�-Ҫ0�.�5����ͯ�P���,'�>/�Opx�uHj���r����9��Žgh�-��*G|�������Rr�w�+��ɉ�����)�?���]5�1�F(�(�Tg}�$��/>�7t�'dx�|�_f#��~��ԅp�M1�����d#+E�f(ӬG�;[�@��@+?9��!�j�6��J֪�9_\��4Vl�TM�!ٗ+�[(�� �< �$����� ���@�[�.�њe~��}-�O_�`�&iN�|��x���� �+S�M��<>ᚙ�J9iF�;YY���0�F�J��.�e�Ss�t�L`����D؆z:hp
qZ[�����Yr���)��d2XI�TI�I��8815ƓY 	 �d+� u6l����s��ޞl�������%�~������f�@�~BRD�xw�\g�/�g�u���CӪ��m?Ӑb�1X���R׾�ݍ��YؼD��8�N e�����wtu9�	!  �fzT�֢nܕ�b2�\܃�kNGB�������	qu|�� ���):�����I�yX�a�͹����_�D{x%7�pV�,G�� �O�f���JɁ�o72��(��?��#�{*\��ϏHICZ7a`r��D�%�.���I#&�5}AуGgv�<����އ~������e�a]J�f���n�E{߇*��׉���(�����Bm�m����:AXs( �9Gv�-6g���7���q&�u�E�CqWk��Z=�pz��B�CHO�*wCm�s7��Gpn"X�[�F5���[�-;����pF�e�%gU��g[c"J��������Z�;���]�YN`Xr��	�l�^h�p�pt�ԧ�o����	�js{��πY��).�u�zv�o��P�I�~��=m�o���4X�:�o�T�[��W�B��Z��LΚ�ha0PS�Rp�I��7bv
��5�ʿ�@p�� ��r"��C�1�$44�)�涷Մ�ov~�?񈊞����`��/��U.��Ȅ�--Y񻄍��I2+�{rGF�K�W�G|�8���E[%��s�%T�6�(r�賟9�,_F޸X��<ja\�Ҁ��h�T *��@	�em�q8ԁb
�/�$����2�ef�O�O�>���"|�~�(�M[��緐��f��3�M���d!3��_���ȾfԌL����2�ly7'���u��� ������*�����68k�Q��]/�)�1pW[�i�/��ʻ�?2:.]wV�:�Y��H N�b;��Fh�t�м��5F?ZC
�_j>��� �6|��	��s���̄�i�j*V��q�H�:ʝF�nY����<�����+?[�|Ej����~�7�9��ax&"��<���k&4��v�x�����dO115#"2bn�w��u �t����{��8��l���:�yU �z?p�#aa���(K R:�VtLA쮤8�p�4�q`�ܺDm����`������J*=�xx�=��>��t66���B�94��N����w�S&|�9Y�]%��;�˯%�})vd�#�v��^�#��"��G�߳7ۣ��u����>����v,�����'�4��8���o�~�Px�G;�F5�[�K����z���4�K��b�Qc�:v�`58��x�rU~G��g�҂qdw�Nm�A����qX"4��`�W�m��� 8 (+{�T�%���&24�L,�J�J*\l_.���c��k�ڇW�J���'v��n����9��wN'�.08�H������{� �c�j���JQ�����V�Δv%�	m��,�=v��u-�py͟��R��/f�1���-K��W�@�Q1���㯜���4e
�gE�3�f-u�:���d�vڡM�����Ґ)�#&,#`Xu(he�@�qV��9��*�f�������!�%��}�<�gr6�E���6WA$�0ʁ��d��j��Jʮwk�a����0a�1L~�\�����`��Q� ĲA�n���G�����<Bp5��H�H
	 �r��U�v�z��8X�h^�,�m9��U=Q�0�ae��!d.��-[����	P+m(��ƶh`J��i\��m�x��ro��f6+�����ٺ�?~���|� Ks$����l���t��HP���3ݝy��^o�x�v��ǧ5��Bo<��oJҗ����< N��V�{�-V�M�6����1�5}?��$��rҖ�-���<�S��ݦ�~x��j�#�;��p�i��z��|p����V����
?,���Ԍ�N8a���uQGXD�NB�[h�x��ҞMV(������iSC1ҹ�?9dG�b��Z^��Q�?=�#�p�3��ȓ)��r8zn���1:��������K��\�^�<����U��y  ����A��{-�h�D��/��̐ڱ�N�o����CpT�H��܎Ћ��>�/E^]ܭj����.��S�x}l����i.nfj��Z_��U�'e�~;�����T�#M���А� `��"�#����b�UI�%Õr��+D��V
�[�o�� %�}�F���ź�KIӘE�FHl8��g�Q�W���I6
�mtyNӃ=�������5j��7tt-0��d����)����L�p����Z+�B�.5h���oPz�Q�Ų!�FyJ��ɦp�긣��ET*����
u�z8�	��m�3��:V-Bq��'|��4���}��R��-��nA�|[�Sd+cZ�YR��T�rT��b[]��Z�BXo�2��>�#5�)��pV�;Qs�S��t�ZEia!�Um|��I���{�g[�b���Z��t9{cZ���"�a���Cс�	 ����L(*:֝˹�����^B)}�+�G,�������V��߁�5�s�h�٤���'��"Ŝ=p�FA\V��Xw�/��[е�m�S�.�r�����pARq^rG^$[p���
�c����EG�O'G~�����;���r���T]�M��K9�hǻ�-��z��k�Fhq�˨*����~�KJ���7�_����$�-�	�K��	�F� ���&�4���Q�҉�{��쎟B�� ��Y׊��R
�o�����3�缝�e�ٲa�c��r\�u>y��~�#��㛻b��X=�B�-hol�5�u$�1vh�۝�������o��vT�Δfj��*y��@{T5M�O�O�鯰�r7w�JN��1���Ek�E��쯽��+�[{��)��$��+����h������0�f��I{���:�^<�J��L�~�Z���G�����(:�(׻���9�6�a��T��+��]���hϠ,�{� �<�p9$�Dˡ!�pzE�b�S�����z�&^�8�����o��N���߿�"�m�g!pCH��C�"�����&ЕylF@���2"�	���վ�y��<�	Ġ�&�?�;�Tm��t��c�;-UES��K�&��8� �@�;��#�N'���}�"R��CKV���h�"�6�����a�N%d�\x~�6�#��^n�tpR�z`:�a�C���n��X����f��N+��д��0��̀�� t4�b��eW�(�h=h�+�iX�`$"<n��[r� ~��[�^��Z�I�+�1:�kV���B�0��e��·�n^m~&r�G���
֥Ner\�s�W��Dl�p�|�!�fp߬Iq�z���Iw��a�2�!д3=���� a=Q93�Z4'sA=�e��0܊i~���Ȥ����np[>�rK�����a�J��M�|R*�E`� ~�ia��Jg�h�.� {Op� HٗA��a�C6Y%�`z`Q>��8��MM/����t���˞1�͎�l��u��گD���AI����z:h�J@؝�]�z�*^8:%ā�*$�`QN�k�_v�Cgr�ï����٤��{�6w� W%�ڬ��?fΟ:x�g��mW?�r�qf�i���i����%:}���ѝ��(0Q:�_�6:���y�%���������(��|;oo˪�V
�����ϒ�T��M+ϷԛS̥CtCP���}sޚ������I*��nu8>轧�}���#�?pX� \@B:G��w�:Y4�[��d^o�U��Y?�7�����u���I���y��ݽW�}����e�)R\�ꌹ,�\��"|q��S"?4������ڡ_㪂E�	Ot%N�[�� ��$-�V���B��=���ia�<sDv���Q�G���� `^Q:�Z��Pa+8�0`S��R����
��UH%&cИ�f)�ɴj�j�u��̿�f��E$��끲��\s�X���x-A#ղ6�7���F8]S�DWHt�;�� �ս-nk�)�Ԝ~^��%b�/|�!�Rt��D|1AF�z�~����PE[kk>O���`���Ւ؊��(#��u�l��ӓ��z��;*��6�(��Q� \�nX�u=��E���PZ��U����$m8�:���-x~�<����w� �ASض��x,&����ـ`�>`�fp%/��\蘊Ԟ�V����F�|�@u�4�d58�Ô�g٨mc�o��e,G��L�u>��<��V�P����t�I��8"�U�wj=�k��&�i����\����O�s.=>�����G1�K��2�Dq\ė�2$bv���I��`5��*�'���:�:��L>�� @�L.�=�"��y�4["��O!s�|��'X�� �A3������p�m����Ī��U���/�?w���W�����r!��\�뼐�H<��@u���\�qa�iD̶ڡc&,my���A��}
]�kA"y�̴Y%Y� ��5'�`�
x.9���s4yK�P�����L���N_��J���w�n��K����:Q����?�jP���Ѧ窭�X�Mnk~^����?��������]#cgYT\,�Т����ѱ��y���+�w��Sy=W���^d/�����ۏ�'E�3�g�O3�S�|	�3Ϻ��,�5:V%x�2xS@��!p	9ص���1H �M�J���Pe̔�V�e�'�9��9�,,��AJ�v���&#3��Qjy�E_�Չ�2>���`�F�����} y\�X��f���g�)VH���B�;|�mVm����͝�&��SlRc02�ez���-�J�9Vv�x�P/���6�R7�=H��쌊�gS|ggZ)���׺oe���g���!i ep�<'�o��[ ��`�j8��X"j0�2�!5�,[l��DB��^�r����%X�6o̒����л�A�-�y������Y�|zK�_o.�p�Ư2��d넧;��W#����*�H�$��je�e߲m�\���ص7�nߠ�w���
`��tS�w����Eτ������5�b��
~�w��5�i���Űb2P�w4�e�F �O.��LX#���� ����������6<�L�
�ow,A��B�#4��4�� cш+*3b|��O�h�i����	����c���o'�L �׸�݁.!��
�ώ�'ľ��k+����	�R�)�HP�JD�=?����������K�O���T�f�w�0�[��}녎rK�m���ūJ�%��l����:.�Ɏ~�}<�S���z�r޴�v���@W'ix��v�.���{޵_nA_RӾ�W���Ɩ��&O�����{a轿��Ä8���3i<���]��me�>�pP�Kq">�y%���_����wy�L�8�{�:޹��yu�ۧb�#4�x)����� P�Q)��Y��w�7��]���[�H��+���z���);�Ԯ�̚�#����J�%Sԇ��W�[�x<$&�j�a��#䁑���h�v"1�sQ[d÷�PC�^�P�n�BX��X�!��:��h;K��'ѷ֠��=�=�7\���}��wƤ�{��ʞ�G}s�����б�g3tF�_�V¦CE�!�-��`.����|Ū��P��\����ʱ���ĺa�#e�Jɗ}2a�L0�[p��C�Fr3���}UNLb���Φ��IgGg=�>9m�1���IРϮա�XK�D}�^"�=L5h`���� biWOhG��U��զ$�נl���_�6���A>�Yu/u�ꠓ��l��t������#�j���0VE����u&0��37�#�����Y cC]�-����t�9�I����}���W2�6�KB\�I��}:��R䇛S�#6RO�m�<�4)\E���͔9����ȏ�k���]���k��m�S�A�X�e�=>u/ 5�ah�i^*eAy�b��Yq��Uڿ�|����%@s�lD������;4F [=����E�1Y����J|�M��gEv�N�]����/�x	:�����W�X4���q��n𿍝�����Ӕ��:U�o���t�a�����?���7y�B��L�����I̢��]�q75s��X ���/��_O� �{M�Th��?�n�ݘ�߇�Od�z�_��-���7�b�H�� 0��=����i+x
�d����m$�aیe��hN:�H�h)��+��ʪt���ğ�fIȷo�ˤ�e����5�Պ6x��g�O�	&���V�;QM4�99
̨�Ϋ؈80c�.�U&Zt�wm�������;�bNJ!����f��Դ�� B�d��KD4�>�/١Z�*` X.Wզ�S��Ͼ�Xŉ,��i�a> �|.͹���ְ����Qʯ��,����+��gF��G��9Vb����e]&RY+l�<~CB�+bݮ�'���nǙ��ř�g�{�h��%"�&���\[J����I���.�D�M�gJ�IDৎ�L�"�G&��8B��-��\�P��b@S�.`wӊ�D�&�KHõ!%�ن]�*�c�����'-�lu+bww�E��U�V�!�-�A�EW"��&?{�x����Ռ	j�h�h���+���'$�F�r�QB+#�X���'@w����;�}w�6Afx�$��]8YY�a��QO�����P,vw�l�.�9R�b7'��K���Ӟ{���V�E�4�@� O����4=��3��)|��#O��cNN�-�"�fi9p�}b�>�i�y�g!�%�(|����3���=Z��ƥh��&�ɑ�.+KZߋ���
q��|���D���2�h"�ӣ{�_��F�~�����S0����<(S [a+%�����2��U�z�I���`�X�G�� ���1�:��L�\��^��>J	-@�i�
�U2_��y_٦�˚K� :���&)�J���������I��#:ԯۚ��>4����{F�Wm�?@�A�g��w��@+83E�Ɗ�0�&n�gG���	���6Vf�_��c�;��ho�T�Y���=t�z�ӡ���P�*��Ç1�Y|������)���T��,�-���F��͠�R�E��)+�D��x�*��}�v�|ߞU��\=�)���yÎ�w��k�{G��9N����6?����v�Q���AA���,�:�NB���,�L�]Pؘmg��4���TP�yc`?h�#e2��DS�r?��<�N�F�t���F-�:(��� u�t��jKT�����vw<s��/��߻�"��|���}��� ��҇�@/Q�9�3���z��P*� �ݧ�-�d��P�Z��a�R�])��0�}|��K�����H	��ƿu��<D6#~��*���#��Ū���
z�������R#u������^��LC#�U�S����~�����l��N!��Y�~x��>�Va_baa�?H��s��ǳccV�ЅȣǞ䩠{w���'��>܀#:�6��m��%�QS������[&Q�%��W�"�y�y��a��=T©�ѩ�`�e5X'���$� �>��Fq���0�ҳ�"op��58`��������*��2����Q�N=����t7	���\Ao��Q�
�(қ2�}	�"#oD6�_1,(���0Nv�� }=B[{��x,n�fb@JJxcn�m�ݰ�SG�f]A�g�E*�=����������p҈䵞��� L�+
A��L:�t�)��8e�B�� (��]fg��}�̔�hfzEmFuy��6�Ve�R�_1�,��OSsj�a�@lՇ,�o�5�g��S9kڂ]Y��0��B����X�>>�^��w�I����oJY�*�����6����N_�e��y޺��En�-��r>����n���̖E����U�D�w_��D�P|o� _D�nh_��y|���<5�Ji������!�7t-_O;;�e5(�@_�>���J�|����% � :��.�8M@�\��"������ja,���ڄ�����vT�*��&��o*�_�Mi����w���6�����^�q4`���"t?�b�<�ã u�m:��:�ѓT�T ��`�x����vv4;A_�}vSؿ�6�\\�%7��s��>Wr}1L�i�E�����&�ȍ�X�Е+��;�ƍa�ݧWԏ�*mh�UR��܍+~���%b�9�Ҥ�<���,�����T��,ZcuP���"ľގcO?����]�=�b��^pՆ�뿮���Wt4�Ns	�Q{T��?{e'U�H^��t`2��{��r�����fzT���D��hUm���3`i��jQ�v7����|��U��~_�� �y�������Xգ �;����s4 �k��⥄����������ӈ��ٴ��%z�4�Et��7l�O��p�n]bw�g��;_eMy�Ţ�9R��?l�Y|3i$ϝ1�.��r��q�4m�[�ʅ�����	��>xʁ�2��jo�X	��Ӻ�>)���P*���?53)���}FY�<�@��G��BF�s�p9����:d��1�[%�P[F��X��-��ך���C�uX���Ml�/�m�"BC�9�@��Yɒ aLO����E�R���}�HZ��?t�r��({2�y��\T�������� m_���q���}@����&=���Wk��2\Mަ���㓏'a�� [�=��[���;s��m��Ҵ���*p��s��a/S/<����B\��q:3��aMk���VVou���m½RB%���E�N��Å�>K,�Z%z�P���/���x(�����<k�};/�p���N�&�����*4,
���Ac$+f�5)�YG�Pn[�J2��t�F���A����6'�S��6���.���j�j܈IG�3���ʒ��Enc��Ot�gC~J���~.|���Np��C$�(��nG�0������u9ši
�.��my���u5yO��2������rul�,&���:�1uI�x���H�j�8J�붆6����Z`P��Af_Xr���98]U$�����o�`x:{�a���9C� �n��?T�iD�s�fʓ��!��yd��H7O�[e(������H>Հ�:�=mb��>s%ry��qݣna8$`��"MN~
'�tx��k"$Ǎ�x�n��8�E4�E?;<�s���&�p���E�0���='�η@��lH`��nn���E򪭗To6^����(������*��Kه{M9�Q%q�ȼ@���9��뀣[H��/]Í �{o�(�60F�w�0S������ㅦ�͑�W��i�gI�E�p�n��yA_K� �-��xW=�3��^�J^���R!#�\���R;����0�������"�H�g�B4�{�۳{��䢠q��E��8�E�cML���-s��6����~�2v��OWs<�ߨ������e�0����JH��5Ra���՚:�g��3��m���t)d�f���2'�����8W� {,� HH�`�̬��l��α�!W7n(7U�Z���L1<P�#�V��v�Y��e�e9<�j�^��A���y�B6��t6�E��
�R=#���1��;��o���3�"Iwh!V�}���_��x�C�q�m�Ex�p����#9`�.��"��F�`��?L����X�θ2MY<F/D�o�>���1��1���t1�����>�m����q��%\.����(�f��N�₆���~��ܦ�I" '�a��W�k��	iO4����3Q(@�	{ݼ4�el���c�ܦ� ��^w����[�ȕ�yZ���w�	���HԴ(���Iu�	NI*I�
PZo�R]kub�)W|f@с̉O�MTQ��%�s�ʇ�[ޫY�m3�Ŝ¤\��	����l��<����7�Yy:������j�N��~�ӓ�͵4	���C�8y����$�����;�����A��=�����ōx?���=����-����du�X�B�y����?֪&�=nӺm������f��_��M5�A��]P��~�A��G��%[]��Hi.yq���%�"��ȷТ� �;f��^��c�U+y13�_���5Ƽ��*���Z��V�,��a5�K
N�<��Vӎ5�7^�HWG&���>�%F���� �~J�f�wyP�!� B���R�H����]�taRF\�+w6`ఊh��໨yI��T��ZѬ�� ǘ��\j�.7xD\:srK��	X"x#�Bs?"*�x��.b�6Z�r�Oc�sD%#i�	������'^�t��xQC�B2	��x����%VD�Ab��X{p�L���Ԕ�R6ױa��.dvےChLj`��҅AR^QRi����p)\ό�9U����u	���G�����u�s&�lq�� qf*	(1w�pJ����!�M��T�$�~j�f8���T���Xc�hƢ���f�w{hڐs��1��OR)g
�Z��-�i.�u���$"�yS��Ɛ@�_�H�ŞnS�ƄB�&�c�f���2�r`qʍ��/�����?�v��Eh��C<u����a��Quv�݉KL����Z��a��P�M��!E����>��.K$ծ�F.o0�b59x�]�H�n�mb{H�1���<]�r�0�K��"�v�Mt�w߼���������2 �q^VO2ҍ�RƧ�������7K�|_t�{�#����!Ԃ��c�����.�4W�:� ��� 9��N�Ձr+]*N��yri��
N�:��Qq#
.$�ᝍ�Nή,Yd�E�g�!���=�Pq�K1=�ti�6��熀H���0֥��$��C��"������K�/�RO� S@��(f�  K��Dx�c�z}=\����4��5Y��T#�F3Y�mbb,ͨc������z:	d�jמw��,���Y	��6�P8��ѣ���r�AN��Bw9�H$�GH�z�m���tH����U�A�η���0&�r��o�%M؟��v�"�]sܲ�C�U&3��pcl��h�	W�(�7�K����&�200�p*�Z~e͘Ac�����ᜑ}�C~�%B��x���ԫyu��Y�S�Sa���ܪ���s'P��s!�mU��^�:���J�v�@�چ��i���z�D{~��P�pC ���Ȓ��P?�PZ����q�B���*�m�4���;U�Ǌ����i�V�5M�ѽ����T���,S��ړp�ٹȿ��f��=ը����DZ;or$}��w����w@�e��X �+�P�_�L�Y���+8������xm+���N���i�/�95��1rM�?:$˖�T��d�B�L��r-@k�t-[n���lZ3v�g5�����S�K�յ�N��险����ޡ	5#�fM�*�J�����( ��Yp����rlr&T~����<?2r�}ݏ^�xq�f}s���Ң����*�cv��N��� �.��,C�è@�~��p,d�_���]x#��h�~[T�u�^e�iq�h��߀@���u�B�k�� ����Ј��P9�)�	rV�λ�>���V��'}�W����?:2(���C��|.�x�7���&c�v�õYH����������5�t&�҇m�&7�ň'*�*�eD�,�ދ�.9�wp�^U�]I��K�����NˋjN9�������6�@ ��c��m��i���|+В�]�������8�z�f��(��6�1+�C��y������ߟ���C�����'�H��$�C��q!L��,ʹ�Y�FtU-���F�#�2y�sv��KAtiw�L��_�Y�b��^9����[oQ��D�r��Zt4wk�b h�u�ޭ
{b�e����#|^�du:7�r�P���DZ��n��GߠAH�ѪHa�����r��Ar�Tk�� i� �a5� �����|.�Y��Ω�=���n��~@����N��z\�]_\�ɛ(Z_��:p���۰(åX���sY�9ׇَwC��L��c��%���b����W���hֵ/�յO��~d������1�<׷�s��=�z1N�ғ��v�@�m�-�����},��{���O��º��}Wf��Xo�L ^h_Ϯ��4���s�yW�"�[�L:�	�9V	D�zq���P����1	�\/�����b�R�"'>15�z� ����T��jǟE��.9	�I["H����Vw��hw��pв*4�oϔٛP:�o�.K=��'�45H�r�mT�柛���ƉT�"\���S�Q,�e���9��M�U#�oʎ!���f�&#�0�Y{g찋��i���@�89�A���"	��?�7�0'r��5�������?zq!@m  �}�4�<����`@D��@�;��1kC���*T3�����&�mM�����n����i*6�ؽz�r��_���#��kf-ֱ�P��]L�l�0#S��j�:屶&�b��bB��:�p��F� 5�	�Ҭ��B��Ƚ[k�(`,�?�b�:	Vaaw<�X�pS�ʕ+�6B30ҳ��=��VK���P��>��';�>�E���5+cg�/b{��͘t�^�0@��2Qf��2��Y�u3[Uؒ���z�h��@�Z>�ܞV7��\���j��\���s��0\�Cc�5�����n!Lυ@+�m�\����U9��aO��(u���՛��{���=ۤ/�m�>{���_zq��K/�Mm�h�L�.���z�X��l��-L������j-�'u:V����ӭ��_��{WG��e��~��?�Ý��;��TU;A�/�tҋX��J,�츜�~TP�M��U/��)�[4�Wǡ�!Y>A�G�u(�ߨ���3��(�	2(ǍC�R婢���K�+,A	'�~$g�Q1w]z�^5b�)6�֌��6}�\_D��{����f]ןw�8	��.��o�-k���t���erh�����{�a�����]�=�`"���&��Qˇ�~59�m��^��^��q�+X�b���]u�˖BP����+$F�*���rzw�5�TO�j��M��O�]]CS�!�CLL���$}�n�Nni��E�D�[*��8�l��b0N�)f���U]v`���垚��r0�%���p�  ��D�f(��55�%X�}�ݪ�/���ZS
:�������ޥ�9ұ=��ݸ���q��Ņ5��ID���ؼB�#*2����#mN�7�X�� � \4��u�o���I[CM(l��q��CwܕF����}�u��m��H[lS�&��� �ꚇ<���Y��;������
�T0Gp��/τ�JЇk��r�M���.Sf��6�eKI�E�"2�2����yפq:��"���E�G
��U$���� O���"�2�X#��B��&�� �8/�H���4X�@-q�_�T�0�f9�V��>�������y�_�:?w�ڣ�;4�e2�:������0s��_I�ź�����3g���0�,.��'����/������ps[ Vs�[e ȵЦ�ǩ��&(LЍ��u��U_]�O'���ban���������g?����c7r�����]��Թw/�5ok*'��:&�H� 9�S�"_�|9֮��� ��4v��K�8��[��k�s��N����#���ɓ/{���$�fG/���Y2��$?�����̅��y��|��y���P	N�U
�J���CӢ���4 �;�c9x M��h��.u*X�����Ԃ�2iP��W�ޫU��|�L���0��昄���l��$�rS��v�B�����#�0���� ��Ҳ �A����-���u�;k�K�1��$tI���!�z)]ʘ�����nyt
�9�L1ދ��ՋWg5�,�œ��)�4�m�&�i���t���������o	��)8Y]�0[�*$o]�����{�ź !!%eb�-}]ʺ@цlD���	���3_�~�$ӏ!<q_�i���U6�@Gd�����
$ˁo�n���<���V�}m�?�oJ��U���䁽itp�
�z��#[e�86D(�ׇ���.g��8���� X:69�����!etNkP�bΰ��E�%���
@�FL��h�S�Q��� (��)+��	��gY���@� ֊���	�~���`.�a�x��t-�eNzl�NԵj���_�X��?�A��g����kg�"l�ư ��F�p��E둕�F�qr�S�\^��xy����:�Ǜ������������z}��ɩ+��4�.Y�@/�����@a�nd�叚͍���b�=u*mJq��c���w��#���{��������;�n(���O<��W��b�����C';�X�X�^�ƭ��nPQ�ОR��5����bi�r���e��t{��(r�+�)m5P��9[M�1��@&��z��!-^�@�i˰ �p��Y�s:.ՙf`��5��w�x/K�;��g��t%�hGw��A�C�R��,J0��z��l3��;\-��_W���.���~���߭��}��w��������+W�SC�oH�N�11H�qc\u?_S(�P	!:�X-9�����ѯ� � �J�d��^ W��e�^98��'�BtU�!�\��ظ������L�;���W%�S �*@�B��M9����@�K����I4����q��i~v�z)@��� ���Rd|�7WР�+ԴSW�M�]�{t��]�>7�l1�tbTsDc֣�u�&�X��\Xн"�G�Y�B�=
��Vaϡ)�ɗ�m��uX-1B0*�T�]ieiũ�| Ƹ��<�P�H�����s�q��=ڠ��F�2G�N�2����;J7F�u��X^ﳸ���H����c3Y�q�@�!Tيg�Ws�pd��fͤ�1�d�i�gf��?l�� ����s�'�rdm�g��ҳq�`��
��0e.x���v]a���J��Ԭ[S���M�c���~Td��̘7Ed�a����kЦR���
k���^�xׅ���Пnh�l��������կ���wv�ٿ�MBؗgW��mnJ<�F��[��Ȁ�[[���fkx���v�|:����8r������|�Y��çV~������K��S����������Y��U �充��_��^}3	��3��עm];�*��~fg�BN�M6�������,���Ԧ�yuo�������a�e���9��ےC��E��\#���+���8��a�[�����Ph(a
�[�.��|�t���t���ZT�;9Mv��zۡ�q�P�$lA�X��H%g�L�$r-�-�{U }E?a,]�>90 �-��:.ߛ	r�O�&��� ��J�._��hٙZ�匨��y��ŕ�:Ir�j�*� Xrw�B:h|�1��:9��uσ�L��{o�����43;�ώ��4oս��3���t�%靖�c�СC�J
�ș^�$�K�s�2�]^Msr�;	-Q���uC�c"����0R��u��J-=�ȣ֌�`�ˈtS[�FM4�!�]��bb�����!����T��.�mb`� պX%��M�T�����S{(�B���u�8ӼsQ ��f0]�z���u�
ѷ@���eؒG�!B�U�	ז�(��G�L�u�G/��@����C,��h�4�7U��9�s���4{��_'9Aǆ��x�N��F��:��C�/����#����t��c,xh\BA�D�i�����8�`#�fԵb�<ﳚ���]�_p��!9���-6O��ļnT,������H��F_X"�%�7`��`S%$��o�N�(h�����ϼtjߛ	�}��M��߰�1t`�>���Ƴ.�*Ҫ�R�gYi�P>�{k��nľf%j������zm�t[k[�\��z��z�:z��ܥ�?�����W_|���/����c/����=�5Ϝ��]�+��.IMH,�ey��A��0�p�+v�!y�n��&�푢�ȱ*��{��5��%@�KA7�;����.��pMN�`Y5 !�
A�5��QU�M1D�[q��) <��������9B\�1q�d�hX�1��O�:)Ჾ?}�Y4���1�(��% ��sx7�Ε,)�'v��!2��˸Z����juP�g?���H��+�p�E!��PKH`gPi��r7$�~��w�xG��G?am����L���A`}��ƦT�&�%9ܤ{��Y���k����>1}n^sO������
48�k�SH�G@qU�G�����2Kb�����ۗ����3��+�=�t�ݪ��e���#��cD�C>8��b'fu{U�0 �yhj�$2�z �-�E�ی <x�kl{)��sN��7���-�m�2�p��b}:� �T	�����vauU�"}��`"�ȨD�>"�&Р� ���+��d��F�a�*��ӛ 0a47�uȁ:�0��6�Tz�/ ǈ  ���Q5���`�(��ЗXBh�� N4i�/�{��y�#,u���͓Mh�gw�و��� U�
GP���:��<+;
�}�a�^�f\[X`�8�`������*$�s:�ԋ�.�����9�������S����m�{��w���/_��n]�ҕ���ͳ��_����^n�ru}���nÊ|m�(���
����\�E���( ��Ya�����`s��ٱ)�ܯm�v����ty���qG{��]_�¥��w^ݜy���w���G�?�y�܅����/�����R���I�������{�7�Kޗ�A��! i�Ԃ(�Eتg�H�4� I~/�6�P���}n��Խ�&�8]vt .^���6��FM٧��V 28#��������3�Q��R��Q0�U�Ē(\��eP�s\�����k!ޯ:;_���Sȭ�Μ9��^�p�@�;W��v�G����c���n�W[���c��iF�߄�6u~��%�!?|?�,5v��ջ�p�k�ȹYD�#T�lU ����4AZ���mͫ�Z� ��_[�2��Z ��x��쓘�k�:0b:>E
�)`�莾����*���9T0׻���m��B���o�٫�g��x�,Հسř�tE 
!�18�3�O�����I�ti �^a���؉q���Z��I}��3�
p
��oِ&��~t��I�L�&���� ���d�l�<=����Q�n��,�� u�4�\t�&�)`��qm6�O�1���4(0D�!�!�nB�͜D<LY�Ua�k���)�Ɵ��^Ը2["�d���˳�>���^��#�/ؾi��\HT���	����*i@S{��ƭfh�C��٭B�yJ�g�}�-/�EU�� |�wb�`�)�1��B?_ ��B�CH-�������[q�g�o���k䦘�Im>�?�*���}� qQ˥3xv	��xΜ�|�	��LP~���H0�`���b
�CO�r�;�xF�p� ����Ͼx��l���t�*KG�i]͎U#hKu�J8���[����i�Z]Z�������DOtO8�٥i튺����~�l�볏�|�q��~�ѳ������_fYZZZuy��ѡօK���]��/<{��^���/��k}w�M��C�.�q}�&C�#9;z9�G综��"�[ٕݫ���� zQe�@���ȠK��H��%���[HѸ��DÄ�/�n�]���^9]8%�';J�"Z�I9:�t�v�rh}��~#��! ��}"�$J���/�O�iT���H�Z��HM����U-�����^�i��q�)�%�)�(����n�����{t��n�)]���0�ːj�cg�V��|I iXί��7Ȁ�C�+#j�H��>�����Ki��ai�4
`Ɏ���}���<k [r��REZ��@sd�Bx.�h1�@Oy2�hbz���� ��YW������[�#%d��Vh��2� Y�
�"<�S���� �`�cj"t@-R��rB�~疛oI/>�\:������ �/;���Y6�FTǘQH��a�%�f,cM�l
1�j,�լh6$���x�)(�j��a���-
X�	�.�C�HE&]�lb�r������ƻ쬪�{�S�R�{����u85^ǣ��xW�I ���B��7tx�kI�^P\���� �M�W}ֆ$PG4Ӧ�C��l��#G��e������GR?�TU�1��EB�+��f���8�D�+�a����P���0�{��E���[@v�,�̋�Cb 8�72��[�!<��<4E����9B�6���nȎc#���S�>�G��~~�G���/�n��Ͻtf�?|�_s���w5}��m���'���P��(��߭�߂�+ ���Rc��T��K쌲�Y��ؐvt�[Z��n�觟�˟�L��mǧ�>�w�5�SF����։ڶ��陹��/^�������zsO�k|O��d���� ��j��UP�r��71��U��k!�p
y��f�m+䑛��Fm/�G�&�jȚ{
qy�J���q�uQ��.b)�ʢ��ށ@uJ hM�A�4���ё|���8~v�%4h��uEQ���Y��an�Vt�9�1�o��Κ�rD�����m��:<!G?R�3꠷������i��&�_�u�`�E8eP4�ژ��E��;8��r> �6a�q��M�kn��F�K�c7�<S;�P�����*��4.���^��ka�t�ԅꧾJ�o	��6:1�9��0�Ì:/����(dCas Nw'�;1!�e�\������c0 [b��*7�`�j��1,ئ܂�Ԑ�9wu�B��������P%����!L �J����K�|"s�7��8�2<O�c�l�y4�7sbì��h�^��,ӳAq�,%�ܚ��{�
����*�H^�bUz�74n��1�j�W��P���~O�<�8�p�N�����s�Ⱥ9�j�*���bߩ�f}U�D�N��c��}�{ҧ��P����κ���[N����t��e�ߓRާ9�����s�L(�[�d��q��% hvthɠrU��}#��w��Uq~}ܫ�C1ǝ$;�ݐV��. ��y�r����[Ͳ���	�[-(F+��C����ە�^���0SS�T�y���g���_���+������B��S_8���#z╙?��8ᢝ�h�	�������S)�Kw���z�X���j��;;]���E��F�9��ӶfqqV@H����������j/��Т��Š)jޑ����-��Ԋ��58���%� �j
���&��P��m��HD&)�A��a��Uy[���k�%��r���&rm���Br���h�A��� �ɉP���n�2T��Q��sreI�Bv�#�ͦBAJ�v�m�1�PMyU}���Qe�W`lP����)M�:��!���p=rN�>�.��e8s	8ӱ"<"����@�uK��#��R�ՄuPE�n�*F�������j�s�V�, �F
��a�
 ���X$ݶa�1���k�JӃ�"����;�Cwݞ�z� �<�=�E�V8X�`n�0;�����#P����f�r�NQ4��!c�0����Q[F�l��d¹Ѯ��R��[�@86:��t�����{��w���S< 7bu�"3��[�ǚ�քlҒ�V�E���b!��B��v0Sݺ~����=W�/���s�p��!�?SefFsJ��� ���M���t��8;K?��ֶ��*L8�1fR�Uf����0�!�ߖ>��f
O�H�����mVl�����
��N����4���.��l��i:ΨB�\�^�fk��!��C��u{�G���{�������<�������r9Z���|�'���`\� �>����P�wܮ�E+��f�B\<����d��b�=�^��YQ���@�l�Z�3N�s��f��0&`��lP�/��4F�W��'^�x�;��~}�G�#��?�'��f���o26�?�4��ǟ8�����詗�}{mp�N�bִP�����G���Z�y6ހw(}�X���)�5��r��[E���%�a��K�,!#i�H	��V=.4yZ���%���$,�&���f!�3�����"�ϩK�{ׄ͟7�;l��D%H�LU��͒��0 �M-��*T�ӭ����N�u��3`$X>��I��#�MιWkLNAj�H�k�f�,�d=ձw���a�v�vؤ6k���ظ���`���B`4 �F�@�M���h���qU��-��5���V5"�W$2ݡB0�b�&��BK�8i���8�
68�jEa4(�=����)��J��nK���+M˖2�`H�����G�gj<�똿��O؉q��xU��;�X�ʳ��a��L�
�-�w�
K�J�C!T��p���7t.����W%�������0g�*���T��R�]�>X��]>sN�D��N�c��)|6�N�>�fp����P7�y����׮^1���1H :a:�������b� �d�g:5?��F�
MY5�PtR$����p��;��M�kM�)�Z��6�j��{*+S�ѷ~٥q#��0#�6��'�ӽ^R��3ʜ���U"aX�V�X>3$ 5,�CB���Çһ��٧n�'MپG�}Rs����<M����o�`���H�H��]ߕ�x���_��N�Ȟ{4������\���10�^/`��/� �� �Z��n�� �C��Ue�e�b]���C'hh�z�^O�iM�D�
�D�z�y(|i�yLs]2�pK]$�<�~q�q��*H �������\���c7]��<���w?����}�C���=~�������Z��v}�5;7ףJ��Y�/mn���|���ϝ���k���&w��u��7��Hg�iS��R��Em^Ƈ`E��z��|���
����I�qy�v�n���3�I��V]��V��P���������ve��q �}����M����dQVl��4����ܪ	!�v{<�tp{R�go���oC]cqvb�@�5�aW�_�>f͌Ő,|�k�R���?�A��{�43��F�ێ�:;��SS|8�G��h;�$T��}����#��	-�	c�1��)��1��BȶbJH;v�\��y]�������_\�ty	R)�뱨[�G��'G�PkR�	��F���!�#骄��W�l�!՟+�r���v����ߚ&GG������@�,�ft\ q�@Ì����u1(4UȆ�
C�B!AtXb>.���Zz�q�'����!������ 4E�CU 0���uT������ �#��"m�����(Ao����F1r+��G��Se����6��/=�������'���~���/������c4�� ���#K0|&e�kT7�J̰_[�W��E9�TB��}6"TC��ǳ��>KU��Й75=#�<0O��L뺄�u�fkn�q�m��<d/ ܟּb<�~ �s
�ql@���SW�?��e���GD�K���ӫ
�1v�.�"S�Mڿ@1��*[����;��/��/x��]<{&=~<�sN��tt�y�7��Ok���ؕP+��
�m�؆ ���d�w�D3Ã5`-yV*@��5<���E?<�4�!�}kg������f��3�C������F=У��Aj]`N��P���t�ۆ6?C�#i�������S_x���/���-�/��412tq��{Y�9����_�z'ֶ���Ӂ���}�jh���z���#�$�k�	mh�ԡ���D�ʁpP���&( �Zi���ROR�OU���kI��שJwۢ|����C8��5i"�{G;"��m����+���C�Bq((*����wMo����r�G2
���
���o��D;��r-��a�X��q��íBYd-���m�[8M�O|��r�E;W��]� ��)8�7��ǽ��̈́$h�J�⊲�S����a@��~-R�?�,�*2']��3�tk��.**6��!W!�>��7xw��w��ܣ�e>|"���:k���+N�)$��g`�X|7$&}��5�4�b!	�j��.!�gD��ij��E�����+ 37�=w:���}����dﺄϑ^/!��:�ώ����ү�c8ɵ�p��38vv�%�Q�6$�: F�R���z\����)a=L#U�	˸E���w�}Pņ ���MM-a�:���/_��&�����ߚV�i��x<}�[ά;�����C�/�ȏ�����#?����F�3?�����E�#G���cH�N�-8�m�7Y�{�x��x���"�QsDv�w���;xPUR��v��_`��KEl�w� @U���_��@}v��"g����qL��[��[�G>��Qi�n��v���<ux[����fc,u�[�X��皀Q��306�Ω8�ɓ'U�aX!�=b�V�z@�$�x�4���j�K�ږt�9����b%���P��N�E]T���$JB,�� ����#�N�R��Q`���j����5�c����F�����
��i-���Xd͹w��+�Ω�Lm%�{t,6	�kZ'���|���0�59�n�=�|�Qe?^M���B����g��B�H `e_X#4}5٤wd�Ca�	i�&^��|�٫˭������JmyeY����>mV$$�JkN$jt�Q�:��^'ew�?��zV�=�hú(OZ^ot#͂е���"ւc$�H�|l��x�q�#W�_�B3�3���C�(Zv����{U�3���K����U-�v��?{{#��k�v�.MO�X	=��}��4,r�Ҥ� �]8Q� �%V�N�]ZP��H�eEK�jA�#�\���fP\0�q��:� �/����pֺ��%���Dz4U������^�h9��JA�-?f���%'ֽ�/�(|�0v@�uZ�F���������4������+�@v���e�N�;�I��.9����O_xQѓ�%���чK�+�k*[`��x��=���`�	�jQ��`�l] �
��(T�ۨ�6�����)���q�Ua��0�d[�Z�7&a��b�L������.�z���~]3�$�x�%���]L5Zq��E�� �%��:9�}�t�=b�v��4�THqD�[N=�E�tB�k���Ŵg`8���黾�}� ��!]�~?�J�����k�腆^��6#�J���6��e�>��O�6�L�qe���Z?�����eS�aCs�2�C�أp4Yd[ꃖ�����:�������O�TZ@޻oOz�;H�z���=\!m>�˦�����Q���i�� �L�Z�RqC2g��Tl�@tՇbp�;�p�E�n[s�3�(���X��e�>U����U��=`ʤ��D��}#iVlO��-�-�_�L�{�i.~���(ݕ~��~>�]��z�[��a�UϘ#�$5T���Yj��㽺�a*u˾+*�@B����J����P@����г��u��1Ӝ��<E碤�;v�q�7�<���s 3��\e7j?����M�r[4����ξ��eK!C4H	81���X��.k��jy��e38D�����w+���
���fCыSr'��@� +��C>G�H�"!��}����^��ya����L���E��>UhF�H� ��P�충�B��.�DMi���E�"�#�^;n QU�gE�2炄�iȜ�E�:�j�ǖ���X������g�B��ٖSǗ�P�`p&�ۡ�{�q�B �b���Ҏ[�ƃ�ɠ01���؀��%�h�9%V�N�^ՠ�Q��bǉ����t;r,��K��{����Mkr@�I��U��Bs�!<�0r4��I��~{�h��-?ܣ�
b�X!&uF֍4m��uL
�c<�w3U���3��y'��svZ7�
 �<R�`���&�T�|���E��c�P� W��a.IɆ��r//9�m�GCW�W��2FT$tb�;]Z��{�x�B�b�ݿ��i�����8�#��7Zp�۟hr�O����������N�jc
�mi<z�:�g�L���!�	l��k,��@8�K�<�P*Y}.PIͪN�	1v8{ݛ��%�:>�%��M y�,p<59��7�g>���#{'�J�2�X�M�f�3�M��9��@V U��}�7ڒݩ15,�熼0pKR�́/Bl��X�O�n��MR��w]����V��l�;�i��P�ĸ�i��yN/��y~/S� �K���w��xK��ŕF����*}�S�R�	���)h�A��c]``�& Ê�:F�\x]@�j
�\��i��g_Nt�Kk�N�"��=�&[�����7?���g�b�ٺ�P����s9��W26v��
c���ye�:�#z��n�_�k��$����d��i�ƌ���
�Q�b�����釼	����|��b��nl�x��2����??���y�����o�V�����{/ �;_-��Z��+����E�aBX�nm�`�i)��8�/g��"�$c��=j!�p���.�n�m�(bs�WHyMC8?t1>����]�'��ӭ�#������I��c����Uw�!jȁEJ>�M����)�]� �4�u}�
S���܄ T���rP��#
mP�fa���Y38�#���gt@0`��I�p:q�z5���w��G����\Y��i1�7���P��>ir�q�r�b�?�}������,ׄ�c  ����\ǖ��9u�:��}�^��Ħ]�9��Y�#��#�˂e��|~Ga&*�l�س3-\&4�ݵƆ������bm����;Q&d�x�b���>�������7�QZYh.�Kߠ��(g�/�G7�����t*�l2j!Q`@� Ӳ�#��S��^B[:6��v���(j���&�F�} f4w�/%��w�l:]���ۤ� R�歃�w���0c��������A�Ic@}*� �0�#mK�#ѿ ���u�z���N�G����QL���^�/��M�$<�-����Fu\���U���316,����;��)����lBD�����tTz��Ӣ����?�>�ɏ��S	
6�\�L��B�� �QK	^�ƽM�'�L ��Xy�����+:<�]
�څo��*9����VʆjfQ���t�ٞ�^?�̎����Y��τ�d�pi^*ɀ���b����#�5Bˇ�lS5t���P8���Z��	������[��`��nly�ՒC�a�[���A���f���倝׻��R<�;Y�p�|�ز[N�L"hkJ��f��7��� S��K���X�U�5�q��r�0Idn�c�y{���GU�%~X���-��8�馐��:ęjERA_ b��� d����s��zA>x���Y̨��ҏ�M��z;UdN�	���X����A��eǣ��K���R}���p�8�9���hx\���k�I�%ݚݤ[�Ȧ��I��9��֨�ZOVZ��Bf�<�v�q?ts�4��l�����y���i��ElN���zE�����ލ��Y�T���@`ѕ�->W�E4%�#(<�����;��u����l���q����9�9����	4�]��;��[bs@eS
����%6^iu��#!��N��^�@�}[ N)����]I��@ˉ	[��iga�,���$���c�-��"��P�pC�7�
0�!�o����fz�;ߙ^y�e^��, Y�g��S8x~i͟!�kR�9��4f�}��J�M'z&X3�l�
�~�7ؕ��W�Ƚ����k%T��.y��h��j������[k�n�1D�E���*�`K �B���*�wHn�>{D���[
�1v��`t�[b~�._��a�nI`�{c�cG��(��x��q;�*����|�Nic0�q �![�HO�K	�I�@�'p��Jr����*�S�T��:6��C]A�Va�j��F�.�X6a~����:���g�}�h[!8��"zD@�((�c�JB���ࣜ>�ETscΡ|��a��n`�x�[��(	-tR��H��ubb�U&^���o��Ui�o�_����@�Y9Z�W� ��	ƁE}YRT��U�R]�(�n#O��$h.efh׫�&�+2��1�|�j����S�0 IH���/�,�\C�
�[ab�u#J��AP��Y_	�H\�
��n \�cO�p_C�+�{�= �Hq�����PX�;�M*���ZG�Цt���Bg~��qũ��Td��g����0 �r�M5�DD�����Q�ٴ*��C�K�(Ш
F��@�)�+�}c]�D�;�ޏ`�����j��F��p�a��ơ.P�!;8=Z�min5��� ݒ��k��Xֽ����n�д���f���}�I��ݷBH�
ڮ/�����~^�O>��3lV6�R��tVs�c�=�
��J˲��y	ʛ��(F��9���ngGV�;�H�B����s-Oy�7rO��+��ԔTP�¬�����9�9�p!��t�^��9��QAS��W��{������v��X-TY\ ���KU�E���k4��(��(H�z�'m��XƁ}ҙgt-l(�R�#��F��~�S�%����Q��4x��y���[o�5�^�v�i�y}?41(���A�*�y�D�$-�E��F4�������WU-}%�}�-�c?�yN "|�%@��z�E�hj�Q������2u�^(e����j[�c��L�U�9��u��Ɲf����Dk8�B5�X'�>�M���r]2�����~2�i�b�Cm)�3F�\N�Gn��9����,�fэ��.��_��\����r( ��L���'�;';0����:���[9735~h_���9u4�Ĺ�|8��_�f�����I�����d1h�;|X��g��q	)������i����y2�^:yF�W#�w��2rX(�q�,��	���>-p�C� U@����&V$�)�J"v߱������\�h$�T]9���hT4Qѝ���v�P�M�����ٻ���	fڥK�)�,5sQ�O��qF̎mRlqbXH��C�0�ZC�~i4?��f�uV�BϙE�	��}JQ�`��� �����hPz�����%F!��=F�B;���Z+-�{!��G��HN���f)�,�j�G�Ύ�GST��T��˺:g������p��h{!' {��ձF^�C�3}e:X���zo�[Il.��P���+�J_C�x]�Ϩ�)#����}>��گ{XT��`o�B��:.���zY���E�D�X��QhJ�X~��b����'�dv�veM��h�� ��=-�\ �����:����Ջ��2тD��>�o�8�,V�l��V �[���X"|ZS�.	{Ra ���b��w̯FK����E�(����^fP!�G>�Y�T�)���c��^kҢ��_(��P����,ρF� ��B���/C
ա�!4��� m\a��jt[�q����׻G�	�5��f�N�p�rR=��P�˧^I�/��>���N�������a*�ܰ��Bx$i�%Hff�M"�Z@lN%!K���yC�َR���^��"A���z6�W�n6ȜU!O���zl&X�Fp$�nj�p0m��l${t�x +���C�\iz�����6�Uڿ�6���%]���X,cc`Pz'/�:.���jَd��z�X���i=\�8(:-z�`�����Qv���ľ�K_�3?�b��8��x��xe ���gr�_��o��~�NO�oC��[S���b�~��φ*�6�ׄ�dKd<�
�\X�0r�����#ZMW�5��F�E��3�`bKء�|��6;�j�=j���ʙ�RR;�4��������t��iD�r��I�J횮Y�4 eX�7��H�s-9�%u�v%[3�g�~���\������F9$�ա,�.e��G�P`�N��G��um����vP�4�������P	Z�B�F7�D���!���"0��Cg2+��sl�tc]�C�
֜V�v����BX{@��
���K0U�:~}C-h��r;��t��R���řn�@_-�X 4@�Js�{�17P=th_ԩ�(��}�۰�]-N_L���)>��;ӿ�W?����ȭ7��'�����g���c����n�Mb���W����~�sk���H�0�Jc�!��/�x�޷���.�)�R��^ENjQN|D�έ֪�?����	9������/�ZtK�Ʊ�nN�}�{�3�>#��B|�=��r	f]��Wl^=�x.��.��S���j0"�`�X��å�CU�yA�ې0VB��ѯ�ބ�O� ���8b<�oT�R�w��DH���5�,��Y!קIbM�dW~�:|D=�&�?�ph�����ds�p��t{b�t�>��e�����C�.��N���-1���ZP�[���ҽ�1@��3��W�L�%��q{���z�"�I�ް��E-"���6I��\e��	�	���K�>ܣ���wަ>{W�yղSA��=jƫg��6/��0I'��
6�)u>K�}��ҹ��������^���4�T�u�g6�޺Fo3��Z�!�\E���6( ��:�ڠN]i�".���F����x�}�� h��(�ֻw����Ϙ�@���(�3(����;1eCF@�d�@�*��ЎJ(4s��������:�g�P���pگ]�ჇҔ� ��A|K3O0#Y����kYRk*a�tb���*�J(��E��ǟ4a�FH]F�����RD�4��n��M]�95����S��L�K)�aѯJ4���]�6x����Wt�,J�k_���}��Tm*%�n�t)�4 �=	u�I��룏�P�8� |��\����B� x�~&pJr��V��ϝ9�{YO���S�6i�;륅(r������΁�\���=�r�83eI�αp�##��������P!�5e��f��8T��fB�a�=.� {l��:sE�PHK�������O�
ǜ>uQz��t)��Z�VbU��ȳg��s��O�����l��?���;�Eao��&eK�N�
=-̥�g.lq�Wԏ�:�11M�.N��Z]S8S��Bt��9b��q��iR��Qm?4�hR�o��؈�P��9��4�=�"�S����H0��i�M
\�m(��*��²6�Y!�%$yYU�����^	ꕄ �2/'���z/}9ds�շ��	9�t�U�L9���m��/�=Q�0V�b=[ڌ�h�VUoHa�>��}�d��ҸB�=�I��C#b�$���;���	ٗ.MO�g$=���\�/ϧ�E �4z�>����~���vl�\b ���1�e�:֣^�l��kda기pu�n-�8�<��A������!{Ϩ��d:02�f4ޫ�
e�l°��t�Z(�Zm"/`��N�l�;����E��d���� g 5�z�a���5��[E��6/�z�>?�\D��[��� ���7,��Ǘ���r���bވP:���p���rwx��h��Q��#.�0b�F-vBQz��lsUU�U_�S���u"��-�K_u�A/�dU�_�@C�gT���B�w�P��޻����f�M���-�d']�4m�r��-�v
΍�+�t����2��I�:��`2x��㢯SM;�&Y`�nX���K�d^�t���wɡ8Ӱ��nBB���{C�u��]w�)0�ߡ��.�/�2�A�Q:�~L�k����8 ���[^ZM���:m�nxV����r��K��F�J'r�a"�����	�
�d��3ϼ�z�Ś��MKk3>��@�m�S�e���h����h$�}�b����h��:�S���M_��Uꢎ��f9�G%Խ��;��
ƅs� =v,-�Yx�;НJ?�o~A�ߢA]��]~ŀuB�=��p����ӓ�=i������L���#�>m}՘��q�(�p�4#����cj9|p��Ƣp�2�>��OHܮ�Ld+"���#5{fTaN��������/��
s�.�|��~0���gĨ��kr9]�f�P�=#�R>e��!E��;Op� �7h�ک{�O]]ivA���ae]Q��܅�tN)���Ǐ
�H#4��ZLoem1oǾ��t��^����(=����E9�p�knf���H����`��O��X@� �p�0k�#*k1��Ź�E�a�-��+��vҾã
U��[WAL�^"ʔ,����cK�c���H�g��/h�#�G�<7��Ph�������@��A��OD�K������0��D�^ �na��:���֠��1�5r�*���ޢ���&�6���������#�{%tJC�H�<�Z	������D�ȶ�r�4C�E�#�lT�Hk���=K�k�ֹh�����r��p壿�,P@�F<@�gAU�d��Bp_Ʊ_��ˡ��;�, �d]�f��Iņ�q�j�FqCv�0A�/H�7
�,k�S��_�?�wT���	C*����D�������Ϲ�z���W���Tz�v�6~`���4�����3j��k��t�X��'o9�:6{���%-����s�������EU�~��e1H7Yw�͏�8�p�L��{:�"�,�02�����4���~����s���R�ȣ��tn�ً>�1tQ@��^vcО��t,]����M���߸�w�r�O<��Ğ#i�7|cz��g�g?�i�3�^y�q�#��t��K�������5��ܼx�T�]ɬ0�=#\��yF�����B@�鲪2�t�tD�L�������ω�9cVbJ�Y��G��/�w:�!�c��^��s/������t��=�2�����f���y��xN��}D��ų���}Ea�i�/�A����R�d��������О��r�Mi����w�!1�z���B�U�>���d�x洳�p����E��MX\�C=؃�n�%�& H��9�6����^v��;n�-=��/:����':�%�)���L�n���˳��|N��a�����/�1O�
����3k����f�&^��"�C�����l$H�Ǟ�<��Э�{�=i���mب�)wl�pZ�|:���K��t%M(kk|r��g�{�!��=궮�K�#���i�BGp����_5�Tn`c����^���A=?bFHP���͇��ҵ��ɢ.fߖ�[1/��"/�~A��A�N�鬧[�H�|����
��.�
�c_���
dV!@�"���PԪ� yV��1�.����iI�NՉ�;��Wl��7����~��P���0�a_O���^��o~2���s*Cp ��_��tEl�O��_�5ϊ�����5�E�{�	��b��l�h� �p]n�C=0�I#���%� ��>;�^1�N���3��V���md��n`���S�Tw�U;34���5/��
��G��i���5?�o��'S�|u= b��b�9K�
�� !�"���ҀH,�t
$�@���-���E��&h$�j
�I��"6��wh��u(Ty^��KD[v���oI�	� ��$<ݯŐ��+�O�a��{q^�刾�;����R<N��u�����=��x�&�b�Ω�����E�>,�1�rp���M��=�,��
q�X�3�+xS���<:��?�ԓi��@���ǟ��q�^ph뀴)�NZru1$'t��% a�}��z<--	<������$��F���*�'i��Y�.�M�4&�O�u�E"�[��_T��lE��K�EM��7J_��w� J}^���M��)ܢ�0N	��ē\�	� M��(d��4�N9��Ys������{���B}���뜯�������ޔ���ߓ����#E/=�����KgӃ�zH�t:=��z�	��,���|L�����Oֶh���?>6��҂f��#��^z�Lz�����{�I�&) Im@L�зʾ�� w]�gK"�=���8}����:A\oKs��ԁ�'����Fk���M�y�"�*6���oV�W�ןx�	����u�l��E���z�g��5V��ٯy�{ҷ��o���!fQ��=w�cG�X�{I`��[�������Yb��@�P�r�T�Am�W�bH�H�t��+�/
|_����y��&ѵ X������{U�u��%e�Ix|e;�����ྃ���~�����z Ι�jl+P��x(�T�|QdZ����X� 6(�9��Ԁ6{Լ������d�� ��l)L!�:J�k�k��Z�s+�,V@cq]�IkG��{S���7L�����A��][���7���tif%�z�X��_������MiN�8�7���̃>�G.'K���zk")��^]fCKZw����%�ޛ�'�笣s�X���G�/g�z�|����x��@���<����?sq���к}N��0�X� ��`gۭ�����X���k����
Դ��J���u��3 +�[2,���X,*� {)6C �-X �C�'�'W��J��)����	�
�����f�mA(uSD�;kI��H�GT�b� �!`�*�Ǌ�-�0 X��[p�O�$�J��q�|�^�/��iPo���d����Pz3�\!��܀վJs����B#B��S�-�T�L97�|��
���Թ��[n5�N�����51���̬��ȴ�q�Ȱ8�U7s�"�%SL��$ȥ��Rck�g [��sCL�\^Ĥ5�	i��&��p:�>��1�'�h���U��qF�����N�O��.�� RJ@��t~�{�������(���'u]׃͇�A���$1�£�O�M8�= M�!l
�a@
��pP��4X�;�R E�h��~��#bY:�A&G��hs��ü��d	*�$�̈́X,� ���y[TH���Ɗs2g��% 
�}2oI�� ��ӽ�48�h&.!3�}L�1�E���Ze6�c�Ӣ������ �5 ]ծ�ܫY(��W���*��XX�1'��r����W0S
�!���(�,�h�0����#-�΂ަ�cQO�63���h�*։g�J�$,�=��Ç�:;�)�Af�������~�5)��6�������F��-x.�A���(�U��֔	�-��.��>e�W=�K
�]R�փ�'�50�����pz��l;v{ZQ�vM=�ԯ�W �=�JenlS�T�K�7n	�4:��LN��|HSE&b��6S��T�-(�"B�h�A�.�G�\��l���~����w��W߼��/Y`�/�"-P��V=JJ��nzU
�I������5�X$���N�H�]'���!� j���G��q��Wquj��?ґ������ήyJU{7��j(KpP�Z8K�}�C�IB��]�WBM�	@�{Se��:r�z��'c����h9�ye��j�cG:�P���j�Cs���E�Ľ��㡗�8�4m�USC����*�=t=� 5 (�;]�G��ͅs��TwF �].Α1bf��d��%��>�R9$����*��3���X-�
sىj���^`by�,����.07����G�u]8+z]�k��߇4M����5��P�5��@���&��Vz2�g����d���q)�&mz @aCYt��~9:@��3���2���bAp|� hB�3/�
��>����Y�V4�Ԉ!(D�B�W4PfJ䬸���H�<*�ɹ&'��"��ӂ�H��r����x�{���\fI���!���U/�<'�,'�y��]��͙�*HO��
�ҏJ8Y�9�{�-�<[��.Q6s����+�1"��Rr�l�"��%���w!�F #6K�_�a5�j��u�;����=D]�R󆐧�kc�,�HB��ss邴L�c��X
⹠�<E�E�Q�s\�)�rN���Đr�%�N@+E4؉��g�j�T�����E��zT!_����/���3x�-7y�_��r2bn/=ۢ�a3�ߜH�x�8���$s�RS�uv��w�s�ΦǵY |`J"k={�A1����0X=�=H��"�Z��� 5�Q�Blܧ~i�-������³���uI��ģt��d36'nz���d�u�=��(�s"�$E��u��%���o��nh����5�Ru=��SHVC�u�q�Y��P;�b�z���\�z=��n����k��:vCi0G�u�U,��s5�pL,Ξ�b<7;�n��f�E��iр��'�o��(��B[
���84�����/j� ���^br"B#cM	;�U�[b �  3N[6�D������j���M�N��jĹ&N������u�5 �Zd��ڽnlj��v�8V���b���%�?(x�Seg�u�z<UW�~��j�p~*2�^����k��rVїL�t��`g��Dqj�Ú����s��C������%q��(x^�*o*M��
�/ؤ7��)�77��@�_!A��4d�K�ӗ�h2���;�
z��jΰ.�۬a��6�+T6n�gB>���:2�)2�65\��N�*I/8.��QR!�|d��~p�0^+�WUÈZ38������cӓO|1���,�	]�4�#zb�Rd�E��q8kw���n@�ٶ��r��|�A��amqO���唙� B 5�{�5�b��I@��۹��k��3�g������و\��nXlд�ܑ5$[�9�֘qm�AF&�}U�Y�ߙ0Y'�k��V���3�ƥ�5��c���y���^_08�����F�>��%���c� �\7��;��.�#��( )J7Q��f�.������H���<?��ۯЩ2��i�;�7휺���J������Q��6�k�Ц������w?���z�K�2�6kß�=H�H�Ɩ�	�S8K6��P+�_iB8�En��Nھ�>�mK��7�I�!�Q>����#�]�@(@��=HdAٵ���J
;���/����z- ��D�e͐�	�U'Q��SL��ڑi7��L2���[>$'ؗ�y�Q��A��X�q �ä́�`Q\��d���珤WG5ޖ�a���������$`ҙZ��DNH[�B��V�Q̉B���a^�Z2cƂ���s����%�:}�;yt( *v�,�d��&{x���C	9B(-�2�U�F��>id�h��u�}��1' �� �Ь*d�]1eq�>�#��ġ�f�a�wT���'�	$��qЄW`��,���Z�G���7���ȱ	�^��ΰ5��`\�b��Þ,�A c��sƑ!� B�(s������CA�fg� �)I�
�ܙBUצ��D��=��l�������� e|希@����A��6�bh�{EY�̗��G�&�K�R�>v�(2n�έc �"+}Γ0�YR���ӿC��z:�(vP���ؒl  S����y`��f`Ђ�3;S=�9k���w�A0��ha�x~�!<�k�S�٦�X��J��mA�����u�6��L4 �eF�7���y݇�m
T���f�yX!69�dZ�w����?�ĵҎ�1䙀�@�M������6�>��������#?��Nec>��S����騴Y���`�$��iG$`��y��jp��Vm���WS=��{%�oJ�7�.�xg׺Z�4������1؀RQ������d�$����҉ae�a���7H���x���?tCc���ʊic磇hQ'�r(��H�%&O��x�Bȷ#�u�+3>�l^\�7�&s�����7��W�>9���w3ͯ��X�̈́��[�ܜ�������`Q� -���E��y3+��,�T��  p�cڱ���n�q���08ZO.�c�G,vktt�U�-��s�\�8ֲ�3�np����b�~��m�3�d{];� c��"���'c
_紨�j�A�;X�i�1qr:|o�O_�<�n�N���	sPtܫ[R躩��#ॶ��q�f� v�d�P�'�;y*�g
j Y��a�4+�Ыv�W�/�X �F��?)��+*�R���+'��������x�2�F�궉5g0R�S�0���/�̎R�N�ת�UP}0y����̬����U�!��9�j �K	[��+V�-j4�C��9���#����w '�^�!�M��q�{�h�mL���"�\���bg~�+�]tXp߯q> �μ��y��īR}��a��* �"�����5�r|7�����j	�2 �*�� d�L]*2�(�9�{��WWdI-W�{L�o�0�:6v�=���]��N��p2��Q����n�c@u9���]~�=�=�닁�d�	�ӭ�R�{.3/XS��X�U�h�O�&N�?��:#P��c�Z#�*��ܓ���V��ꏤ�nR�Z�^����������ߦ����tǝ7�����?}����G?�x���KE8�K7�h"�������9�Q��VsK�dӅ	�!��V�pA76b
�G����	$@��+�iS�±cǵ��*��x��M����3�^㕙�b^/t�+�8�6V�4p�m ���jw^���+��c�#vY=���P��agG؁c�T>Ο1+�F�솾_�BgQ"�%��?��MJ8�4#*��3���tt�'�=l�Q7��iA�,B�葚�G�Z�?����Q�/�!���\�J\K]L��������/�+Ph�B�	¢>! ��o��@��GE��ﷃ4��=�^P�'H���6��K�$v�f��w�jnݑ��� �S��\4��e�_,0�}#�� T?!0$��rxF��,�N�x�8Yvv�hR(9 ͔� ���$���,�Q\]�;h�0!(������"�=�e��0ЉƵnJ* [��D��J��s�� Pv��JC���*�n�j{Q9F(jOMN��q��z�|�"d@+�\\�6���95{W]3����A �h�g#�	q�Ց-�h��]�K`�hx*�K���ߖ�Դ~�V*� ��|g��+��QX��#�+𰪐@��I���_�5,篪�E��xƢ��������S��%�ı���9L]��-�mk^Q7,6��B(���(�#(��ϛ�̦�d� ��,n��4�k�1��CL}�=w�.�*z���1Ӝ��ZWVY?���--�)�S5��Lz�R�隵�.�|6�\:�nW�����?��u�Bjz��~,uJ5e�R��Ǜ�6��P�V��c���ּ����zMO�����n`l���ŮhH���[S[�!	�P�����E���z��k]J���g���Z�͋�w�U/���$�Ź��+��� ��+fح�||��F��g?����A��x�t�
H�����������u���ɱ�@�� 
���P�&��#�w�-��:���v�,�#����ET�p0-���x���]��+��A���z�+'S�;N��@�G��7������ٹh�\u;u��@}��)�������8 �1˃�z��~�M��N��2��Զ3mZ�XlQ�~�����A�
Y�*V��XTڥҰ�V�ɚA�c��]�X� Ж�{t3V�	���o�Oq /�J4��热a�Xo�{��Cv��¯u(g����fe;��`Ć��p��ꡕ�>�$����ju��^ )Y[��ҍ��U�ul;4H+4Q���|�!�Lc��ap͜ �	���������!?�=�3b��J� ��Y�=, ҂�zc�D-��
���Ǣ7�5��f"օ`� ��(�K�M7f��q�~���C����Y��<0��c"��7@�P�x1�
�m�S����W��k��䚂��S�j�bv5� �lx�n�!|�W���	T�q�/M����Z����	������2��z-�l�����c�k����CN���������/�L��o�]��u	��u�G=(h�K���"@�7�?�&]����<�dW�9�~ۊY��J�@A78�0�0r�������i���.,X,t���Z�a�|���ko�៵H�]�N0Cw`�������^	v��r�,�>�#�G�
����y�s*�����*�\M�k�A�׊���y���-�=/�i���H��=! I]Ǧx\�?��ԎI�w�R}�H�IKa40�:��]@�ԘZH��n>3`>2�B 	c;B�#Q��O�\*�G �:Cs'kl������gsp�B �
�Q��{�SޡFgm�h�ն�v�| '����3���}�Ҷّ�N��q���A9<Q1����_.�� ��k����>��b�pr�8i�� ��{:��񘹪X9dj� b�]dvˬA ��u-���GpK�,�������� %w��V�����ED�ss������O����~��p�\E��z��� ���sP1u�^��E�Г��A��9��\Va�G��?[��쮬!�Uq(v�z$2�"�	&�KZ�(y�&�Nr+v�Z�R:�8��(�����T]�5���h�|�+���y��_0D=fNSd{�06}�{%2�h��<>K���U�L��<����>���я}ʡ?qQb�g��魴Gw�T������ J��-F�v�*!�������O�gU��&���M��GT?죿�;��q���߭�PF�J�+s1�ɘ �h�<|M������x���me��nd���(4���ŋ�2�!�ƙ~ܴ8�v��A�������노�P�{ ��ڭ�Ʊ����N>����Ԏ�ÅAT������@����A(���S�����<D<�f��Wny7�Y��%�G��G���S���ZVZaG�%�oD���6X�lĪ���R��cf�q�;p�P��� ��[��"؃{qxR��wQ���M��C��w7�Y�>e�Iu��"�ܣ���Z�T�!�?����^�Vs֢�Nٙ16��|���<&U���T̀5` ��sTg'����a��Y�| 33 X�n���  ��z�TL�� ������!�Xv��(^HM_�O�
���J�gF�V�Tw�ze��	��� i�zs�߮��_�q�X<��N��
'�ōT��ܩ<O�;��d��
�
�G�*�/�\��/!t�W�' ��F!�T�*_`{��{蘢�+�J�(��1~�z��y>�t�O�; +%�9u��J�3Ĝ @Y=��-���~4h����۠���J�8�z@/�&��z�G��WNk�@�OT�����+�!�z�;�zS��U�?�$��
MN�ێ�ǀj)��gYa�Q��P������>����[|�*M�j�0�ޠ��[���0k�ϸW����6�Z@��]�<R'�X$a%H&D�߰��@8���ӗ��uA�70�ޟuA�y�^0���9B]��Z�w8����_��_C�gRi�CC���=�]��� �%�Cw�����iŅ�$�`�Wy�_�8�� ��.����E2ĴСu��:�ߡ�!�-����L��n!D���J����Z��S�A�����Y��G�T��E�AF 	E�2�tH
A0�S�T�=^L+����b ��lv�E��札�?��Q�$�+�fj��)�r:_ճnU>�!�D80�f�{��v��X��g��X� �h;�*܆�B� �@��b��k-�BQ�i�b��D����C�D��vE�b��e�+0��ư 3%iM������"C��P�u`� ���eJ4�\�.T04�˜EU���r��.���2���s�9�s��=8�����B۳��V�b=e{�tm%��m��.��Z�e`�Ƈ����&�/�b{i��Fu�j�dMZ:zg��s���1�L ���5ޤnU�N��<�z0 k��;����NY];��@g�l�P�]���$�� ���Kz��Ҡ �Z�l	,�m8:qo��{D�ɶ��k����B�ϧ�S5x���ծi����U�W;�餸·����Q�����̛�py^�y��o��/]���/_�( �؋�!2���B�]$R42��EeYB��y�*������^��}���b$�~��, }���xy� �+����G�%a"�s�^�ݳ�=�N�<�+�ʎ�k�I�C`_�E�(.����G�+R��y�v��u��B֖�MD��OX�z��5g��������&v���8\�0C*��r/5] �!���6-�Գa�cLO,Bh�q���w�Z����=��� �/�Ѱ?/��_ΒB��3����1��rbLpN�3��	ge���˘`[�2��?-��d���F��x�tXW�<�Z)������� ���p�<
��$������b���b-64Nd�p��A8ƃu3kU7�Jg�)L�k���N�ah�jNȆ��\ȦZ�c����+c�0��	�� �^�����<���_Fx2XK^����'ol�� ���*8����d�t)Y�_� һ�`P=���`�u���pb��K<`���W��+�Ɵ뭴B�����D8�Ў�an� }M���e<�ޔ��1Q��W��-��ੲ��"��V�2
*R� �=��	���8���e�9w�!�qe��U���ǞH��P�cbxb|(��-����H/����S���S/��o>���C_������>�ZHL��6�VT�r�[����~G��U6!Ɨ�[��D��jm�`�aH��Q�!�X�</�_�m[��[����i�� VO��m�, �Sv���wd����j��m8vw���/;�|��s��p���X���Ñc�X��ي)�n�b�u�e�}^8��[c�(!���R�O���ϸ�Zv�A���Rz,��w��L�7��y�ov"�ʐ5�� �0�=@���~pB��PΪWY0�I���3�Y0�/�uX�96�C��q�슲m��W��h�����0��E��"/��ٮ��������[#�6��m��Y
E�"�j�E8�T�(�3�xy̮MR'���}.��Dx�q1;���yFc[�	Pv�!���c l�K�ܰ��b�]���w������}��	��}f����a/��P�X�����7�RM-;6�X8)D�����z��쒾���ܬj1e�n�f8�e������+>����󳗻��>��: �V�h�0�+Д7j�� &���&Ѻ�HK��?�"�0����{� ��� ,��9�ˡ�T֨ut*���me�u�!�ҭ���[���M �b۹:{<[�R���������Y�Ϛ��;�����U*����~�JSx�Jh�=c%��ܯ�aSz^�g{�e�5������Hz��ϥ�O~:}�7|M�����a���H{հ��3�%��]�.��R!͖�9,&p}��:��fgws"�Ҟ�Ǒ��H�`m8J޾�B��sX��ʱ@A70�b����Dvj�Z����a�-��wC$��\�rm����1�	�8FZq ��^t	����T?
����?���~B�wv�~���8ip�[�H���8q(htU$�2��}�Z�n��v#(��"Ev��v��P����C ��DQ�������0A�; �$=s��$�uW @�6,�؂�3EϢ��rc����^��1��L��rj�r/&>��w��ϬL���AH����$C�0����c�do� ��Z5Մ��Ɍ
JUx�c�6�� ���@P��F�}��0�ò�uS���!b  DYU�dν���`#B�l�g� %g��T��|UP�خWc�]hQ���d���ۊX�E�b�6���w8Xq��ae���E,����2��L!Ć�'Bd�x�0hy���Q<S{fs�У��`�w 
~2�J�Y`@ ��I�7X&lN8��"��r�ޡ8��f��ɫ����3�A�k2Us�S�����}���� ]�@��F���흡��`5�2��a���\���w9����L����o���BXqe���>�5+�k�I816����>�9��:Y{�y�"���|.�-�N�S�ĥt����g��;�D�f��?���o������f␒��*G/ϜK��b���F�[�'�֮\H�c{t�z��.�a��"k��(�bW���W%z�yh�vTF*_�b-P@��ŏ<�dh J�	*'��v�*Ȉ����ݰ׫v����Z Y8��)_c	�q\,v��+����q|���� T��w�����[hГi3(oiX�F�����p}�(�F�`��:)8�\Z�EH�+�O�Km�N�#3X(�ƚ[.�7�X2L �K�$9/@����r�1�i���p9��a�pX��ݱh�� ��w���"��n ���g���}1_BZ%
*������b_Z�-��:��C�N���T@�V�?�F�v6�Af��5�}p�v�w9ę���T�-�����z����P������s��c��k�=�dܶ�4���O�;�!y��kO�ϟ�kf^��:6a�<g�O֥�����G����,����JDϥ~O�c���}سhIr���PT1�c]��d���|��+��L���W���b�}����^��m���@�ȿ�� �s�H" D��</�^�r9P��cG��)�R�'��&�k�Јjw��r����<���ȁ��?�G�?���N3ϥ��qO�'�׿M�<���J��a��?�W�w}�itl ��?�'����ӿ��O�ob'�y�0 쫠S���bp�h	�fr�Z#:{<vz��T������`{�(�D�t�~��ơ琉����k��ݹ�ﳳΟ�#m[���*��j��gX��
��� ��r�.�c�]���w����e;ӌt�l�VxD����P�:BN���v3�!>^��d���Ǜ�V�� �;��8qt2���؟�+ʎfTUfI��E����p�.������l����B}|6���x;�g&%t!�_ΔȎ#�K�4ؖ\K��f%8��#��]����jg�vME��]xv��:wY�G��+g���h�dp��(�;��2 �Ƥ�g�\�C���w��/�J�l�>��=gJ�����אs{j?���y��8��j��5@�F���z�����"���=,WU@�kʡ8�*Ӕ���ڀT�������̸0N��lg��}�5__�e{g`���������E;j�����Ξ�s��l���pc�?2��!�&������_�m|:�o��� e@���N
$I�S�V&m� g�ZS�U�`e�R���iY�g�sګ�?��%�ӟ�����1Z�<t�	�W�Fu�T���w�'��o<�Z�
wB�-��-��Ԑ�󘯊�Lj7�v��IL`�T^o't��J{vA<M�2��Ȉ��o2{�z:���Ũ}Qs���][��]�S9*��8F6���'��Ŕ��"w�vh!X��c�A�+07$�Uj{%.�h������o��̠�㤚v���q,.��G����ݮ#*\��z���i!��P��δ�W�q�bprd��{r�C���uBUZyδ���`�||��Z�ɋ5�t��l�v��N���%������w����PSe;Gb��[W����k	&��fdG�=��U�ZT�_;��E,�|F0*`G�q�]�3���<U�I�f���������Y>O�_��8�R�#! DnF�_�u4g28�X�@(_K���}�2@����S��X��A���b�2C����Ӟ�9ڵ�ϣ��lH-^yN_Ϩ������Ή9a�G���r+�/�|�0��$V���σY����v��k�6kg��!���:!d�M%.P��[k˅��s�=�z�^_�������g{C�������:�����ӿ�qi���&������'T}],r�v������Ks��JX=�������C��2�$��5����C5h�:)��Z�X*��<n�ύ俜�\��ֶ@A72~A�����9[&��*QB8a��^h�䅟�U%��`�'c&S�m`(�C;�l�Cw�M��~[do4�k�9��z��%RdQ��d&�_�bݍ�F��c#lT�Z10?�?�^~���o��2�,/n�}�rF�C3�"���]�v�R9;Z�M�?���I�Z��G�\��3���(h1(B٠��vod�j�Ɓ���z�B�%��0L�E��#L��:��x��y��k9~�w�\��Z&���Aq���ö{p�w2kD�̙j�Ai�σо=\z�p��<�# �����^�Η�v������D/�-�>\{�厪0bv��[(_��<��9���<��͈9H��k)��X��t���ܱ����g(�_���/^��l��L�#D������u�^ZZh.�Bׄ��Y�L?>ü�=��B�و��q���<����t2E����'5����T���ֈ��u\}����\��x3��{��
���q��3�m ���y��I�;����F6�j�#Y�Z�\1Zz.jt����>Uվ�������m��Tk�.��첢=-%V4	�S�[H������2�������FLY�U�jC6��Bz�����+�o@��c��m5\��I|�u�[��~t��ŤK����k�p��GJB� (ov���W�
����Â
�o�U�Z�^��B�Pe�x�Ks���f��n*�S�+;$��m�bU$�XY�I�]�r��S�ISo�MB	I�0� �Z J�8e�ә��
0�:��}����N�N�v�`n�L-�Ut<"�q= �@tnc�����Z�Wɤ�D��T �k�K�CF|Ζ>5ObQgA��C�s0]�fL��*������<q�0-v8h��69��w���|�<��� ��?�Ϻ��w�9�9W��1��2���l��=J�'�M��EA� f�c�(�r�^�P�'Ӎ+�˅�48���C��*�s�,�\1��%���Y���=�Q���{?�a��!� �U�r����~�#��Ρ�0�ưC��{f&�~)��s�a����i��$����ɽ����0!p^��z��g���x��hZT�΃�79y��ƢP�։f�yn���������-gp�pf�8e�9�Ky����P�'�J,\o7�ٶ�p��z6���*�]�-7I�Xi)�>��j��GL<���QC\���^HT8q�ѩ�óʜ��3�uakD�qT}�Ⱥ՚5��GBt�Ue�=�S�(����t�5�e뮫���O��ށ�jk���w8�O�(=���ɖS�j&��Y�[%$���+���n`�]�ǆ�k�����(�H�|�6�v��� '�ȖKl�5�E'�>߂c�,����V������E�`/��m;�H9��7�ќi��E�ؙ��,k�1�	zE�Z���@h���Z�����,�)�NV��q�
}��#b^Rh�3�H	A�.�3�T
�vyv�0/f�9pO�~P�BdS�ɺ��j�}�
��8�e ̡4X��D���9;��1�L�흮�ag�C��}�踕���5�Y�p8��r�j.U�7U���^P�Y��"2Aa�.�@s�Kۡb��r�9���a�k�s���qf�<�"�ʫ}��Gȶ���|��jKgǜ�'��u�T���sw���9��������'�S\��!�LŜsH���Ffo�D�&나��ޓ0D��������2�k�z�.��'<����&F�!�x|���U�W�Wf�4��a1��W����g��EMK��rTѮ�:�Cy|�����ꁹ'�Γ���S�и��y�WZ�.�p�4D���IG��sZhc9����t�-��w���H���w&z�҈��h[@gG5�:`�7�錊*>��K�"�]N�lߧ�iSi�0b�Cc�1h�S�=S�il�xz������ϦgN�u�X�޳���T5��̺��(���.�{k[���7a��QTl����Z֑uBժ�~j����WC�k�}9���p�_z��Uq��S��^G�{�� bfF��A�!����bC|H;��z@�j�T�e�"x��H�%����Uub�wC��)�hc�ʵ ����)��������q/tg!5��������n��Z��* H؂]7bk������>�� Qt���\s�F�q����O����-[��i9sث,"��q�륪a�Չl1��}~�C���4v.�K�&�F�0'��Y�g��cG�8�qW��A��r&`u|�o.֗{da�-�6�"/�@�C��p�赢�|�+��'�z����}�2�j���Ɏ�g�7 �����p�k���R�Y�� 6!�e*�ﶁc��
��T�����v=� GNq���s��0&��k 6�箻����64�７1�S\=��)�8߻Ǩ2fhŘ/h�\�gו��"�.������g�eXf)��.�s�{Ό_imx������	��4��>3Fn��zAhv�ldd�R����{��w��Kcb~'�G�g>�4��8��ݷ�P��B��?���@��;n��J�h�߫jLs����ڊ�"��-b����)qف�o=��<pO�V���z��ОT�<��*F�n��Q�^I��Q��L���җ;���ߺ( �Ʈ*W�nC���\U�#�A��pp��_�I�]���>�ŧ�3�_z������9�+رR?d@�b�z'Nx,RU:&��Ml��X�@�]g��=��Mqo8�\���a(m�o��֕��w�(`Ȃ�N�0:W��"o�&G�K΢��PW(�E�ir�ܢ!gj�� ��\�k�εJy�ޓC/�/U�%۸��iw�v�m8�ރ�u�����3��]!�������{J��3��H[ �H��z|e0�GȩЕ�Y��,Jf0��FA��dQy��sD��1��= $1��C|��P���7�q�dV�}����Ο2
��$�2�k	�G"�n����:v~&rh�lY�2�[b�۪ @�_>��� �
=y|�^�N�2�`;x��O���z-���1���ܔ׹6�s���2��#h�V�l�2l�5�����٬ |���Ҟe�{ܪ��̲I{)�6k62��*�)*�,H�M��N��4�d�	eq�x�c#B��U���J��������������[��c�	ZO����l����c�~���4�sZ�۫�Ѭ}+�J�P��m����|z����<�zǦҠjK�=��(�ZE*�RFj�;���@�'��r�7:�����( �F�O���B�YO�cY@�v'V�W��|j��������}�K'r�{a9pZ�:i�.�� �P�MgW�R,��e��*�2�X0�㇓��[A��{v�xQ�)�B�+�Ąi���=����1S�uX�Va�c5w�X�V�u=���g̰T:��H�����0��]����sv�����dX<�:���F��s1��5r��U����_�{�ﱑa��6���3 �nt�4j�1!R�:,���u��s��Y'�Ӳ3����mƞ{��'9��E�@In3(əKo��ɶk�d�o2X��Dv�y12ۘá\C�c���� +�7�<�.g����A�k-��p��e������&&��Ŗe]U~�x��_<_�����E¼)�]/b\�}3v�;�v��J���%�N���y�SE�����}��h����)���WM�c�!���Ǽ���y: Kd�*³k�K�Ra�(w�7~�7�G�|z��j�XYW�c�;x츲��B�W��W���z	JX}uz.]�zE��H����耲�.��J��M������SuX5�:h����u�ֺ�O#{���7�ڕ����5�u��|m��"ݽ�8�v��7:����R( �F�+�UZ7"��A��c�nn���r !^�lMv濙bQ�V��d���vГ�z�nU��k�Ϡ�pJ(�Cג��P��Q�:@HN��*���k��YK���ѫbuz�e������ ZZU�C�C���Ř�1@:O���l�
��b�?��_�)��4��(�2m0m�����g�9��V%
#U��2�$P
��@�1��l�G�uL^��W�OֺXoD(���haQ1��i;3��З��~\��v-�ru�.1f�S��,ZdD(��{[,֎��l��Q���؄��qrϙ!�N,��tݙ�����t0�E�K�������dp�>gہ��\{fX��8Ute9�
�GO� ���=5�9R1{yNy>W��^��*t8١�����C�]f��v͂��3�����e�����+vK.�Y]���sߖ��+���D'�1DCG������wD��vf�k6���=�f*��5�#z~�Ħ�V��M)7�}������V2Ӫt`���0o�UC��)���3�H���=��`�V���Yg�޿_��GF�����)ė���H���P���� i�N?��G��.���f.+D��^c{�hyM�ohCﶦ�w��M}���3�����z^���K+�*�^O/]M��t�����J/]�����*2��Z��9!;2;k�}9�[���� �aN�5���o�X�5��� ���,��_,�uA
>X�W�|�ICT��w���0܂�n�z�1gMƓ9�}u;yb�ľ"L[N=R��.�܎@Y,��.ޘEW^P;����N��.40hk���ڷ$h��`�6��4�ۢ��@߀T�uD���Jݷ�:fcv[nha�q�d�H�����Pz'*튮��#z����7Ů�zk3hԩ���0�*���Ԕ+W/,/�!���+]�#���]�Ȣ�` �	
p��]{$�CE��*�X�~��B��{tMjsВ&�~R��DcXgV��z��"�2��l�a�3�3�<]3��z�U���U�� Ե`�B�0A=�n����XON)�#����[ti���!1.ن���Fֱ�@����=NլW>6,��� K��m�����X�e��я�{U#&o:ܚª�pfܲ3Bbͭ`W*��ff�����!\�V�0=λ����j:�k�ޖ�\�Z'�K�]���*��#�HQ���W�&l2�l&�,�Ě<3���	P8BH�gW6Y�Ƃ�����a��h}⢄�jγQ	p�}^��YD٢�����CG<�n��k!�ݛ�{�Ζ�86���ٳiAa*lb��6��N�s�Z�� ���OC��;�Ÿ���~!}�?(1�������[Jm_]ZI'�I��#��4���"-@�o�^�G�.S)�kLU�WӲR�;d�~��U�&�t�N��.i�&�>m+����t�i�؉4<�H=�;;�Щ%�m���j��64M_�������߿( ��F��j�"�ˡ����*ڛ�k�D�|i
����.9Ț/yw�����ô!~�.f�PJ�-�C�Y^"f �FD@�B���om���ڵ#���{Mяǎ6j�X�]�`bWkڞ���-C#ғ�G��r�ⅴ�^Qd���S;�ɀ(�y1%_�o�T��*�d�Z�oto�>�y׍#��[�NO_M�OO�Kt��f@,���
5�A��W��i7U9\�!�ٱ�rQ�и����-̾H�	p��.���dG����U�0��"k9�ʑr<7��f�SV�O��S�Ք�&FN�ά���Q��?YKE=ܜ=Vμ7?~\;�%i9f� az{w,v��7�������-s0��x�Y����"kX+^�|��)��}�Cfb�#�fM������;�
��53K��c��RT��[i��l���0�1cn�&��܎ۣ��}��F�sW ؙ��]0���A6+A��˕7��g�:\�bZ�d{J���o��oN��}�e* ��S�BsY�o����#���du;�������PGJ�%}sm�w����!B���g>�~��~L�X�;��-�++���]bnв� ��U]��ŋ�
�t�]w�!�η��ѣJ�2�h�+0pb̯^�I�
���t�7Ž���I �/�=[N��,�7{媎����oJLx�*fh+�6WӰ�*����Ӓ�ua^=��6Ԭ�G��Rw��N%�KȤ^���j��_�( �6H�G�	�uo�3��W��p$�<�ηS�E���T�8�����رq�0"��8j�IU�Tv����~��ZY�0�k4y�1�D�����p�Nd@�ܢ#}d�D��Z:�w��}�{M�gMC79��>���*�߶��u�Z7�f"B[����2 bAǙ�����Kit��n��Q�`Ɉ!,{�`��c��m�h��-����XiQ�r�]���p�r0R�11]��zk��?�i���Ύˎ�� Ӗ�qe9V�l+����`��М����9��q����}�;#�l��r�^�Wr�^9J�J���6�`�^�ۀ�'6�T`C�0&�	.���������w}�w�f.Qp3�$���x��y�����[;k?,Snw���7O��7�?���@����-k�r�0�١!�6�fi&�o`H����|�ؘ�ߎ�̡!9���]�zw�_��#�ߛ�������Ӯ+�&��0<W��|N�@a�{��y�	��ʛ��}��;p�������7]����d�Ǌ���/\�ܿ�[��Z�%^�银"@G6�#�<bM�7~�7��h���F��6Ŷ��ы�@E�]�1�7���@����<��X_z������ϷZu�s�lR�gGzƁt�������l35S���k�4���}�0S&Zss���#�z-���
����Ro,lD���� ������]`!p2���%��xs�+ǥE��ͺ(m�U^��3�P�:����'ӷc��p���Jt�'�� �����Q�P�����*������_U;��x�0A�D��13@q���bސCw:���[�
{ 3+� 9N��`�^N��|_z���ipX;X����	�  D���3�K�Twg�!��,�`uwm���[������p����O��?V��;����Ä�e��9),�x3*�ŎW;`6��a����lH�2��-�}��O���O|"=��fw4��w!ʪ��+S@�-�P���z5���$�sc�X�C7,&l���[^I�|�C��sߟ��m�e�t�^�K�.�^���Ei���xv�j�|�v�L�g*>*��� �(4CX	���ރӥ�p���59�V��|��Z����`�ٜ���PS�I��n���tp~�#j��mzF��[��*�6(M�$W� d�E��^���t |]\T���(�������.\Z�3����y �����?K��P�z����=�q���}�������[f��U�bC�u���[�w�T:~􀚪Ω% L:����sS�;b�-���v�jg�3@���
�i�6]��i��1b�R�C����s�!����O�m���"	z��"L�X��?)���Fmg���e�&( ���sx,ZZxs�=m�<���X�_ ���_Z���𲣮��)�8s.�~o�A�'4 $x�i1����t�}�Iԧ�⊳�ܺ0����u�2*}�'\�g�ӒRsYH��k�&}��|�ŨgN��uf�s��ώawW�P��a��w��E�ŕ��
[9�xo��ᵤ]h��[T}��j��#_��`P�KQ�:��[�ȶ𢻦ٮ��@C{K
��`����w����ZD�otIPuݙ��3ϺFM�N��0 ˵e�c���,h��xe�;��4r
�y���4�GB6�����O�9��^�v(���뤩˞.Pɼ�ޭ�i>l���}�]�/�~&��9�g
�����Р+L3';|�?���	q'+mJ�-� �}���+S���#�vɀ"_weF��Ie4gR����	��^I�o��t����ҬCG�����R9�����ML���8o���f�w�����;q�Ҵ�9c��c_L���Z��=����^ �J���m��	�X�j'Qu�LP�Q���V:
�nT�G ���s��F� A�U6��r������~��ނi�c<K04 �?�?��t�w�Y��B^u�J��K���+.����w>��i�Q������1�����Κ[[k�q!�F����W�]��ӽ�ݫPۢBi���Z¨�ز:�SChyI�[5^�R��rZi����v���ꍸ����i�ʹ��`G������6�@A70��o��;^���ڳ���k�������@�|c�^��^��W��y�� afK���%6[a��dĳ�8(T�D#�LiC�9���#��8d' "L��P�3�d}rT�m8kI.i���l��_x����w�ig�vf�lvh��?v���v��b{��bQw�����By�f��[o�9����w���?��:s�t��N=�}=�B���4��Q23���W�A.��5y�����,�n}���Jw�f�SO=���������-�����x�w�a7�Q�{"ٌ�Bt|m9D�ٛMi �4+�O'�˯�z����OX��cv���-G�� �f���B�U"V�-ɺ9A�+��)\�:�^�������ΨH�%�|~����������wλ�T�F���v�0f�=Ö��"ff�~ה�h�Wd]99A�0ٺ"�b�������x���?o��o����!�=}���������ܸ&���A�������Y���Z���a�?�����J����t��)����+�����HO�8��`�t� �&�@�wg<JϷ�Y/�\�~��Y�K�B!����N�^�2x�Գ�6�����Q����|������~o���|�����=�d��u�h�Lv�6<���(�}4�TK�Ad��]��Z�أM���\�j@!+͛˗.Z�`FC����-��r\ӈ ك>�гt��	����t{��J��Wl���}�/}ʎ�@�0�G������� Ͳ��?�cwUu�ӓs��f�����` Ex�
�$�$A	��������a209�ι�+����}v�3=��L��?�z�����>��{ιg����{7��L޲�o�6z�����p�?���ge����A����w�r�P�Ŗ]��r�{sq5��X�@po� ��c�GcPŤ��®ҡ� e�Z�>�b�2`������V���92@ۖ�\c���gE��ػ��U��H.�}j1���pQPv�ZV�n�x��y������c��򒗾�|�/?PN:�$-��eb�ds�w� �����iP���Ge��
������Զ�2�~q˽���QI���>o)�׭.�~��ʕ߻���������m`0��7>���?���n)��0�O�� �ņ��н��/�+amy�{��0����1~ի^��o�fRk�L���njdD�8����$�7�f_�%C��Epޣ�>�;�O|��C�Pٹ{Yѷ�<��*O�姗/}�?�"Qe�"jǟQ�Z�+�i�Z�iD���dL9b   �)�	l#��)a�Qrý�o����7��|�ӟ.�wn� �����Cҙ(�7ŵ<���܌$Өsdcj�`	�yWb�v2�;���c��s�5ה���_�˯�ܺ��=����xy9�Q甯~��:z���M���;٧|~���9_y����F��������]��� ���\nP����9��{��_'v�!EG�	L7`��)�x���"WW ����ϻ�ȕ�AkƆ�,R���}�|�ӟ�u��Fz�ﾠ<��Ow�����7�7e�r�0��D���Sc���zѧl�\�c����G<L����>�պ<~�[�^�֐pѹ�46���ͼ�����K����� �� }`|o���r�-7�1=�]j����A1��{U�LݲO����eU��H���vn)�z:Z��̝�7�y��̎�_�;�7�{�䁡Ѯ�ˇ%؞�Q�f�=oko�
��sV?3�9G�-]:%	�)X斞1�0���w���90H)L/k��ŶM�)E�Y�ҠiV��g�:N�d�8��uP�]_V	��	}�ލ��ض���.����ꁀk����	�%s^�{��u�гkqqH��N��Hj��EhQ�"����"�� -�]��yR���{`��q:Hn��kWy�w�o�;^�6n����@�>�z�a�)����_�0u@�1Io{��yQ��<X�_��xg�n�7�,߁�O��l���^w�,�\�벀��q���AC��7)eㆍ�������(�Ʋa���w���q�Y忾�������Y�%�'��,0g��yِ�����aCW't��܉��-�|�3��@ h��QY]^����a�;��������]u�gZ3sZ��l`�6퓼��5���6�ȵw���iW�x���'?Y>�5 Z�r���}�s�)g�,W�x����]�I�s�2����R�8#\�b�9���k�d�E5~fA�
�x?�)O)'�|�������s����r������=w�`՗�a#R��1�Q� ����O�>i��G�t�l�pls����B��G?Z����ҫ�9��򲗽��Y��ܦ�y��u��J��2A���P S&l���.��VKP�X�:>�3=�.��2��8���EP���-��|}���?���=��e��NLC�O�A��M�^}f�(�`�������:���7K/����/��^�yĜ����ny�����#�K.SD뀑��<9�)���a0u��H,{�'�sĦ-t���Z�tTEs�ca�����j^S,��DX%�L�����i��l����,��T��2�	X�j�-+�^zi�v���7/����S��KK˃�z�X�����o,]-�=m������ۚ������ͱ��M�M*tR"r��5���ԾwF�ш��P��wN F�;��թZcg�'iV��h�פ���r�c6����bKZ)4;�ci�d*��tV�lLl�>�ߴ����;{P}�P���5�����/}�.��9m�O=�ԫ�>�+�CM�O�� �0F|^c��P��{���;�{[$�������TM{��6<F_#�K�Az�F�(!��wP�n6��,�?�9q}.=��d}�Q�%�d�|��֮�B�{���Pn��E�*���b�0�0�$��A���ǜ��^_��W� |�_2��7������/g�u��$cs��+|<�m���*�n���
��ݥ@VÈ��}�{o�R%���N?�m8]�������=H�y�\ ��B�Y�@Ȼw� b�Ƅ�h��~���XM�U�N�K��q���x/��r�]���w�׼��e���2�������=�l:rS��5�h�骰��1}���_C����#�������� ����rĚM�w����W�W�9��[�̦��B���d���_A(�EEe���qM\n��	�(��E��42Z�bæ��S$�P�z��c�)���3�]��������UX�𕯲�Ρ����sA�O2��u��'P������%[c'훘+�͜���`�MoWoy����x�+���!O���;�0� etW^�=�9��w��R䍉�B����R��Ѳ}�v��?��﷼�-n��뿖e�׫4Ĕ��p	�O�*�n�p�gA�y�Щ�c�o4\qfv�ϸ����>H��s�����?��.�eT��]��qDs�R%���r���[��5��h�y% �V���4����l����vq$t$�����:�`��� �y��Kӽ��%���=9W�"͇k������H9B�չ�>�\s�5嚫�����	
��9X�%�����꯾�%e�e�ms��g'$�l���kmk�`M�RL�S�}�\��w��v��ܬƱ�t ���Ҝ�̜�g3��3���xN�����]�6s:fN� �&m���� ~��zf6�75����Nj=��'=��#6m�������}����_���0��O�WA�����4�zḿ������{�EŬp�n�mz���U�'��~�py�cD�G!�3J�7I�0��X8-R�y��6Q6��߹u[��p�)'I��;|��K��c��I�T ̤�\nZ�"��6U�W~ �R�u�7:��Moz�싾s�������򗿼l�$���3wև��7�\�<9ћ�w�t/,��;L�������_e@.��2kN8����w���r�)�[n1xs^��%8d�%�^�}#�<������#�wja�'랓j�;��)*m� F��IO~�ټ?}�[zv���ۿ+W_}MY�c��$C��z��  z/rN�d�</ݤЁ`����X�p��6Q^�◖���۠n��b`y����o�9���.J
�6�~�H�9	�i/��ߓl�e�&��dKg�FRu  !*�2�j0D�/zы��A�>=��o~.�k�xq>�~>�^.�&��ZTXs Dx6�,=n(��M7��{�� u��@�s�����?ݶZ�x�]�����Q_�:"��$ &z$\���G���Qn��A.B���.�`�φ�we��|�Ϲ01�_jX��g{k�2�9�b������?�s��t3[��J�2(`@j~�8�21;�l�]J�1w���r����+���kָ3��v�~�DKp3N��]e�`�p�"�_��֖Ve��͑
�Dݢ����u��?��;-&�r�U�/�vl-S�=*��?���x�1eǖ������\d��Hͷ��+��ڿoN�[D�4�uv��u�x_��5I{47�bE3A�<��rF��Ts*�ɵk����Ӥ��\��m�C}l��S�6# #��J7��A���o��U���9�E!��a}4�N=����O>�G�����M��}[�]uǌ�ϯEt���b��$R�i���@X�{|)��=�?tq�/&�����y��ު���3㢡��"��t�@����9+��E�J���&"�N��f��M�s�N�u4����B��%���+F�W�1;��2��A��-R�<8(��}v�K����b`q��U�Vڨ:^�җ�=����n���VLǰ��a�%uR��
��I��2(S�!l&[�������Z�I�v�j����K��h7.B،FÖ�+�q��V�)�b�������q)��(�1�hX��*_ Ӥ�\y��~����������f�?.P������UF�j(3p����M�V8���r�/�vW ~"j�E��v�1�KUy�촓N���V~�)?�]+n8�"���v��A��L���E�6��(q��\��]��=�E��Ι�X� �8յ�y����c0 ��8|p��)T�&���|�����=��]�Q�t��oZ��
�ݤ�C�D� �I��a���]�l��K�� �
���ҿ}�u� �,�Ò��}Fs�%�����W��k�q^��g>�:\��I~�(l).j�W!�i@��"e$N����=�صx�:�X��|�7��ՏU~ƅg�1Kw�-��O�y>��~����3�>\+F��c�ZX��o��\|��z�������[>���T����v���� �Ѯ'] �_����_�)%q"����g��eҰ��,k�u�c�*M��u��zB�����ȁ��n.����̌�<�]��jͪ=�㝽KF���)Bv���D����.���葇wfF �S@��j.��y����O��aN�O����j�Ӧ�jQ?�h l���6������S��K��i�jW�~�7B���u-�7u�c{����ƢYk���'�x�>�G�C>_A����Ԣb'��HZ���V�k�w��K;쵨�'l�yy�3�d�}�B_Y,��1��,..@FwZ6e!�H�ء�|� ���916�ZX���.�k���Yvn�M#����2
{��uJ�=H��=��`�5F�6�rqӈ_��|���[�������W;] z�$�|�+^)V���;���ZL34=��Gu�%=J�z�;^���Y��$��P2�#T=�"�9]E{���4>��L��駞Vv��N�pT�۬E���Q��ɇD?�ֱ��q�ӎ(��;Z�,�d���C��:��(Na�P�N )��s����/~�\w�JMp��ĥm�;�6� ���5+�8�>B�N�U�)�Q�"/�� y��Uv/<��s˳�9��7+�x�4'\����-ޠ��2D���u�"MIv��ġԎ
�t���pM�t���U9dd�	E9�.�j"�RL��0�-�H2��n�Zz�'sSOh�`	8/._�`�hDJ2/ �f�@̙�#�U>W�'�Ͽ͞�?\�������D�x�1��nW����=
�)U�9�Gf̘/5h 3fG�e \���ah�������@߀;���/������1�^_�� �+�J�ad��H��G�gua����U
@���ث�ӹ}t�۴� W��MG��Qcܛ&j�m�_yy�=�q���//;u7����/~�<���v����F$�)�x��6�M_̨� �{Cr[�M*��k_��ǋ��㞻�a[���w�܄�Q���t��^m�Vo(�.�:x�ƳM9�V�9;E9��^��ѳN:�?����(|�U?���" ����M݊xY�U�����?Z4O��m�{V{}$j\��q�G�9�$�����uz_O�^b�[�<�]�ڪ睷c�B��	��t����3N?}��������v���zFv���s&�� �0�}fl�yv�%U�>G�y!0v�'�C2<
cB�{�X�Bg�lR��o��g���qP"1��5! D(�X�v��e}�on�
	���U�hQY"��Gn�v�
�2d����d�D?��*C{����yO��3	�z�����S�l]���b�^E	�
�/���N퐹=���TbqB�D�!S�j+�vьLkGv���)c�F`��J�j	i�c�B���U��->�]e^�CTvC���
mN R�����R���qF�x5F�y���	'�\�ؼ���k"��KYF({��([�f٣�b�����Nډ
Q���ݸ�?�o�S?Kd;.W���$�,�BH)0�62:]� �}h��N\��1�2!��\;� �qjfL�$ˮR���Q_H��p�EA��aZLaP���M��'�~X7��Ssc��fRV�=�ɣ��!�9� ���9�&�H�<e@?�L�o:e������H��µ���� w��g&L}�.��ф-"c8O��;�z,���h��sB�"�:�(1f�`1e�f��Ä[sR��V !Q6�9v�Sa�sN��P����=�r�F�۸360"f��'�`:��J���� �=K��$������4�:":;4�y�?�9�[ fV����/�^��%�sP��nX�	���+��,�˗��;f���@��Hխ�b�zB��2���˩��#�]�����Ĥ�}l�tܚ�G���{��}s��f���G>�a�B��G�{���|ƕ�׷�I0���$�mry��R�h�	x�J��lE�~Vλ 1@ο"�?�&��n��N����bug=r��X[��i�*]☞�Y1���G��L��ڴ�����O>�������=��7��b��������)?^-YA�1^^2XP�����Q�ÀN��W�1L��s��/��4�\�ݻA=�*��퇗`J[��(p�\Om66M��o,���&Y�� !�J��z��`D�$�!�2�C^����.�X����)�9���_��UO��ya� ��;��^v�S C-� @�!@�����F[ �@��	T�TT�����DG��3U -�a#�r�ɲ���� T��-�U9zB��1�b� ��w �����e7
cD?��r]-X�H*�:�_Z��ႁ^p�jk���伄�ʘ�=hH��ف�� ��9�)�׮8�(J+A�����
v����+�������zFet8*�WfmWh�  D�*��E�� �)��U��#�{D(2��
�{ڗ����uyk0b�Y�䅋C��G;�1Ր��k� ��<�Y/�$�!�7��Wj�RK�|������Wf��]�ʢ�p/�V�x�`�`���5�HVI?��D*��j��!��z1�R�!��}	ۅp F4}����   IDAT��ȵ�fdTc�ry��^�Fw75��;�^|��fLp]Პ���؈�pw	�;j�6=[`3@��*��ȥuwII0{�x� �������oܚ�����C�neEV�!s2Q�R��{��r�uוg��3�G�9c]���[F�}���z��o�V�'��6�<��1�	�A_f c��g���z�-��OQ��Xtm*�ڶL�H��jF�R��n��!�<5*���1a���i�Etx#�U��^��=T�G]懂 ���R[��yJ������E�l��ܦj�]~�wV�)���#6�n-ڰB M)9�0�x*fԙ��EӋ��<��lU4ǔ.�#�٥Wy7n� � ?���v���Z���(E�C��%,~x3Aj'T>fT�����1�H��X�7���N�|LA�����Ź2C�d� �%͈@�%b���n��ϫ>�4��
X��31��}UgЇ;���9S�l`-�/t1$�P�bIg�Mqo� '/ra��]a\&e�ڕ�������(s�.��.�5��V��)��T���R�R�i4[�5�Co�9nڴ��OZ�� ]�I`ڄqI��1��:��=�r�`g�y7*��W5����$�Б��"q��N@���L����H6��*�M�V���H<����R�c�oW�����3��W��6e"C� �k 3�U~��7��|j��<Q(4�5;v&x��^��C&f�I\p��H�5�H�hw����(N+�c ٤��+M���:�MJ��1��pa�6�9?�q����%֣9��(5��`���q� (�sb�`�j�i�	��}=����c�z%�~X�� t@-�l��w��]J�U�n��W�������t��+N@�7�c0��'c\����>mtT�L�$���TG��A����kS�T=�btG���J�g����e��yj�Ij���OM,���j-bɵ�xY�
�K��E�*@��,�;w3���šY�F�A�;QS��y~AeaܿOy~n+�u�(�E��P�w�X�(P�!dmv��2;�V�,U�V���O>E.�=1E���hTK
Cc�g �A���Ls�?�7���QUH!$!�Љs��
c���*C�>��]O(|��a� ��!w��\*A��E�AuX��̈́l+���#�#��� h��4t&n[�l/ ��$zYl�(t<�Fz������b��B�;�\�Ղ�̑7	%V����>�63ЙUԞ .
>�0��;-s�p-'�������꓈`���j�"��7s�[�#�����p��]�� 5��	7i?�����\�Quj+F��r�F��5�| /�4��0KT�Q������)�Me0��Y.����l���{����@��!��Z[p;�!#^�e�
j�>cd�Q ��WtM�7�3_�$��"b�dY�|f�L9��g��.�M8�s3�d�Ft� HZG�;ˀ8����O!h��2ĳ��sTm�L]�w��q)~��D��h����?�Dg¨�Zֿ������� �c��.f�6>KNe,Cbg�����Tʊ6��ڷ3j���S�	��d�O!�׵a�xx8��vɅ78>��\*�*h�
$�+^�_�u�-R�6&�Z��:���e\l�"tv������q�����kA��f�\��esa?�74.��vM,SdC��creQ��u�Xt`г���c��8+�* 
�NMg["��O��R�^��[�k�+�߫Eh���Ұ��=h�u�9稀��f�>��ăJ�ȇ��A~�[:'׶�cgk�1-h�0��@�C$D\��B�6j]�����6���X ���@]�C@�I�&��aq��Q�X8�}b����:�� ���rn��	�<�\) *
�E�)�^�kdHh;fG���j�7Y��?�`?3�*�dd��R`P7b ��\]]h��>��U�dUG�2uR<��G�*v�$���4�e `#��耘r�2�H�QD�ъ�Bn>�3�A�̆���`4��0�#� ����s�|_�W @����>G5�97z1oH�0����{�KLFS-����V&��x�f�)���B�X��G�D<�9�ZN�5���=��,�|F�6�XW,ܶw������y�{N��?�Y�{P��������w ��abn;5�cF�����dA�J��/D��f���{����u�y��p]���B�+��&r��e��AT�;����R��]�g�7�j�w:ˠt�����:�+q���zmJ_"
�+w�A�?T����D�Vvw�9�GA�)#���K����+�vPE�>|%gT��4qm��p�)��@��Y���1���>��䨀��T!¬a�5�t��C�էr����&�Ώ�Ո>��\�~����%�5��X��֯3� �T��������o{AA����'ѲY9Q���^(fT�͊�K%]eր�c�*�B��pW~1�e����W
���CJDYͫ�r,�a�c���M�UBs#���Y��f��h	��]Vƙ"�0S,�Q:� ��6�8\�"�òTwE�؏�&7�Nh 2���F��;�9��DD�XlЂ5�}(�/�~`b��Uf��>c��3|u��ZO,�5���n��*��
`��]:O�Y�	��F�[&C�.2��0H����E5��w�h"b'Jm��2iWe� ��qz9��3ˊ��cB�	��,�;�GbS׃�Ǻ�`�t~�R0K�S��߰-�:�T�h���b^h� ��Ɣ�w����s�έ��;�,Y�����TjT��L��k�z1@����{�,�k��u�P���4T�/A�YT���Wd��te?�3yz�h9j�6� F�8���|�M��S��A �% �ov��� I��c����Iͅ~�����0��d�&!��ilzڴ9SZU�P��߿ҥY~��^~�!g�~����ʐ���t������3XfO<�w�QX XZ+'�p�O�jo&ꆫ]s�����<�S%�n-��8P�$����UR�A�16V^+�v�6�U$E-Tg�⯟�Xd�k��(�4�^D2�p����#ռ&�����s����RP9�p��h2�щlB����p��Y��Q�'D����17& �b�M����hvh��ѰvSc��Y��.����0#����d��n�ܒÆ���;�&+D�c�Xܜ,��A�~���H_�F��04�F��"�J���X��ŁB4	�#r	��H!]�*@Ӏ>B��Z7��ɴXڸUMNFq��#D@�T�
#�9Bۓ!��Vm�����̔tOji mD�0�� Ȇڠ��6�\+�0����`E¥6_c*��0q��<��"�3�^1��O�������Tc0�G��864-�� �/ے�@#�A�����s��xL9�3����>�le�~Fy�C����U?i������T̃|��$t?��C���@�ܟ�j�`��B�7 �v��X���>��H�s��{v� ��EϺc����-:3��x�8�ɂ�
��8s-���v�����Z� �lW^��R���&fs�Ϗ�Ž��e�ÏY<~��&�<�w��9�!�ϱ������:�(��1��h��hk���+�?#GV@�k�G�o"��3?�ĉk��g��qY'�ED�w�����Qf�E����ٷ�������;���u�l��)�o�6_o|���:q���8yS��tp�6 ��LoZ�|�e�����L�a��x=�aXb������8w~���Q�>3���nl�1%�z>�By0��ڧ���V%�ӂG">rgP_jRB�Equi7�����o��"0�]��(�� Ǯ�X6(�F�v\�Z�o��z�v{gժ����B��?FA�\_�x+��	�ɢ�D͠q��i��+� �=.*�S�W�V��G"�(��ϵ1 DFQ*��M�@;<B��u>tA��tYv�Zxq1�y?.���ʈ�CV[:I #J�ȱ����R�&������ �Q��������Y���dd�]�lPB|�g�Sʝ_ù)�}3�>�������B�թ���i�7Qpɮ.�M0.�����W��>�AAה��]�����zֳ~����,b\��w��u���!ȍ��z��8��O��&��n�lG��1C7S7<��TG��P`w�\qI�-0I��}�߸�E8`ڭӍ�g����� �pfu.�gw\F<��������آ�0���>������3�{0u@�����y���n��'� �����%��Ч�b�f����V�*.aAz94��/��Y�k��~�Ck�9�O�������2�3W����H-3_�a�Q�eY���UB�%��-�il��6��P��1m@
֗���kZ��r��c{H!m�Q��� s[�lw�@g�"�(����\�a�"Y�@�M;��9]D�G���6"5FԮc�0W��4��^b���|���{`��k`Nq����@���b�F(F.�C_���[s�t��V"�&_�Bx�|�$��M��ain��cnZ��2	͠ȅ�G���ŤO��֞�t�r�vlDfj��L���)�� �����=u�[P�t�M.�� �*��;��f�%��,S�� 
��_��`���C��CaF-zYu>Y��1��`\P�D��ygN�&Ј����Ε���{\gXf�}14�:�$?���'hS�IjuyY3#k��P-R�a>�)�A�[<Z��v*�Q�� �\��ţ��0�f}%&�ς��"�P���ݔx��i#��(n�d�<O�6܀�­���|r�Ufʺ��J�=/>�9��tuw���v)�����#�OI1o���S`d�4B{��ا�s�
��
Q
�΃ԃ
�-yoЏ1ga��p.ړ�&YϜ����VkV���=�7P{0R2�
6�l���n* �Ne!87mc|<_*���������]&���\6 0}�{0Fzܰ�A�����}Ŀ*�K�i������K<O�����[���Rq����sM�z~��YtA�o4a�Hh��F�繃:G�;< �ni�@�P$U�zFѤ������y�7��DGح�oʬ0����QE�H�P��ܪ5���*��D�_�jj"�Q��ŵVe5V(G���Q��K\>*P�u�H:ʆ�/��/����7�+[��i��%߽����o�{Ri֯�:�M�XO��i��W�C����*�a�ܤ�aQ}v�����1- A�e�� -��� �v~7��hr�]j��3z�[Z���%!����Eƿ�#L2)� �uƴS�P��
hav��ܖk1�x�á��	�C+��P�
�w�$�h+��VX�a+X�X �QHS��I��|x�f �Sp D�2�J�n ���)��^�2�.����<�!F��;zYӣv��.ڋ� ��v�2�b}l�|�X��F�9ޠe�����6���S���8C��vH/T�C�R���'��5�@�u2:!���]dc�v��v#�R����W��V@�q�0�w=2�����K�M5p�u,�Uw	}�c<N:�de�]Qv��D����]|��v?Ў�ڑu�	�� c0y�P3�O�bi�Z����4� ��(���/�G��e��p�Et!�������-���i�) �{>T&	pD3}ܾvӆ��� ���{jk��h,�1�m�S���(8�+��s��]������'�#}���XF�`P�%�\�VnB�c\��0��i��&ɜ���(L�$S(�n����9ah}F)�C9�K�tTnz��s�A\�����q�K���,]��c��1\��F�"��S��q�>p����׿Z�UY��N;�l���T��%�sܹ���i��^�U���O���L�a�q�5��� E9��ٛr�vd��§�"3k,����-������x7It�Q*�w��%&C;+�o&�9a0��D5ô`Hud��9�X�z%T�i/w���we��~ة�q����)@C��Ek�Q�0 �s$���8"Q5��Е�!A!��@N��j�$����ذ�"^�%�r�Ο���~5�DSm�"���5��zA��1pVae�G'��)�$?�#�H��@*�^�:� ���Hq��pof�zlӳ�Ny�r�]��iGc���d�0Zb�� ��
�ŘQ��A�<'l�j�=���l�LP9'����f9S��	��5D�q"b�\;M�י�f����nL�<"�&�t�:A���fX�2�Y�9�h�6B�q�!$W��.H���V�l�����0ٖԝ��rm.�O�ie��N@)Z�Y�ҍ�&���!A��鈢�3�A�L-�j�+H�K ��� s�9�9�kOc��G��(?�ju'1ޞ�l"
�MTٚ�g��-D��Cn
��� �|��7� ��,��q����.���l^���*�F��1�ٲl�
�A�td���SD��t0��g�Dmt�I��XJ1�&���k#�W�r�맽m�#M��`&���k��}��R^��=_p�M�h}p��&r�0�~���%�������YH��]�J����ig�����+����v�ª�h^ZK��pZ�V�H���a؊ů���E&�0�F��)[f�O�燩i�y�#�8~��3��E�B-����4�;X��y�aт]�8Y��!�E�L�^%�;���S�-��z=y����%�G�U%|J(�(�)e�V��q��9-�,�$-���c�,7�~��ګ쪚�a��Mq���ʡ3*�t��˪�8����C����ۨ[c�����;..m�\���~�G$� ��(2@��( j`��(į�J�\2M�H�@6�ӂG��nh4?`Q��2��ԧt #�UvY�!M�DٷG�?���M(d<ht��"�,�unZ蝹�z�wg�� �@�v�wы �e7�O���@?�B;y�t�l�1�'��L�5\�������%�:ҏQ�+`-�#�*s�DԺ�i�S�ש����<4c���n[�'��v�C6t��k\3�i�	�+D��oGQ�ڙ�M=*�:)f���9�+�U� cءy1�Q�n��Ʋ�e�-�b]��"�0���,�Mt8bdGj&��Y��"�
(Q���p�.�9���'�v
�G���sűT6Oc�k ��ѩ�J[�9�v��<L@�����^�Q���%U*kn)��`��fʣ*Κ��'z�ρ3��(g���]?N����O���eY�̺����$e|u�V��c���p2ʇ�Ϙ���B�iPX��SJUt)��ʜ�ɉ,%$G�?���hS[ft!^̥p�(#���J��C��5Qɞ�1�?�3{����h���m�:u`�6�"����J��m��l��2��5��'@:�cg4���!��Y [[7ͭ����|�\u�b�����_�6cZ;�` (km��_��Y����"tCV��E@���?�U0UmKLK��;6N��#_�C�r�U?P�5���~�g	mfW�,�+���G�0���"����
p�����Z '�e�t��n�#�Ԃr��7�uJ*�y�rb˦ҹTQC��3��j���阘����K:X��]��!ؙ��c
�5Ô���Z$���J���~"�0Y�#�lZ����!J�~��+�r���iX߹��ۜ�xRmb�O
5�+���:"a0�>oU��
��a�yj-MK/��|���$Qi�y8F��mD-���o��5�G4�!�˱*.�<�.�ta��m"W���2ڴ���:�0����M��sN"�y�R��GT�D��n���@�N���� V`킄�r�^���p�`�Cfw������b`���΃��o��C��}2�d�$ÈA�~����w�v���2�����$%�c�G:_��sϹA �	p�n�f樒.��� 0Y\���e����؍�)"qxչf�,�� T��b
R��V��0����"�>�aD]�T��}f� �75�-܄o������=�F`z(ܘ��� 70��bԩs�c��)� E����1"!b���#�$��fb�?'��6�a�**l�u~�tJ�]֯f�Y�X�)G�+�B��Y	��~��)(�"�̳�<��q����5�;�s�u�63\K��`�d��%�p�;E�zLl�n@{�Y?�_��j^Sό�%A��V#p`�D��s&n͉�Q����R?K�D����W6)O�*�ؤ��ގ �M��B�wsm���(h~%���c�	:�1�3#;y����W��`��Q�O���7z�ͺ ��]
A%[-�r���~�������}2R}�\Љs�9����ZDHH�S��]8:%Hm/va��٨v�-Zغ�1jo��Of'�5���c�pQ�R��	W
����h6�� �R!D4$�cwR��ZA��'�oF}
r]2��q�m�U�Ͳ蜔1��i�\d�-΄u��w�[��1�\����PV�n�͆���2l�!���C��mAj��e���F�s��`��ϺG�H�?`� u^q5���9��K�>Ǖ�¡�J̙�Kb��7��Z^vu9^Cc�t
_��YֿRI�-~��r���hǽB�O1FU�ù87�����Uv#���Q�*���^���hG�D�	�F����ŋc�$���7�ol��/�����4�8'ғq�ֲ�o��׫,�$�L�0hjeUw>�oS��: ��L�yO�$Μ?���炙+��6��q��w�¬ߕ�t�'��o��a���8�tK�� Y���f�D�	�����2�ų�3�s1�VZ�铑�9��r��Mб�]����7��-�ɑ�~�j����y�`N@��qk	lV��2�Z7XwAX��[��U�ݴ��a%�lW(�D�P�sb���P�VT�'��7a�gt�ܖ���ƤGnᙩQ�h�V��Ea�K?I�/2A�9��_����B{����c4�@?\��b�w��6��8��&����v�h2��[�c0<c#���|����q�������.D�*1�*��ev(�<�m2�=�ϙ*kǏDQ����NeO��!�Ɯ� ��ؑ�1�Ckbwn��(�Y:���	$�c�ć��!��.��n)D�S���`���Ϙ�b���kW{!&Q����H���е �Z�b`�I����ar���6�3vd��+i��7̂� $�7bC���V���^h�Bf#�P�0İY�*�>���@PlND�D��S<�� �=Mh������P�fڕ ���Q?��q=-�3FCͱ�/m4�P8� 6�2�YS��ͰX�O|�S2t�˙g��q�`]�F�Nن>���_���__��A�KD^��y�J`\���Y$.`ˏ50���lT�K�1O(����)F�c�`~������ �1�.�u�p�dɌ��m�=�����`3�#�ŋc�K	x������fD���/!��l�*��|��
�׮B=���	�b�G!Z�3�!��������f���g��V��
��=d~,�h�c��	�0����M�RIV�ڼY�;����;����kw,2'{%wW;ωj}�/W��и���ݽ{�ֺA1A�c	 զhQ���>fX���k��}7��Gsp\�3&'��5�m�f(`�����LA*!_��fz���ô�?N__A�1Zf��Ө��;��!��Y����.���d���`E0������� ||
q/>{��T�&tW �?�y��=Щ�1�z�c��\+K���zbRt��9LRE!����{q�`gE$E
���aXj9f^K%�D�aw@	V�
NG��&��Ν;j�
n�������85�k\<�d��AY*&��0`���P\���4BZ�%6(�@�f��U��f����axj���z�[�b\޳b�M�{�mF���B�@�����d����f�N��$YG8�C2���O�+������t.�U�Q���w7m:� j����O��Qd�>��m��r�^hI���Hc���b@с�������v�3��_?��5;ˉ'��H��va�����_P.���EJ��d�0� (���(ے��1��6�$�\x(sܦf`����F0����� ~�H���W���g]��B>�f;��2��(E�W�l�D�)�yN6���^�J���Pdr���X��8�0���SG��:^v[R)����xڗ��X��AU|��x��x���/�LF0�d��O�!^v���s3��֘O5����� ��iLp�nX��������v߶us$U���L�p�w�֛#�?AA�r�o���mykY&`�k�N�X>;wl0"g�)�	F����C!�Z/n���#�;�t��*�PE���M�UǬך��K;��ZF�g�^Z�ha�-����� �0F��@̻��U���pe��ra�nd�~D�LQ��ع�aU8�w�,��4f%6���tT�a��$N9�$�49d�����1-ڰA��Ds�o(�t�	acH�?�4�-�u�^M�E���������H{���E��5F7��Q���lD*����k���(^ ����Ȫ���8��r�"=n���؝�;�fi��C�Kc �DY�m:`W�V�?��0$�hX�A|�E`���l�F1� X�FM��-��LP����3:#��t�ѩn��=�
���a�aÅ[�蜚Lcc������ ��A�v$� ���[т�v����c���0IR��40�N���H;}w�2�M �����@����2 @s�1G� ���6�%������ng� �x�%�:�&��Am�~1������S�=.�v�İ�蚍N�h��g(�*�G�j��6�5����'��s5A(׶��n�p�;����`'��c��t���PS���<uT�"�)�Xe�d���A��s�l��Ǽ�儕�5�8��)� *���R�d��zew�څ�'A9}i$���c'X{�C�ļa$r^�Z�������T�cWy�~�ERٶL�5B�Ӷ��,��~q��ݿ�ŠI2J1f�W딈� ڷ�?����b��G�ZE1�Kz`\;˩*�A$�)�?�P�m��i��P�}p/Y#���5�G.i-Ǯ��9�w��������1�R2Z�p�I-��2�����I��6v��H�\�x�d����3���f�hڑ:�X˔4+��yZk=h���mo�)�16�JTeG�-�Z|=�XA���=1*]����c�z/��K�g irw�;��|jw;�C��T��z$VHB(��+�biƴ�_����vl���A��أůM�m]F�A�G���"�:�g��:�����xr�6(X�K
v��� *��`!"�pDu��TE�1^,���p��0�G�t-\$��A���f��CFXt���p������]e��E6��G�#����/Ԧ"��s�P�^�:$'~� ���b`�:)��7	���"�j"�`b)��u�L��1�zd�%��#<�e#Su?K����n0|��.�6}�����~w�fԚ�k$�^m��F&�>1��lOʴ��O����=.�V��ރU=�#�M��NY�!�0"��D�B��;!󸬔jA�s���P;T+����|���g?cƈ]��@nT�(���f��<��d����H��A��F�FȆ��S�Ǧc�4ޅ���'�H���0�0S0-��z�=����?�S��_��Ѱ]Q��=���>�	>b�N��%v�Sj���\2/`�h��`#�F��Zs��0w]?�nu��V�9�?��V�<Rޘ��lD"�/N�~$� �2����j���J�ϊ�JPB��W}v��7x.;i�j�Q��<@S���scT�a�'�Q{f��8֪	=�۴6�yםe�j">���]�Їx�B�i��ε���厛n�i�\\Z.W���e1���%�	�����*�k>v����t��������w������+���O6�v�i�seF�	���l�(�/�mr�wv�	,�"�mY�'T�ar��XAr���4>��&̓f~���Y>���Gσ�x�]c�c�g���{��}��o�����֭�d^����� �~u��Ul?	����#b�Ch}Z�%�����
��)�a���������
W/ǠePv�Q�c��=ZHY��g�zQT�o���`��!!�a�٘�*\S�pSC��#ZN�-��i�/f@~y"� V�(Wr3Sn�sk�Ff���~��s�30 ���9կ[��«bf2��{�1�1!�U��Y�M��m��b���A[%��~�p�e�9�pBٲ9�P��!D�AQe�]��KE�R8?��2��"3!p3.� �B�Y�S�M���4Q�ÌX�1 aͬ��B����r!V]?��Q��R��z�Ȯ�B��Ex����,.y�ZPyU���]96�D��0$��o� `�r�`��A#����NY�% ���� ���q��N���`�y�8 5]3~����`e!�yIC���V�]��KU����>Q޲Q$�E�����E��C�Ir��W�Y�]M sZڝe8\�������k��I-�󽸿��u�M��Zus�A�6Kj�(Λz�dar�Hp���\K���������;�eo�<j~iMp��3��6����q�Yֹ������i��u��Rx�`a�5��gրSN9�<��/�w��U\�c=��m[��%dr�W?j��������v�˹��;�,�.mH!��zV>RRPv���=�ts9r��r��e׶���պ{�{�FĊ��,K�Ԭ���=hfp����c�h����ޣ'��7�L�U��Y=�3��Csʍ�����*Ay3�Lx���G�,D�KӐ{5�cѤy֤1֣��$���ޜ����={����Ϫ_��w )~�f�,I�65~��'m�z>�l�_8��f&����>��"��]u��\/z�S,�7ҷߎ�	��B�O#͟W�$o�z���C�ª�	B93�;�,%�Wj+%ج��>�� ��-��"*p�,�"3SA����uN�6Rj{*+�ع��_�����2���Xpt�R-�i���f��1��f�,��z�����[,�D�X�����YaW��1I���Bx����$��}��� �FQ�@�o�����^�牭@ŉu����|�
�=����BM�v��lw�r!�}��P�`" ��11�6�Du�1BN��� T����'�e��$�~YЭ��^s�ϕ�GqU��2�`!Gƿ�E�P��M���.�9�׀ň���;Ŀّ�&'�����R�D���ۣb�0�g���/���̂�-R$��c��]��H1q>\;ˢ����e?A	2+�r������FC (uX�^����0@�1���C���&56��ʟD���\k�v�k�7B1�	�l����&�~��Sl�\�lB�>}�k�Pju!�Ʃ����P����5`�{���}�K�Sܢl|�'�և$������։�p�`���7�0�r��R��ti�_��ؠy���� j����G�
0��}���O)+=v@i��ե���NI����σ "���=��rm*_�2cM_H��d����K�W���Q�|����="�}w�"#�X`����y�⒋ڛ�g&2�r��֞��&1�M]��M�+�^��ѓ�4{��=8�wL ͏3��pe�9��p�)������G�L��#[��FS5��_/�����f桞�qM�s���J����qۭ�/���(���g��u�f���/����a��/�C��t3���|�&��\��F��ޚc���F��{�`�Y�u�A�6еt�YQ�����:�墎@TWg!.\52f$�`���.}����(a��u�)\��+n\/,�s�Y	�'��s*H#) P���.��[jw0���B?אav�XO��'g�K�8��4B/���}�'���X`�ѽ �F�3�E�.�<D�D�9�cT�m�FF��-bp!C�^(\�c�Y?��Tʂ�:.h�n֒�~�J=����J
��!�r����.���X3WN��3��1�;�bX1Xb��Y6�G��5����D�״��%1n* n.j�9�Jk���LW5��/��a|q��( Ee}��c�x�`7"�Hԧ��*��ME����p���ۈ�ͱC7������y�Դ�{��(ߒ�X5�O�p#s�n�6y��K�K�r�{�m�λȜ5����j;��b��n#���4�bt�����I-Tc!�!';�s�g�kTc�yl����U�]�I������ Hce��ƀ��������r��m�hǈX��{:'�"Ƙ��X#��n $�6z�	��� ���?��'	�<�"v�g��-w�&��z
��C[����+&Y� ֨\����9�bgר�R�!ˀ�9��(�P�d�t�4u�@U���_�H���%�*��'��Si���9�3���:��έ���ۮ�٥�V�k��Sv�I���MN���ܵ�u��AaE]��)L� ���.lV}������B����:�c:^�j����푘�q=�Sz�E�D^�0�@�yi���;F����~}w1��=-�|g��.�o� �maG�'=}d��}�5�Q���6�7��ޮ�e6���L��
U�d��UB�̭Z�z��wꁇ�=��	n1�Z��5Ǳ�ڙ�j1bW�}Xa���԰U��={mb��r�E~xv���홁"���퓗�<gb72���� ��z*���"�3N\';�q�lk9�\1��`��$������N>k+�ǎH��������a�N�a'�Ӡe��Ha4���o�v�<��Q�� q�
����oټ��`B�/.���93\O�E�#���)�5�S��`��C�		L���i��2X܇� i	*���Ǚ�TB����@;>cl�MCBԣh�+C�D~�Pr�(�6�1!��=C�����K�6��+C�>8�5�T��f3� ��lP���lq4nf����_�T���p�nC��
���6�Oj��d�0ܩ�q��\�w��$��ݩ��ڎ����01 ��`�]�{x.�������nV�}Οs#�,E�K� �1�q�<E0�� 7�	2��W/����-2�G���B�|_��7'j/�6H�� ��{N�����au3 H����sJ�Jn(x� H����n\w�u�r9N5�X3wn��4}(�n���\)�Ї��J�z����2>]e�r�9�h�z�X-���;��N�/����v�TT\�+�������=�����ԧ����
�Ö���3E����+����7I�<973���;��ؽkjnJ��-sJ͡�unJ����a\hf���gi���&����I����Lͨ/g J9_�r�j����������֏�j�����o�����9a�ZE�k�$�W���6���X|ݯXA����~06[p>�L/$$C�������].@(��=�P�} y@��s�ߴ3�eJ-��ј@�`"@!��,�$�Nh�&wZ���+�ɕ�_c����q��[sd٥R#2J���r��
dAC{���l烵Ц�2���0�m�ŝ]L�o6Վ�F>B����#�}�_�����dOfv�9%E�А
�R40�	Q~ ؎�Y	��b������ט�H9�Ō�W��Ϊ�W�-P�����-��e�M�?I�a� ��0Ҥ�m���x��٭51"Q6%
Fm�ۅ{1��Q�o�k�K_S�=��,��� I�/,�+�{�[_�83'�YƽKF��3�x���#r�!�U�^�~��JȺݮ�*�~�x�T���D���1�0��)!:�������Y@�P��p#��9�Lח�ߐ�j�H��Y����g�* ����w�սH f\��_�9�>s�~E�߭�c%v��;D��{�Q�CT�^������ʫ��G� �'�`���� ���d���@HX���7솎c~����T`�L4��cC����1��殻'�c�����q���zp��6か
�>����q�2��]��M��ǅ���.Q%�J�m
9g�F�C���w�Q��r��ǔ����9��E����g�"
/����ȇ?̌���|���\����5�����u޲m�J���1�u�Mײ���s��A�o�jW\7Qg}+�	ýLAc�U��nrwu�M<἟Y��'������,<4��$��":��S>����fB1:а9� �)�
4��Ր���~Q]]#���q�b�a�Ij����:�~,H����
�1� ���u1��B�;jn}L��2-�r�Ѧ&��E��vO_iV��Z�Ě��TVˈ�|�lA��sfL_Yx]hSL��3�mj�A��Ȁ�9�+�	�O�vU����u���I-XD�E]'j*!vh��D]+��V�}ø�q���(�5,����]�!#�Ga�,�d�&�G�#A���V������t�,��RV�l������ʡ�Ӹ�^ppզz��p[-ފ�!���&Ѓ�i��A-��qR�^�@LYgF��`ȴ�ӏ\5���|� *��%6Z�kN�^�H�[Q��lR��4�}��ic��(T�%*QQN��Ui�=�ZT\��0�  �*���;lZ8�I��
t8t(�]�� �»���C�NX׬Y��
�Rd$%DՏ@�����A�&�W�~&f�E-�UUH�&%����xRbě��41�S$z��ʳ1*���KpB��!'�=�n�~|��������Ăp�ԝ�I)`�S���6�H��:a�HE�KʸØ)���A��u݇Kd�H�; p�x�Rp���\�t\�,���g�t-�U�m��~��z���l�K�賌R$�r��o�И!�Í�����E�1m::�ĭ�`C=;�	�]�vX)7��ğu���+�+�W~��5ɥ@5�t�i�]�$���zr�S��q����&���oH��Q�Q�'�Y+0:��6���|Q��6+}��q�'��=JܸO)%��?�׊��|߫2+������Xq����>sfa�?f=��c�`�����0vQ怄�5ח_w�D"�Ljb�������kMGDJ�Gi�)����M\�n�a�N��:�DD��'�/v�Ӕ�Htu�_���9�\0EW,��n�^�@����Yg��Zv�~k^B���O9�!�VL	�����������3,�2 z��MU�.1�� `<�����ȒL��
�߸�|@�̌��9�c ���E8j������]�ڟ��G>�����C�=h?F��	�� 1_V��>�Q�Z�ЖK{aם�qGya����Z��@�{H����t�߰CZ��2�P�#���Wax��& �5A$�Xq�Ї��1"�����g4Rf���
E�	Ɩݻ�zڭY�GQ(Ww�"���N�dR�#3sɂE(��EF4�I|02�P_����_]`��o�Y��RG8�b���`��U_9c��F�!�$���EuUq���{��%���E��WIW?X�ԉٍˆ�^;�,��byX�5��(:*�7�6D'���(��� �\�Mmh�6q���l\[|ϕ\p��&
���7�G�/���2�\��]��s���I�s��y��#�<�d��*��sr̅��۔;�_�zy�c'O]2%�F	���=��~M9Qn3���A�(��:\����l��������ԍs���wͳ^�Kl�Z׺tyYջ��a]����~�Fk��Vj�[������ڴ�(�G؝���A�a��>o.������:_��`-���O���K�Ԩݸ����{6�6(bL�v(�ho�arp� �D״Kǔ_�{��`d+F��/F%� ��xY �s`$Fw�28:b�F�\2�-b�L���.WH*�3��	�ЧqC�Q82�W�E��^~|'��oY���� �ES��i���}A�햱�z�V*�M��.-�,��p
�-[��]L��1��R���H`��؀\��j�wؘ %��������~ZY�Vn �-b��  /e��D��ukו�����F��U
9'pH��h�uN��܊�:���Y�	�	�3��X�aX�$A�C�RM�5�W+��6��$EH�q�ܮ����'@^�fK���lW�p���� v�G����-P�AtD�\���t	q�4M�lٲ�Y�!��=Dy�`�l�a��7fNqU����(�q��,��������"�4 $bޜ�hY�)�1	�8��B�s��:i���2z>ȭcM.��}�縌��hb���G)�|�]�'�t�57��O����7�G{�8W�����z)VOV�k��Eغu@zq�s�y�Hj^g�!�v�]E���'=ɹ�`u�%�&�'?����}�s3B�^��NP�O#��vn�J�0��y�c�Z��CNi���	�X�Ʋ\�7�>�hi�FU��*/�p����5��s�v�_��aΝ�Z�@th��>�&6isb�F�r6��CG�蔫�˕(�p����C{*�Y������������":���0��� �&�ҹC�Q�0a4�`�{a��`PhVh$���h���g#;������jË� ����b�NI�(�H�^,"Z�v���z��N9�e(�,�L
,��+{��R�
_��\��ػgo���z��"���oVE��N���)2;���4v���i�^�pQ]�u̴��v%��8l	��Z��KeX�1N�j߰n�����fu����`Y��;`����wA땺�F��]:G�y@L�.19�(Wʄ���=���˥�^"�q�r�l��a���%C�>%��6k/8 n����]��'�- 7�d�#�7eIb�)� |���"@��"^E�Q��?�A���?g]F���^1Ǔ}��T��cN�D��<ĺv[yΔ�n��|�_,����A�~�ܮ�����+��a������fƷ�A���̂�+�3^�:EZ \Dοd�� Ap�@��O|�Jhy����^6K���c��?��r��T��ps3��ݬ8�[�·���ߩuJ��<�/�^F�e�E�
ox����k�i����v��/��G�N�� I&��s&�I�'�w�K���s��O��f�*�F;H~�3˜��۽|��_��_����s~ٺm����g�ē�v�aa�z��`� (h�8n��-c�$�6�.�d��{+Uje�uڨ(7�zs٣5g��b,��y-�94�[�}�=I�Dz�a) OWeOO�<H�����vP+n;�oFa�d\_�D	�3�6���G��Y����=����M%�I!,��tdT��C���x%�t(����cTS�T�ֺ�蛵p�x� B�(M~xP����~Ƞ
���W�\CcZ�����@a D%r�m!+@P�&�KK�dN�׾����x��y��>�h�O~��(�'pСE�Ą�s\��;W��6�$�]Q\F�@���>�	��E?�x�"�F�W@�ý�����]P6m�Tr�C�7ܨv�6��я~�|�ӟu���64(�@��e�=���Q0SQ#A�B�x&��q%��J��+����YgA�$���הo�;����.�[�6+Ae��D��Bb�l,��a�vb�I�X��:ܰ�Ox�C�p���y��(/��x�.pّ����q��j��s��\y�{�+Q�v�t�%��\(cya�+jӹ"��K��(��Yើb.� q>�э���i��_��r�"������|�;˷��-�܇�)ǞR�:묪�R&��t!��Q��p�|��B=1sF�N�ӣ�>��$#�n���}��o�+����=���ɟ�s�{t��W�^>��U���o��\n��k��`^Υ�a>�� �d�8ֆ��¨�������o*�{��̚|�0� ��Y�����5O���@��	�
�D�_\Չ��P�y��׈�c��|�����|��Y.���b}>�����_(^|I�� !�s�4>�@�mĦDz)�>K5��EF�P����ފħk��c��i�ֺp��7I4���Yܵ���E	��*�=�vz>�~F�'�>�OaZ#�W�A)�G ����r=��dL������&�{��w}rC��̪/�ǡ�~�z���OF,���G-d�dy�YXT�25��(�A������Ac?�Y�0��z`��<W��֪��L� ���x�a��%cW��(����;��ۋ��c��M��}�-�Eь��f����ɚf�3�(\ﱳ���>�Ϟ�+�RViW7������{G�¬�N�?t3vi�v��L��Mh��*���q�л`lm���Q��;E��� ���/��\tمe�c�O�'=�g�㽫����)�������J"<9Jg�� h��s���>����?�:�s���} ���W�,檩���b����~����o.��r�2�����>�<�ϔ� �����W�0�E��Sb�N���8�7�Xd�V���y��p�J�N$�E]T���>*���c��6������� P����>��t�D��p�Ŝ
=�ua�IP���h`�4�� N�[�9��L����*���»��.�3�:���MZ.���2:3R��x�����=��h&�mDv!��#`�yp�3�׬��_���9R�q3Sl�c���-oy�ٯo����o,�|�9���//_��r±�;�h�X
'� �]�Y��dGV�ŸD2�2_`��|>V�X�/���z	�/��²{��r�
�����q��%%�
�;�|���%��N�Y���$"8+@��H�2�M�ܴ=���sIʉ�E������|�_q:4i�T��y��}��5��	6#]����o`����:n��W�Ĉ���S�y��̒��:a�fs�D�%~�siwf�(��2��U�N8�2�,�o�Ԧ�U� ��@�d1���Zs�Y�>ǂ���)�Et��E}F���S\.D+�?-���$�3X2���Wh)j��y��|��j`4'Iag���G$Z_)��|�B�ךw��|�h�FW�ő:�^ #�� 0�����X���v!�۵��%$=u>��0Z�����1T�޶m�w��׭+�>�Q��o}���W#ˮ�Ӟ���{/�]-����P�~ja������5Qf����sF-jb!��q챻5���\�4��З���r嵗����m�*�-�)$�?�6�+V��� �4Bڳ�C�V#�n�
T�'��t��>��{��q��»\yQ���/;���3�(_��ʍ��X��������/��8U���W*��܏����-Q�Q��@�evC?�n�4������������Շ���T��'>�	�ÊR�lذa^��C�n���`���p��7ㅻmF9��ah~��'�\F�b�)�p��������90t�Vm*/|������Z�K*��� �3�����A��5L�X�t�)¨2�¯v���tDy�K^b��[�EW|�lZst������聲G./X=
�f�-Ν0�"�_ͣ�  ���o�Cߥ��.�Z��t��@�s��g�ּ9�s������%D����p�&�.GRD��s �֯��Nm��3���'������ek��#��-�� 
n�g�E��O�W&���t����]2㙿�Lύ�r�1q#�U�h��-��pR��w)�{@c�};���)��<�X�?e=m���|=�w^P���O+���i\�����y�Ѧ)8�[�<=l$t�ZFHr� w��+��?N=��s���(1V�>�y�"2��Bñ ��
���F��7"ن\�,�$���h8j���H4~�0�hm��ūߏ>�L)�\}��XY�fU9�Me�Ļ���j�Y?�0s�=�Q����+_i0�[��L��򗿬<뙿&�i\�k3jwIƛ�<`,-���87�KU�k�:dkn&����ҭ�Q�-n�׾���6�ַ��r�uז��#W���!��{v��zY��%�J���+V�Qw��zP���u�+��h�P�
�K�V��w�m9�r���_*/}�KZ~�U׸H)������@,3̈́0<j�����D�!M`�;}��n���a��o������ovx9���J�.���lF�x$ӕzG	��Ꚑ�(�T��yE���fH�� ��s�u@J�G��g�g��g?�.J)�v�Z�9	q:�=?�*�k��e������a�O��3��m��~���屏;_���o��mxO;����W��\�2���n�A0@�`���"{�y#���?la�Sxm�����YC�t�a����'�׽�u������g YƈW���:Q�=Ϡ#�"��8�"�^��툣�>�y�s�� `���������|�|����&[��N���Qr,����!�223b���*#�m����f�����кW'c���x¬c#}���B��2e�?��1��~��Տ�����-��vq��"��](��FVYm�4S�70B-�h����,S&i6�c1X6.Zx�������XA�7X�0;)M
ތ�v�z@CC�����1�����)wL�4��ra�A���P���C��gA�-`aA�!�<�O���'��c�._����������� �T#ڭ�u��]U���ᢘ��Jų�+�����׾�<�)O)��r�v���EB�5`�ڤ���Vi�F�f�$p�!�J�D������O�)�B�۶�Gi7��?z��Q_}�U���?J;�9plV��i�ltL�L�4���թ���e' 2#��L?�+ƵO;ߓN<Q��A����<�)�U�z�uS��}B{Ө���ŬScU]f��b8�_�=�[�7ƕW����;��y�'&���7�����L���N)�5\�>�e���Q����f���
� �t4#�~㪠>bQ#��`��@�r�<��/O����k��N�㖲jժ`��W��2�!�1��Kw%�]�js��H����I�.F�?�ؾ�i���)�́���e���H����<|�1�k�U��������g��J�� �{�_������8��V���W�O��dܸЮ�$5Kk��_�j�]��F���
Q�\���$mUd܀�9�5֮�E��k��*t<v�Ƌ�y���eG� ���Wq��|�@Q�"�D�j��$�ޠT�5����r�r6FN��} �b-��Ԉk���v���K�{Q٪����m$�Zy�z�t���Kz��c��]�'����j���XA���bLv�ս��,-RH�Z "��������@��?�i7��S�4o�ݔ
0`sXib��ѥEN�,�{�;˙g�!�+�\��;�nw.
�N)�N���FgU��]��c���n�ŋP�G?���m��#�X|qP�#�8�l�r�Ԛ�Hݡ�~"�������
����V��b5%��
N�>L��E�P�nz���v�a��u���E1 �}ܞ��%�a<#<�b�V@Ye��wF��C�uP�����c�H�~�`a=�łq�|-aX�X\cA�i��`�^X�4���䈢���>�*���o|î�
��B�:�0��`gޝꢛ��<4ڜ���� ��U�v��ۑ���`<��J(H߂ȗ~�I�1����ZD�NnT��k�(s3�3�,�w}�P�y��n��R�Esf���	�a>r�5�\:r��r�^f!2lz����|����9*��>+ǜ���߇������8�h�F�q��\�Թ�ݵ��b�����}���Y����D�)W���с���h�����W�!� (j&R�-`j�6�ʚԓ��H?��<�7)��ǟ����6ou�V���+��Y��kV�&�U,�˒�J��{D��{�z��?�.ߓ�Ɍ���08��j? K���� %���N~�Q�]����_���1ю>��ث���k7�#֮.�ܹ����nk�.N�hmU$�zp<Z[D7.��=J^� ��ڔ�+��C�Wc��;����+#�E��s���hG�����������;v��Uu��ԏ�J�to��7�w+�GG9��ːč�e�B�^'�d��9Y�O���sb���[&������8�@p��p�R4h������O�t5mc�Hُu#s2e( .��`�G���\SEZD�#��T훝��yPٽcgy���Q���z'r��&����Z�T\J�p�e���˖�{��	��;��py5�2d2B3��
�t����?B������nAeܽ�?.P��U�7�7�M9��f�ʈՙ�������O�!�/��@`|0�����.-��a����~��}U�!��V�5�& C�SW�n9������#<\��8�0@�>a�M�)�F��0C�b7���b��&a����5T��7��+��m���r�n�D��Y@;�̾�� ��9�����x�)������-�@�|���U>�W����;�<�ɟf��>�r�񱰙�lxl ��s���^��Gc��Lf�IkwԞ=J%���E/�}��� ��HGs��7������Lb���6Z+��D�r>e�p�M��Q	�a]���0�$���d�fܡR-Ѕ~��%n엾���Q�>�����.���g�>lg4@�j!���R"g�ϥ����9X{���r�D�9�\��&@�`��q__�L���R6o�Vz$�n����C��X�^v
��:"ti�W["/$���L�����WJ����7�������τȫ/	 [|���":��FX"��=D�h�70�.�0
���߬v~$�?Oc��c��,���F��<�.�C:{Xv���O+�=�Vt/^����N���q�-�v-�hH��ޮ������qS��KY]��/eFm�Q�UsRHD��7e΀[���*��J�`)ιC��n)�ַ�?��?�����w}@: ���N@��?R�"��DEA��\@L�hY�]��N���������WJ�i��3%L��׾�E�.���f�5Y�^%�C\:�H(J�ȅC����WA�{�\1���
 �O �����ay@��G�������Z.a���o�^���~��ڟ��g���R�����t�2*������
1O`G ���W�A]�DY_�#0�j����|�ϕ݃��	G�P~�E/*��0�[F�+_���P�@����b��`���	E�����NJ�k�r��:@����P�åyC�D�Q��8�fI�������S��d���_�z�K^�1�-��w�y������6l�j�v�b���B�|,A�1.O@9�R��Pz�Y�?�hū���T����|�3�g���7����;nuH�Źz�)�k���'��a�=�@��	 ��`��S��C�����o���t���e/~i�9�������hJ\�_�җ�7�PN�p�F���u�^c��Z!��Ө ~�� Ak7�9�ŝ�Åf��n�Hv�M�^0^��V�C�X�}�k�y�=߮�W����VQʀo�������E?�ݙ���P3�5�������])�s[������������������4S�G�K׈��\��q}�8�7�ֲ�@t�۾��p���ʋW���r�� �6��ԓJ<׳0�*
�s��y�a%����A�a���Gs��)�Pw~<�a�Q�;��7]S��
�x��ӭ�,w���N�:dG� �f�%t�(e�%�=u�x�_��'�jG�����;.��k	���NHfbbT�e�s�q��c6���S�i�>�B���(_a���
��� )UҴ>1@�U�pǎ��L�_�������?Ӯ�k��/UD�[�t�)'�e����˺Z�.�S+�+����r��LJ5�U�b`���Nѡ�h$F���?p�~�#~�C�+^���'<�|Y����u�/w��p��?$*����EB��q��&��RV/�h`�X�c(\`�p� ����ժ�m۹�,ʳ��[��������c ���߉���w����o�v���m�������˺�X����<?��0v1�j�ժ�Q��믻���#�ź��g�f�%E��^�Gv;|�;߱��Z%�2a	���Q|�+��`�\��/ ڬ��ss2�v�B�d �Ec1VKpt�ڧ� D����g���e��!	䟾�O�^\rɥ��\v��N���I�� �� �w R�ƜhBv�/Q.& �7$�������a�TDխ���?�1��/{�4Q�ʕW\��I��?x��������m ֗a�()ӯ�~�-��<rn1vu������jT# 
��l������C�:[����D>��϶�mo{��Z�	�spۭ���֊�"8FS�gk7$�`	��L ��{�3�j[�k��S㣠��0D�����E���V��;R��8��.�`<��qJ�Ԃ�0K��$�&7}r睛='tփ4Ǘ��%���`m984(09��P�s�r�qh�hC�9�rg�ah���Iz�� {�uM j��m�����+��Gʵ��Y2�kc7�����9�&)3�>/���� �0�O_�p�F�����̀
�A�N�{�[�M3��3���f排��ˢ�?�E�[o�N=�+��`, �U�:�zV���as$�X�~eq�$z�ݼ�B�)�`#4W0\vQ�����s�G<��7~�Y�x�p�1��/����o}K��eҥ��3ɦ�s�b8�X��.�;Ys�y�h3�E�$��]G�E��uQ2���4�v"��:�(�-g?��J�xC9��W)r��22�wlw$���v�T�G�Kn�X�3��� �G�?F� #���1�ʓ�~�~�������v��;���_��[7��~���ƀ��8��D�s	c���ꀬ�vs�(�:�g�V1WC|+ )��N�K_��W����S� �
:���+^�
�w.tDz!����[�x�� �s����LMQP���2YM\9�gK�B惎�Cٲq�!C����w(_�-�%e�"˙�5� �ח+T��5��mZI:�bOm(�C�
�+�D\7�'�%�C5x�~����׼�5~���9���?��#���W�D�p��)/C� �n��<sV?�D�֕�B�˔�q�>�Q����|�����v�;�=�O*����f��Fy�sQdX��E�ab�5��8pa�0.N�Ȅ�� :�s��ҋMS��ՙ�?��d��="�8�5\�h�.��b��>�_zu�s���p����'�p�7i��q�#��{��u� I-1D�T�]R��|v]�7ma�P��2~��H�:�(9�B�am:�]��֬��CC�p_��MS�O	������X���#-�~�z`�`�'b�	C��@�n,|�Z�겘��=QP��Yh��E}���>���6 zX�� PiZ�C���[�a�tZ��:�,�-�d�v4���%�~��*�b���r+����;/v���p[�m���ؐ#���-�'#�J߽��?A��s��\aoV�X�Mb���V6�2Z�ΪR���QIQ�"l Z�%���%���H$`(���P���<S9_��^֠�UJ������S�?($�O������T�q���J�8\`�aa�"�md�cTH�3�9��c40��-���1�?F"�#�R�s�dzYg�]�E�`�ey�pyE"N���yFL�<�P$^Υ"�ӝ��,O��':̾����w��{���<䡎�!�w�����F��|]���{�O�hv�2 ͻ�������$v��{/p"D��q޼es�V׀�qM��RGMP���q	0+��n�T�	�3
���#a��*Ր�:m �v�΢'s�f��݊��y_�D� .G5
ppm4-� ����i��2z��@��#�=n9W�B�G? P̧��x�y�JuL�����Qp����  05����M5�=fVt��N�1gYWߒ��.^��h�����p�gh�R�}���v�#̝���Ĺ�`�@0��s�B9B�؀*����A>�� �?&�C��\����&�Eg��LXƚ�:��!3��z���J⇵��g�C��(�k��:`z��el�D�r��U�����L�?6>�4>�'i����� �Fz'*�|��cQbMB)���	�7�!��Kc���H$b�db�p�r��+�6��qhfp%i�_ w�>�}����U�<�%�t���}��^q�ŕ��N
V�.,��;L�+Wh'�t�,����a�.M̙!��~z�����B�'����
<Xl�F��� ��)\7z9"E����T��ڽ��?b�M��~� B�ǔ��,��2��L���𰢣��.Eōi�I��ԗ0��O�u�K�=�x�8�
���x-W�V�c�b��	Y�=y�&�5c���w���v8X�{L�Hm�o�!���fW��M
�����HװOb���G�h��"�vi�	��V-'L$�#��#��0��*�4S˄��[���[2��燎�x������cj����fn����Q͉ A0 v"�2/�(�y�Ffm�45� X�է37�J}�X�)����> ߵ�|�	��@0N�MhL��qf��� ���2�	�v%$�2���A�ܙ���I[̇ ̐�B�j�ؿß5&��YȖ1��M���戂��q�����Jt@A�ٝ[��e�Ll�S'�7�&����1?�w��)�������и�g��>f�����ɕ~�p�r0Q�囪�G��cUw d��2eCs��Z�t��&���W��*�1X.��rNٛ6i� �������p٫��e�V�Į�r� �6"�#��g��R��ĸtO[�����5=�C��
pc2-�_6.������":�!����l�{r-���n�����t��9���8ޝ	����6�4&^�����xSx)���:�@�����&J���N�hOSC/2��|�k�co�%�Gdg�5��%�h��h10~�e�r�h�X�K
|�N&PC�@!�����H�����Ȅ�P�\�rx�������Y���)��\@m`��,��GwM��tT�ay�U�v�;֕W�F��y�m "x��6ch�RcJڶrx���.�.��"Z��1rfO��[ ��jL0�y&���+�`9��<�h7�@k�d��p{f��.��%䱯�1!}C�p\;�� pFj�0���,�4m�	W��M �;t
�"��j�	�]վ�G;"l;��z"Tֹ9�c;��*B�)����B_G�� �����\�9�9���!�%�W��F>ª�O<f�N{0���5a��&�y\tU��閲[G���?]{�\w	\q����dv��y\�y�e#�'�lK�=m���pvm@n�mh�iQH�YO�8��8+���K��pң��=�� ���l �k2��� ϊ��EYK�ch��M/0��s:r!��˼�T�*���>�A�%7�W��߇�����	�צyE-<�w�ޝ.��W�<�o:�E�Ş�_ ��ۍ�0w��˖�S��ψ�Գ�v)#�sv��4+y�]G._�~獷s��7�g'gf�Q�l�h�li�5#?Z�F��]��g[5�5�x&[�u��\-ad3u<���g���yr_��p��?T,���C���rO��"
�(jZY�t���{���\<Q�)�Bw{A�h1�7���Xd��#y���"H�� )�$l��`k�Ң�-���(�97)����eK˥��3�h���)�V(.F;��~h��P'���w�͂�b����:x�E�0"T�Fl�:t �6�&�ȶ���܄�g��a�C�̮��t��໬IDw�ؙC�[/T�C�&�7��nt��i�W�/ Z��Um��0�I'��y�[�Cl.��q�c�${=ae�_T-�� ��(q��e %��� ����=�F80,�h�ˋ��)-�h� 9�֌/@��XK��h|�0n62�r)�?�I)���+C�q[9^R��Y}�k�e#����g��^�gou��Y��*(��\JÜ:�t�eC��1��f@�4�W� 
���a���eܒ�3˨�H��kFPp�8��P�;�S!���P�,�+�}�o�4g`)���r���*1^ ����n���> @,х��}B[�,�cP��S�M"X�x�B�,}��>�˽ N�4`��u��^�vݼ����pO�7��iS�u�:�tS�
�x�mr��Nڻw�>��8����.�Z�����((A��I� {�;���_sF�kk׭)�y�RJ����'�)4�w�ջ�v�l���)��H�/^���/�Wm,���������W/Q4ٙ�iG�����jmj3��F3�E!�M�OM+��&Mk�4��0ݦ����M�?�z��kVϵbP\WrN}1-Q��9/�ֽ�+JoLc�8BJ���1)VSt�dOg���s�nk����6���������֎�aٝ���W�����-�ց�0e?�_]Ap�o�7����jL?�a�̏b��.�{��p�4^��:��O��4L��G�I����r�5g�bâ�]����
�;k/�=AB3��D.� 5Me��:ch��G*{�J/��c3���/ᦩ�A(j-fֳ�EHu��s��JhBT�=�:��a�n!i�v@ l�ݺ6:tF<��4�S	��u섄ڴ�s�7���w�n�
�! �k��tR���C�1t�c�}`Z���0 /���ON"�V�MW����`�~Kf$��=Ɉ��2� �4P�G�n�EZ|���?���I�.������� \��С0�Y�
&�����&�g �� �2;�a� ?�f�1���8�9���{�o��H�c����0y�q]��\?���id��9y�K'(���_���wf�n�y�d<�ېJb���$���;��,�#X�(&J�16 �F捿�N�Y�-昣/+S���c?��`J=H����b����s��/#�`WiO�DĄ���ql�~��LJ�"c�gn��"A"�G>�>-���V���WX�GAT������5�K`����u(���O^��*S��=��d(}�CU�1P�ʭ�3�� ��b���P���`� lK+�:��&�,���6yy$���w�q{�����ܵ+�ꤞ���|\�Be7f[�ȸtQZ����M���ilxpE�����VLu4��j�X�1���* �ǈ�l��J�6�Ƥ�sOb4db� ?n��-�ss�L���M�qff5�4��f���J�ߥr8����Q<��QC�y��sV��Y�z�����:����,���_Ѧ5��.��W,����]G�{0 ����=�@�������{ � A�OCC{x/���Z�F:=AP��Hbw�k>Z���i��`Ե��������\��oc3k�0��ᅒ��f��j>FCoe���������j(r���	uȽ�{�u"̹2,�wkDD��M��-j�S�t�^$�� *M��w�y�܇������V�<Dh-����O�c.�c$d�_]������^��9U0�)�M�D�Ic`�*����>��4���ۇ{G(�
ظ>�k��� F-`���HX�­�a�9ҝ���J_3��،��γ~z����Nc�ȅ�����`�5�t�L�}���_D����e��ڬ =@¿����2]p��o�D��*�q�@��xc	��c�}g��=i�pAu/ѹdx�+�����!A!mu~J>�0-h��C�S(�:�<��X��p_�F(�\R�N�`6-wF�q݅CF��<�;O�p���>u-�偙��������ј���`�_R!�Q��J�:L�~�`+��Ql�ꜭZ��T֫�TO4�p�_�V���\�A:K	�8�?ֹG�uH7$׹/�\h����n��Zbb� cb���K��2Q*�GJ||�[�)w*�ę���.��g�Z��:N��	����_9�Z �=��|��,�l�]��}@��srtBd_GG�ܧr����=g&pz�)�<� �ʺ��\ϼ�� ���<f��͐]����:�O,Qn)\O@�ǽ�,�kF���}���Z'��Z��o�c�_|�>��"�O�t�aW�vl��4�@w�%,��2D���7�	�hI.:<�Q��� f���صZ�"�Ц(���ף�Ŝ�p�B|����v���w�e��N������f�� ���&��!��̑��7�*�S�T���]ka�VD�z��n�i}֦v���umNXp�Gϱ�nA2O����Q&]���O��1��NLnTF����9G�ՑY�޸���������̦���ۋ�o[f�&$�����ٴ��R��t(:שF�sY�+0�F�Q@Zۤ��H����(�a�W;Ӎ�@1~2:.k"a8.�0�a�X�C�5���}���Na�r���ѷ}r��W\FP%+n�x�[�c�v�v�[)��[��W�^�q��>%�Fk\�z�]D��wiI�Ř#h���� ��M}�J����eZ�K6,����$Kb�
@��u�<ȿ���>���쇜Şy�F��ĭ��x8"K��ui�#�`	`�`3l�
է}z���y�h� �0�c�Hj(�����|�䠿0��7' ��좋�y��Q2�ߑ. "��6�{!���߸Ϙ��p�X���oJ��=�}�Q��R�8~D�d �1F�J�h���N����$�}�ވX�r��(��M���/[�s)G������۷��ؽ�ܶy�A�I����>�6$���թ ����x����H��%K��?��mV�f�VN����Jsrv�E:������z~,�ieIP�X+d����1��ߛ3MaJ4k]l�&bnvttnrj�����Uϑ���Y=6�*������Kc�{��&�=�[�>:x��\�c˶m+{z���t�MԿ����U�����[?��( ��4��!�9����[�Z�o�O�n�6PD��D[���=� ���%?�<���`��o"%=zv�l���ʲ �PH0�諕;�a>�lP������Z�0���h�csy1�
����P�ι��*��Y��ܷ�'�|�$j�a`6�^uY(�b��ϭ� 䗐n]�s��`�O�.�R��>�5����hR��<����f̽A�� ��,�����i�k���s��n�-s�F�)B�c�4�����ǘ3�{��¬��^F��,������r�l��s}@�@���c�(����}�ͬ<�ݕz�������+0)���x�h>Uu�3!�q?�d:���s�8X<�\�+�M() %��v�c���܋��ȿ -�Bg�*��U���*�_}nh�ѕɪ&0H`k�	]�@��Ww��F�4�ݷ#|46_k���d��?�\g<����#p�����ɰP����F\�&*�|U�7@R �n\���c���"���X�ڗ��.�-���2N0�Y0��ʹ�d���pUF�
��u�h?נ,�Sq�ޘ��^vi9�ӜHQ\ߛ��|X �(������;����w�( ��v��Qe�7��nO�t|G�ɛ4�lǝx�˭t)�]�=|�yڨj~(4��Mt<��r�)RlF�.�ы����][6�ݷ�i��hZϵĵL陚��gRB�I����x�֚&�f�:�U�\i3ۦ��o1Q��L��w�A'W	��ix���M�3y�	��
]��3׻l��1%����t� ���Z�w�0�\Gw����n~럽u����*o߱����bݿ�"��u���9�hT7Չ��4U�?/y����7'JF�З����G�"��qg�A>��ߔUD��9�R�")p��
QY��â�wn���+�b�@�*i����L1n����ؑ�B"�v��O���R��0FDaq�v-�?�3,��6x���&��:��BR�Ӂn� 7�lZ�5�t��2PD'�7ax�c�0l, ,89g`����ݧv���0�ܻ��x����ݬ�.=��#!C��r�z̓=c� �H�<����x��y�.��Y�p|� r���r����l�f�[��O���ܗtvi/wV�����iCAfv��ĥ�{��F���p���	8����ȅ+��0����%'CJ�)ݶG���> �ǐ���{]d͚��א'���s��8�Ϯ���ܰ[T�(�P�J��2v�T ��V+���Q��Ԇb|�tP�`z4�Z�#�"
,���5N .�?� �!�$�B�n��Z�Zc��U]P�q�]����'+U�o�����5����Y���Pb��zZ:/����02�>��0"�sa��͑q�0�r��s^!�1�g8�&�m�Z[z� Q��"SN�A3b�FT��4�t� ���޲��b^��
��OP߂kRm��r�-�O��r�
2���)O|�T��(�ץ�1�N���a�t\�Sd�g3�9��}�� v��Ng��3�Ƌ~#�&%zp��k��HC4���)J�g`�&��ظ�5V�]UZԗ�
�z�����Ǟ���֦z��I^ׂ�k����n4��̤��M�O���7�� 6�Zg`�b�0i�]����"jKԢ9�K�jh�ĵ
�=��U��.�@�9m<��z�dwWOc��=���7~t,���G�z�v)L��b�5�'����_�ii���f5Ɖ���t9���ֽ /��7�n4��j��XDxNà����"AZ��u´�A��Ov�z�j-�wo/k���#N9��ɸw("l�έ�̳�p��	r������/�4��W�B߮��42Ƹ�X�i���%J$*�EtF	;�ZK���bZH��ު�\�����l���)|'��}���]��Z�`�� �'��!1Ȅ���h@�o1��++GB�9��^Չ�G0���`mt���ݸ
���E���M�� ��I�"�}�]$����lۈ�act̰�H���U#ѯ����U�(�}?��psoD-!���*A����0Έa�*
�93�zU���.%~rX��^E��ݍ�S�9r��xh����hK����׸bq��D�@����ɸ��$���#I�(pe������d�k%¬��Т�x��,٘� O�h-��.N{��\/0Uu�^&�A ��{l�yf�"�ML�*�@�R
��d���2�#�>� � N�����'��eH�,1v����>E��H@=��`L6�jd���'���$8`*���f2{6ü����L�r1�)���;�|GlƜ��?���7d����?R#�a#Z�y��P��=�y�#��ی~e��T��'����(��L�Ђv�$�=z6'��0?�>���
�ɺթ�3l�p��z�i�"�]wp�U�+��X���ʯ��T�F'٧m71*�t�y�
�t��;�)�b�5��ɤL%�-�z4���MO̖�#x͊��҆���2.W5��1��R韶�ܫ9��)�}�lKSk�p|��X��yP�C�y��e�k��E� ;�#�]�"3c�f����\@�H��c�RT�q��%
`¡l�}mN.��Np�hK���p	̃�
�,�s3�Y�q'��w�_���r�QG����o�cV��=;({�]��ǚof����R��L�����-	��A0�]�$( �T�I����j�s��|�u�T�/"giFt�=TmJ�S0g��c�(']�#��)��ΞϪ�%Ȍ��ܩZBv� N%��� ��YÂ�'�JF����p!dY���@�����[�0#�����$���ƫ0��~l�z��7>F�U�9c-`kw��.�pO��=�q}*J;��q�n0�	��[��t�����C�Wא��4qs�#�O,g�q��!��Pv�T�W��e�ve��Q��8o���U��\h�>� �����qF"B������,p=3��t���6�Y��2����e�gTs!E��'��GG���-�0_�Լf�ý~d���b� �r.x6�{0��#ڐ��|F��vPi ـT�84@0��>�jm�Keu�l2Y�!b>��m�r�hS`���r��~�;���~�Źs�nϣtq�e�Rϻ�
Q�B�X\�f�6;�R.�f3Y�}��$Z�V>���(����Y*��y�:�@����pX��W���wP:�f��1��?0<�~��9]�X��d	`;�Y��Ir-�'h�"���f�������R	0�c�3$X�C��X�����53>�?�|kGkK�X|�T�����?�r�n2�]�Ъ��{��;�Wa����>]�G4{�y�W��3��id�Y�M���e��/W��������׾�\�;��}ʲ�\��]*�x��%���K���͡�����,����DF�pz�����0���+�/�S���a+� `r�ȖcYd#��Zb~�|.$A��7�g�`h��qI�u������LFHi�
,�%Z�~ff!�<5=nj^R?AGd'k�*��v�~j.��i�ÛkVh���/ʲ�<Q+������V�j�|W�J�3p�ErJ��{`���|�`�8b�m�d�Ȯ����"���T��s�qB���P������ɪ
������gq[�}Vn ����ӧ�#l
cn���v���2GM
j�KΛ��J�LH��'vT�^�i�t	�� ,��� #���滙x0�gy��MWZ���vr��L��85A@��q���\Y�H�8>��l}�w"�s0Hb��.8�8��Rk�nK�� (��yfGs�,�\�䍸�����g�O���<��#�$�1�(C�������)�>=Od��(�&J�gZ�y�;�s��5�D�� 7�A��h*�"w� ��_d\S�P��=�
 &oD%2Z��C�q�Pр$`�sS'�tR`~�V�̵�?�,/��y,��� #�2[�W#P !���i�����6#C��<Gw3O6�h��(8e��kWHV���A"����MG������m�*���W��R�WE�[��lF��\��F6��:44aT�
�
(33Ca���`f�pD9�����`���� ���,�hKԧ�D�F߷ؽ%��D��M�^#�j�4<'j�u"jTjH��rB�q;M@�A@��:v�+C�3�s7������ �C�
֊vf����
p�4�}C����eU��@w^���Z;R�5����C�Z��6�Uw��V(�HF�:gT��UU~_�~�ڲ_E_��nh�����?���I�@ ,єF۠
�%��V��S���:��#���V@�h�} �`��1��J�@p�}�Ѵ�#�^��>� b[�6�r��E��7��r����ՠ�K�=/�`��0[�@�v��H��2B�ӦM���n�%=�Pw>�Η:$Y�W2I�+���;.Y����Mmwm6mn�h�8S�����LS�?�7�s83�f����p�n�\K�9qe�s��o�UN�fm�V{~nSh;l��7�,�nf�߰�Q����{��O昂~"=>����b@�(�(o��$�JY'���"�6��Svj�6�s�g|Vc<���-��9�_?M=���h�4kQRГivW�F	w��ŧ�:U/�Uא;�\��O3�n��O� ^1ų,E�� ��������W} �%b�.T����
�d\ݠ��ZyE1I�R�d{�6��{e�:��>@�i�\�`D��ˊc��-'��r�ͅ��X�����~r�r����7�u0�|�����"M�2��8��HC��(���1�ac�lE�~����cXls��龎��n5Y'W�;\��PF�OV'ٝ*V�Ҷ-��Ic�ƕ��}\/K$0p�Tƭ�pfi�"�q�Xԉ#ÐEdQoB�e���p��}��j1ͽ��ۧ�7���q��������A\j?��-�N��?�2��[����z߂i�	lٺ�!��Q�@_�`�����(����ka@r?B�����L� �t��|�J1oӵs5�4�J����c0��c��W���-�E�'�g���"1��<���H7����T��̈́�-T�qnBpK�EC�<�.��K$�H�|��L��������:{f�A�uE};�,׊�& eu��>�t�9��>�ktЛ���!!3����;��c���UXh/st떭���.��Uש���Dc�U���ci��޸�C��Q��U�Ba�N0��P�ճ=FrC2�K�?>AnJ�Dy!�4�"TW���_� 聏��@s-z�%'q"L��w2A��n�L���댙���J(�P���w�-��(2���@X�b�r��%"[/MQ��\t35���ErP�-�݊���]gr���AJD��XT���Ż�LU�٢��źJ����k��b��pa��
� �%��п�{���O9CH�O��}h9��$�^�H�D���<�h�������y�Qdqo����ܹ�~ K���-����>0(�b�Ƌs`4�DaT�!X	X/"~0�yO�fg�7��)�e&��nk���xF��
;�yU�S�g����01��+U�;�9�C$`l|����w7i'����_���d|�\W�Z�{�XJR>�;'�$y���¥O
I)�:t�sNs&Y�dW�7�u�J�M��Ƞ��'�K�{K�"�`�s'��\++�3W���$�LSf*N<�$�1Os�-�U7�`�1J]X �V�[�6	��!�h����\��$�*�/n(߯�a %�(5<Q��N�66G���\��g n�("LٍА�π�d2�����ϙ�����=߽V�7c�w9c;��]�x��;KE��>�Liؖ�y� ZbiF�<�g��'6!�&�#�w�{G�Q�p8Һ�N�u�8���Ǖ����T�C��Q�Q�G�K��_���m���Y��7~����6/���� ��W�`U���Ñi8e��F$Z[/L!��>��Ǹ��H���k���n9�-���.JbE��*�t�_ީň�M�Mc eo�n��7lX�Z=k��v�̳� k2q����ga^4Q$3v�ro�#EN2�F?o7���#�3Z �ó1��� �����v�E�Gj�>L�;`���!ȕ��r׎1d׊�)w�!�U!L��5cH�<�����qs��w3o
;e\9�M:��4�
F�,�@�T��x�u��GD]���	��{�J�����v����Y� 4C�3 �v�H/U���Ũ��Q���煱A�f#�Y:JO��e0�#�0RT
\�("MȰ��w,��U5>�1�6�
�� �>�7�U��?�c�'@Me��F&4APjz	�wj�K�2�']�K(j[�g�z}V�t���yM�$��|���&��ۄ��|&�0�Q��qA8��H�G��O] ��AK���=��މ��꺌	��D�K3��]�^��p��k���2',�w [��;6(�+J���L7X�9E������/��9������˳����v��իW��N=���S�R����9�xDy�k_S��ǖ�|��J�y�}µ��)�7�v�o�ʘ����v�^m��sOt`Xd'����k�1UDf�@���4���ch���s_<�M,F�=С0�A�Vr��� bծ��6���ڨf�^�|/ڤ�����!�uxxB��Ouun�7�̪��f�0���#��L��8(wҖ���	ǝ�]3�iІ���0a��2�-��)��i��\w�,�)`�d�C�)h-Ad��Y>��z���Øu��Zh�m�x�MS�$����0;>/�����!�����i�K?蜸N u��a>����
�:)�9��)����U��]��R���dE��;l@�ݡ�Q,0r�J���T�B��( ���g��޽��h�Z�	���Β|0�(?X�HD{a0ƕP�	$ɩ#P�ѡ?x٠j�$`%�L�Csn3B�`#�k�N�b�uRj�m�Ů��r�۩�NiX�e�n#�u'�7� �Kԝ���b�rӯ���Ξ�&���|N�0��F��Y!�͈�=�BN��Y�q�y@#�E�����@����D�U���	]k��mkF�Yg�4�h���r-�1�FD��� <�����NX�`r���W�缀j�)-���A���xv���W�˦�2 �am���^�(���oh�"zrґ��@5��ɒ��Z��<���F4\��lh�x�6n�hWn�n��|�K_�Ɖ$�0��+��ԓ�)�>����_Y�<?�ڐ�ls^�,o�\`M�2.�aD��\���U�(���i櫊�����En{��]�4cc-���D�1<?��Yd�����R�����1�.<��|8��<P���6�+��d4X�����N�x��Ϊ�׈�����P���"-�9�2X, �S�}��E~��g����bM��1�����ڐ\��a��®��r�	� ��횯
���'��Yޫ��H��L�:/�G�5*+D!Lt�v�]t�Q�h�p��06`alc[�\ 
'مԠ�&q!���E8�1��['�S�H�ƥ�<��g+Zg�<k���2XQJ���|?vOx��0f҂�	��ڔ��/D���Y�7��q 9�+�_wݵ��~�.[ج�PqJXv� kv�w�q�˯�_���j�	���X@p��W�Ez� ��H�Sۓ�FF6�]?v%����6pOb��7���<s���ΕA�mH`�����xS�Eh<7A�|ޞ�R����4�rY����zX:�(�B42�1ܼ0B�9�XZ����F��7��/ܓ���<�!ժ�E��z̨ P���l��L�Y�s+]�#W����bc��s�C_g:�����W��o�Vey�9ڬK�|���eZs������n.?���GM��/+�����*�Wܴ�͜�樲��k�E��sĜ[�k�5���J��ҥ~�����H
ݦMذ�	�&kڬ�Yڊ��{�������c=��=ЮtR�l�vyAw���6�G��J�BR|���QߋE6���"���>�ì<�9�*'�t\y럽OƎL��%&��uʀ���g�񛔊��r@I�f���F
V�Z�Ij9�P��[O�sL����?�]�8�~Ȣ9.��@̋�h�q\�
�05���6-�U��1eOypt	�>@��!3�̤�-�U� v&5�����S������@��<� WU�L{�ݴ~�:�ÕLF�D1�3�(��_�$	/���Ds0T�ci�[!H3`�.3�- ���Ťy`�̶	a����D��F��BS�4P���{�SN-�|�#�\@�h)k֮.6�P��\|���i0R"Cv��1H���bu�o�=�	a�JR�t(;�<��<=	�2�<�I0$	R��ioj[�ա���Sp���Q{ӥh�۹�3E[�MLA2T��t�W��"�/�QE���Q�|U�ZD|����4Z7Ui����i��3S]�m�o@1m��7ne\n��ʄ�[�d�\�J���9���r٥�5Ks�ǘ��H �oc��Зըˬ�\�ṁ��5*���Q�zT������E1�w�G>���g��8��1�)�M��ct�ח�|�[�K..��Y#fH�Y����ISVe��)��O!܌}$���T����6:�18��P��
)�/���p������w/������{`=�!d����f��0v�0*r	9��u%��]���}���K������H��4;uv�,N���w�W^U�Ĺ2��2� '"@i�¸~�r�-���-g�ur9pp�CT3�cK.�I'~l�=����^�Hw������cw��L9�`N�/��<#խ�;�f�G�p�TF$�H�q踒�Bࠍ�٥����� 9��ΓU�'��å��"�Ti�w^�I�1X.�!��kV�I `>iu�� ��0 �n"�"����1��.�RF*"�B�E�asn��V�2c4^��K�>������$ߦ�D�;�\�h����s~c̸w�'�a���`���qS ���_��cv��c���'��Rf������~��V~)D����r�" 9�1��ZU�`]�%�p��U���`ب�΋�ѷ��i�Y?��Z�ψ���չ�wy/s��2`	���[8c��H2�G� ��Z]ɶf	�d���cT����,����A���"����wfm+��g����)�Y����3Y�!ږ�,*����r�E���<�bA������o��Z:�`�g��.R��b4+�:��>F�=:sA}Ja҃҉�~���ѩz]/|��*2�h��'�ɹ�����a��5EO(/~��#���򊗿����Yt\��0���q�	'8���n��e��4� �c�=o�?Z����VE�]q���_���e��3i��̡	Z@��i�]<�ǹA�=꿨΋VEi�� �h0P�����GQ�f�%O�B=�z��i��Qĉ�,ɸB֯ۨ��l��=2P�BZ�ĨM��g!����.���N-g��`Q�se�����M.��AIڪ{c�n�/��{�Nh�)�@z~���Re�Ɖ�����:K��J�����#�� g��5"Q/�?����i���Pu?���u��jakR1�cd*����ݫG\Xfd�kE�+�2�	�5ە�vF@�M�t���0I`c<�q��4���[Ɓ� �I��[9����]�i��/\���!P�M�Mԗ68Z�'&IN�NI��8AD���#�kF��r*�@9J�2�|Q��4������;��A��%�|2��.��o֣�"�*��W+)�Iy�����?�� �e��O/k�V�[o�Q��l߱]�n��a|\�Yms�
x�U��O_r_f�H� �&�T�)=�6i��>���vQ�!��v�7�C�D������h����~ m/���$�R��Ƀ�3Vh���x�(wrG�,:#�H�j~��[G||n�#t�y� m�ڥ����� �́%r�ڭ�����oص=�}B�ʂ���p�X��%��Pb���Sm"o�����,`�Pץ�v��{W^q���A������S9=���^ JPKK5v6*���ٯ�,p�c�=�J���\~�����C4�L�{�ψm:��%��I��lV��K4�>��O����-�~��+_��K��?��ҖY����z �{�E�:�@O��LMj�#uv�> �r������J��).~�]��-�+M��Ӫ;���J���맨A�l�Su�f�iղ#YT��`��Q ��t~������0^	x�w��7N��<�ܡ̬��EZ5��e�\&ZԦH��«�ӊVg��,�nW���ejh����r��.[���TX����fCX�����
����~�9;�Q��� ��ݞ^�?�Od�KA�0u2�T���&��	m�� �&�0yp��>MV`g��Q�WB/�vЂ��S�	���D�������I*3袴��w*�$��Mclw'�E�!-�T>GЬw$�kՂ�ZJ]�)�c*Q1�h���D� ����IQS�\�]��Q�t��b:'F�Q�P��eBQ ���մ�$l L�j�\c��/4#�+3C2��G�&�d�. |���
�?&����9Y��0W\�}e��ڎ�����(�E�D�U��#�в�#����^:U�Nî(E��!ͷ�졿i>G��I��0 �Ax�ߙA�5�Y�$=KRO�{��i�8�L}U�̙�a�@�%���!�+�v^�
�8��Ts��f�/��artg\3�c�N�9DS@�1\���� �#'�$\��+!0/g�gKĬp�{�l�W�4m�UD3���1.��
�d��X~(�
��o�"!�� -�N��ϪU�a��y�� C�U/�~]g�F	@Bl&\��`������V�u��w��{\��[�o�<`t睛ݎ��:��x^�6�c�:ʐua�@��?��_�%�ξ�q�3��H��D��K�lN� ����բx�;4��XݹT�\�����ƕ��6�̦��z�c�l�^���fT�Q3.H���OI,
��@������w�>�GP0?�.5� �w��,L�>����Av�i������;�;et,��ı�-c}��WK�x��]i4��0�.|*�3���2g_���D�j-غVc�EDQ�a�=#�['�0Q�
��@��9g�&��ĝZHDYc��
��e�\*�Č�/:���hV�'��r	s׵<������;P�;v�>�G��4_����@���!�M11��1���8z�� ����H.\�m�jf{��]@��Z%����3���,����T$6���r�KƂ�8?Y��sλʜk%�2��c9GQ}�Q�>�kP�_�t��#�BP�BE1�ލk)KJ�^��-yf1j�u����B/��0��#�ÑV���uּ����c���֧H���)��ӟ���ֈ�Uø9Ÿҧ��f���cT�'�&=��;����I�����m����,]�����q _N����:o��,���d�2.A����3�Z�y��:�s�2Wx���#w"k�W����}���p3F��F��mN̯��r91/�C�ںu���o���.fͱe�Mv����۲e��'�VX��FV�S`o�����������g?�ܥc�D��6	���ֈq�Iަ�����P�%��Lu�Z���cr*�h�ԥ�e����srE�j����63+�t�Ĵv�����Xd��Pk���qF2g/TwO�SC�z��a>47P,���`���$٠F@�2��⸅���f��"F�G��Vj'�e�4�ٶm���ڡ�#.~H�v�֓ஒ�b��S]�����K .���.���0z�J���]��������3�3�?����"�pUw��@������am��`42�p�p�D�.#���A*ꅾ!:y�|�fP�=`90��YD���MF`���,_ ���x��j�0��Y��d|:Čp��)��l^��"�a��\fc�Lک1�R?��Ȱ�����j �=�po'���!HrC��EL�v�s �0~0Im*J��o"�\@-M�$h��y�\ߠ�j���*�9��"��<I�b9�H���e�{�(,��'C��鋨���&���1�莸��?���K.�:7ʙ���k�Pi�s�ŭ�*�
`g6*�;�!����X����ߝ���'�4�eɌy<�S�@Jn\|ߺg\�fq4�̗t�s,�9˼�vtY��6�,Eep$��eɜ�Ṡ=K�*���&�&����q�b���B�\���.���D��>�;���������*aϾ�
|X�qnes�g�6�5-)�;UFc >l������[����|�(�77�8.����Y�i��:�1�S��	m�ȵu��t� ��sIY�98t`�R��-�sJ}�[qh�hW��T_�r�,�~jz`=����W�uGIT�o�ㅕ�H��@t"Qk#�� h!,=@ͽi�o0B7s�8ɞ��~�4���Xt��#]8�Ek%�UT�2�(P�΅h��e���d�V�X%�a�,��]���������0%m������o��~�ca��,��Ļ��棖��.=v�D��sgq�dօ�8F"C � aq���F�v���E!�
� �����L���V8"H0��6���C|����rX���xA_3���v�Ez��q{Tm]�� 3�]w��Ԕ4F�9t]F��s��.��,ӌ���-]nvg���b�*�J[S���8���D��D~ M�j�j��0��Li��VsF}�+��_��U��	)q�ے%��A���=�f�-��7�W� �d�B,��X$�\����P�����\c��%7-&�̃G�P�y�7,���ǚ��ZX�
�/� �|�_Ѿ�}@ ��|�&�L&7C~�v��jɒ}���.�#}��hf��v�7��{�$��h�O��	�U��ʹi+`&#iS�"><��}�KPdrF洳,70���r"D6#0�r+:y�ژu����f���y-�gnV��}���v��G>�b%ʖ�p1�g��
1@��=�v��~�ʿ���?�g����I'���c�W*�ǈ
�H��G���H��m��)�i#�Z��%��̜D�곎)"k��U˺��[�p{"/�~*z`=�a�a�;w�O
��:W�.����?�dq���o']f�+�Ʈ�gk�L�^ AZ�"���uk��O��ʄ��@Yrک��*`P�V�ͬ5�@� ��5b�"2�ňE���v�PqF#*��*�E��L���!���K��'��8\��QM���P`���U������M����){vc\U�[tt9��m�C����'�BAi�9Q5( >G���bQo��2#��WWS�aq��ާU��i&fO��ŵ���^p3�c�!hi�+2��t�"C��������$�CB�>�Qu5���6u����\ �&Z�r��n� Av� ���X�W�(0K�c�8���x0hcƵ���K]-���<��
�e��g�;~�x�"1�p=5�E9�p���-C�~��1g%�ձ�K{`ҍD{x�0��6#z���t�.i}"�LI��p\5�\��}�^�>�3�<�,P0\胂ť�N��3����&��\��E]�X t� �rʬ6�" ��Ͽ���|R����Y���Zh�̮DT!��T�	
��ؽ�`�\D�؆ul��?��C��zV5�hF���.�3Z��Ҩ	���[�~��y���Ψ;�*A��q&(� '��Ji��cܿK�{��n�x�*`c�\_�֬пr (��-�3~QI��կ*�\v��SS�L>T�<����(�LrD�'`ը�kX�B�ވ�c��ٵp�z^Ft?K%֢�ڰ"@�5-]�jtfr�@����w/���]r�T��-�� ���Y���Uy�֟Y�Y�o��̂7�)�д��S��	M>�xI�Zf4W�[�~ǏW{r*���g�A�m�ņ����{`=���|f�MYT��
� �=
o�O^�3�MJsɻ����:�)�F*5!k0��l���qtJ]�x�Hd��"�B�e�G�ƈM�NǢщ���
k�c1����e���!�"�R�#�d��Ι�cM�0<ZP� [N���L0F�2���K<����c9p��`���h�!�(�����5������W�#�\�M�a��y�Aمq����E�+Y�S�@ꬹ��;\����r� ��:�uY�#��53b��D1J ���7 �SQ-�p�&��<�Ŭ����G7l�·Qw�o'�����,tAD�	`�с��l�}�ƍ��E��WJ֗�aE���5R�X8	_��/hς��� A�7�[�Ȃ�5u+Nv��K�]'=�#��~�̒e��E�ʍ*� ��#,�s9�:�b�0'-b�U���rS7M |D����]�k8a�A��2�[l[�P  @ɐ�	WN�����(�f0��i�8�L��ܣ�վ���Z΂6p_��h.td�^|�"���Uq�D�#}�����4��k .r�1��Y��E�zn"�G�Gb�I'�l�\g^u�����a����)�5\W:�BԪ���%�;�Ĉ��RM� ��͹e��}������.')/��&��(���W�^���
�ԫ����R���Ǘ�T/��w��aH��λ�,�����#������	�SoUj�j�q;v�(�(���_#�NmV�}[�P/`ܳ������:[O��;{������˛;�:��`�Eji�v�1��kij�$�eNsxNk���V 3�-s��Tb�	����M�ݏ�� G@�� D���lJSlR�������>����뿲�[��њ8��Eӟ����4)@E������9=�S�ө�����kVi�劌Ea�u�z`ݯ�Z8ؘ�A��b��
�*|��+�`��{,A�}��	p�zj
x/ĮQ�'�����&q�K3���hؕ��c��"����6�v��τ ω'�\��DVZ��֒c2=��H|hL{ئ��&�+�a��Y����p�NWN��|�u̊@�u�rp�(���*�����W�8er!��*��P軴j��pu@��dKs�����t�R�� �Ѹ�����������.2g�óuo� }m��E�w��K�F9���7��_��dwϹ�_x����z��ﳋ���<~�?jv�}��U٠C�j$�f�K���` �B0r��qfgC��#�q��+5jo�r�,�����?�?� P�+5W�b�v ����C��>ùNu� I���+��R~F�p��0&�vSٲm���׳��dy� �N�{��;�� �s��="�l�u��Q㣎9��*�s�]���`�)^:�9�8�}�&
4lA������quz|��LYX����I��F`7mdY6�ӼD��C�����a�m�n�-��M
�1��,��A�=Ǽl�$E�C�2���F*ܖ��(M]�$�ݻ� �����s��\�\Z�a�>p�D\�z~��h�M�s�"�G�[ν]��˵�{$���䖅ɚ׎i3	c����i�֮Y[�R4٫^��r���f�X �$U%���6Z�s��ru�ީ������4���=��G*�gl�4�.��Gu�+�c�Ԏ��]G6�]���ܺjzjNI�ۚU"
tV��g(;J]6�����'F�gD�"S��bd���5+g��h����>�Q������8���ig�qїf�"+��m��r('�{����n�K6��o���s|���`��%7����g���B<�����=���kO��q��)��h�M����G�S���Xf�m��I�f���E&�;�h��Yw�)H]����@Mf�#J
@4ƸG�ݨ/4"��~-<�c����8��^u�D�BtV�_֭]gC�%ѻ]7����8���*�}(�����8�M�\\��X�p�5r�`�dW)�ߗ���J�xFy����ъ0s���.��)��!���M7�����-Ĺ��Eb�H�!�Ɋ��.F{kxԖ��dD��|����+�(�y���6���0,�c�A����Q��N���kVd���\�R&�����w0�>�>I��(w�~���]cD����� �r�-
-W�]p�bV�6co�	��xp~���Gm�a��Z~t�U��`.���$� ��AEf1�  ����_>��f�֯� ���2.v��[�Ns3^��}���s��E^��;�ӌ���:r��&���:ѫ������7�I��G��n��@hㆍ�B���g�
��B"����]C9��ǎ�:d���L|�3��&���3�E�c�s�?�Q�C�P��[��Y~㙿^���'��3�U���ed/�L\���)C��.C�î`��toW\~Iy���]����w���������̜ݠD���3i"Ӏ�O ���)J}�7�"��[�m+���t�m�(��ǟ�T�0�Y�9�!��k���7�5C�l�sK'm����:���.���O�Je>�����.){� ���s(Z`��z�H�m!c�s��bZEkOw�55-iokY��35;95�f���1���l��� �\񘅚_Զ@
?�f�=�����Y.�E ;	�}Nt�z�p�U0������fm�i��V�Gk��ά$	�W�v�ԉg�~��yȐ��_�<p�j���� �0�&��Nv��%2�f��?�u5Z�����P%J����y�����묑�p�X젆{���W䀉�:<�&O�X�4ȏ��,p#2��+���'���$��|��f��ŭ��hHFmH�׺#�Z���P,���hwyAy�;����LYٹ�>~7��S�d�H�oq��� ���4�R��o~�k��^-���T�[���jg]~�[�Z^��ז�?�g�nw<�mP�A�V�C�!D������ �F<JZ��8��  E2EΕ@sx�L���o�zWWw�������,��?+W_s�2%/�B�Ї>ԟ��Iב!�0��1A�=A�Z�'��re<��,�N�`���'�]r%�������s��\�<q��g�"xe}
���c�D�fs�@���x0������p���Y%�H����}�/^��姝rFy�+^Y�h��S@l ��LCM�`.�����z� ��/|W9�|Ԁܒ�����O˿~���ŗ]\���^^�җ���)e��@\��2"��������1F[��`&����Fr7�����gRWn�����<��ǔ��;O�㧛����/?����)�_o��g?����d D�.���[�顇�NųPۑ�B7�3G�VdK�VN8�1�|nڷ��m����"`����/7(�0�[���T���2 G�FBH�k�)�9Aw����t$$�6�80���	7#�0md����;��FH�<���,�|��5kVK�����z��t�4k�7.�q1T-]*'�k�T}P��1ԦO�1����隉���o޶�����O,l���.=�$�?K��sP]jQ+�ӡ�쇤�U�_�!���Z$�-H@���uJhJ)f%�G�꿦q�,�\[�d�@��s�%-�[յ��Uʋ��&1�Mڔ*�������EΌ7ͭP���N�ؠ6�A!�\|ݧXA����� ���Q�U�����L[�����l��W��n6j^EG��W�0�6�����ʿai�\�"�(��:���)�(Hbh�5��x�1�S�u��Ț�Bn����b���t�A�b�]b|?��ϗ�k��S!�'{\yƯ�jy�c��0Y��S2ر	ևQ&)�}�-�_s
��b�Fj�Ҁ(BI�w��]峟�����[F�Mox���*��c�w��Ю��~��_�N1
J���-\��w1,�M���﨤�9�h��\JΆ��~G׃��U��O}�S��`����7O~��o��o����P�0�s��7;Tw�����6n��1�l�w�(ѝ�9I:v��7,��_�:�A�Q����z�<G�v��U�o2`��><��$k����9�*���R3�p}�D���[���1jGy�J9\Z�+��s_��tZ��R~vy�+^%��,3�DQѧ��l�A{QǨW!���! HˬD�	Q7	%J�& �(��/{�����|�|�k_4�x�@ �����	m�/�5�3�� L(�}�.a"@�ƅK<\���nUN�}j�E߇�OpG��QɈ��/��Mo����/}ы�o<��]�d�^%��;�f�V;�ě���E��\	�����v_��.�j<b�._�W�����{�k�����g=�\p�N�@0ޛ����c7��tEE�f���EFޭ���&��Q�ct��ro�_��<C��==�����(�'��D5u�n5kss��ʎ�[�B��|:��qf�z���v�Ye��#$|.eUg9z`E�_�Z˞ܾSh#*�y���F�ygg�Ԟ��wL)#8���ۥY�Җ��`�R����t��^m��8�J����R��n���C��
�*`Ӯu���Z6ϵw�L�(�F��S,LO/���X��4ף��hS_��ζ7u��gm�T���x�C2'�v��_�� ���Et��,����0�Χ9R0FD���}���>�A	|r���?F�J��Q1P��F��2t@�����@`!���U'O�������ߺ��{�x�i�'�F�ta���X���u���r��w8iަ#�*��v[y�{�S�p��	�7�?����'?�I�]Kz�Bʑf앺�8�Ǹ�u~Ƀb,뽭�?ijD���0�P�W��6�����˵W_S���w�?|��G�5������け�#v��=�U��]>v�q��f���1��Q}a��44��	eF�WYk��|����r�i'�����=�}��l�S�����W��`�|5)(޹c���:w�I�9�`�i`�'��:U46D�-����s�9�%/y����֝[�>���O�����	,�r�-e@,X6�����Q�,U@��o${c��@���@қQXV�����ٟ�o~�>�)ǟR^���_{��wV�����}2�u��l�"MX���H��T@@^��WEA�
�Q`���.�{6�d�'�$�������s��$d���/����i�߷�{��<�9�9G �Գn��qt4REc�����5ϛ�= x�!�B�㔜VҏyHB �6lfֵT�<��ԭ��qLz�m۷��o�)��o6v�+_��i�V*,v��a{�8���"�����X?=;Vh�6 nm��B�T|�WB������U�
��mo+�v��!@���b:^���/|���"U��ߝg�Y�d�&m#3�� ����(�}�`.ќ8�e�|�	������2=���?��Ŀ�1_��/��������o��y�p��sŚ5/�{�C��uk���M�'!ǂ����=�ۤB���'��L��ic���T� ��ฺ��:�4=���h�l`S߯\��2SYkv���j�$�j��~��B�BQE���6�Y�\��='��:Ӷڊ3��^�׽���?���Kw'~r|pH&'L:M�s�������$C�$��=�mzJ��(-oa��2}t)�&'���bB����_����$N�Z�ʻL��C�@A�\o6�a�>��Ԉ1���DS�E����m,4��B�U_�ܩ.��-|�9��8�E'�-��N@A����F�~�����[K�����p��X���b"x2+)0(G_��2����1�P�#6}a�:�WT��ب Ԅ�}�R�C�"��{X�������Z�<�L�?>��Ϛ�MZ�y�?����#4]��j��эZ��6�.��b���$����6{-jHN	'ѯ��ze������W_}U���ß�����Oz�Q]��o�-�},�
4�Yt�^�M�@���߭��uFX0��# ��m�7-�����Y����uo|����p��x
Z���������X}�.U��RJ��ߔ�����`l��s{�̨�2mN�<s�����Έl>k١Ř6�~C�z�W�c���\?��O�O�&�(,��~8'�ɣ16�i�TNF*����pČEt��"pxpƷVh�jE������r��,:BcmSذnCx�ަ0���~�Q0 ':��ލ,�����bȰ;�
=o���x�C��ט�P1F�b�,��L�5"p�q�i����~�{����߳=�u�]� ������Q^ &Ԁ����%v5��6��AIF��}P�=����q]O�2�w	;w�1AK���������
�u�c*Z��
�eL]�[1P����9������jD"^�;c0D�X	̭����S2��K=�% �Y���!!���X�
���[��Ă�
'Z�p��&�@<'<���lN?�q	���zV�Q�k����;�����I��WBimhkX�5�84V
�L�h�e(�7X]+18���W麫�D���2�: [a3�p4��ֶ�0Cp�}Eo,��T�i����*`t����z��Aj���P�Dˋ���]����o�@AK4+,�V���� �8�s��|�e!&#��������Ђ�c��]�)�����`�0��!nR�k��#̻��7iW�6;'�`��h1��M'o��b"&���J1�q�&�x�#��C�S��v��	Q�0!����m��N �}Y{x���������`�d�j��{�S��r-�	�
  �	���W�N:�|$�J*�Grue(���7�Q��!�mwtt�w��]���H^��b
eX�'����}�� �<����`���!ާ8C�e���_'�Gv��Z/�y�o�NǴg�>�5����6���֮�HBeez��F��Lw1��i؊�H~:�cO�0^*'K]��}�c�G��V�-��@�bZX  �.�kC�l��Wҧ��O�V�g�LN���Aea-׸<S8�%V$o����#�/0����N�@<��0�ˏ<<F�^�%Y&@-��v?�v�.�[�����/��𪗿2�џ��i�(`��tl?;�����>>I�d@�h�b5c��,-YL���Mp�ҵP�c�ٻ'<�9�o~�,͛�%�M	5��d���_y��^RB����VX`����w6O��x�R��:> ᳔�H��^U4_)��@Mzc�v�1`�9�i	5��!Ȥ�[�f15=����+|�_�_wC��j�|���Zc�E��E��*YA���*��Yi	 �F�QY�:�)���7[� PT-cW���lLo�Cb�j[B��u�is9W�s+<W"�H�om���h��?Z�nU�)����_bd����ҕE��C"��e"h7��l���`���i�����pH5���*6z], !2d���lڸ��/��:�֨h:�CG����[mݟiat��RQT��|Ϳ�vX��nl¹N?�t9�W�g=�Y>�/T+ �c���D�q�
�%=���lI�G��l_��2��Z�'�2G�S�3\pAx�v����`�V%���h�x�'!p��*ɀ*kc���F��[ ��X������&�>7H�0%�8x(���_����H�3 ��.1Գ����m>TҎ���Ђ�:͉����t���b���s��}�mZg�r�SGȣV m�Hzk�i���4��ԥ,5?�	`(^kb��Lꁅ։9F6�O��իW��un����G�-�D��/!�;�}8m2�$
H�n�Rs�J0�,O���/W��6�����p��m��yn\S%�!��5 K�cU�� >���%���3F���@�zC���3��Ʊ9MB�+��2�1�>�g4W�p��`AGSa���(�a�j��Jsg1��J)뎎�d~����ג� g�<�+������{FG%*���8�T:֦M%����IB(�QB�Hy��X�]{wk*S=�6+����lEE�;�}
��ޥU �M#��oL�h(#!���]k
U
5��.�0��o^����[T	�^��AkN\*S2V�����s/8o���XɯG�2������l8ĹI����L�n".R1j��|����<5���.+��E����)ۮQuA,�]E��Vm���[�p�ֱ.�)�4V*d�*ۻC�:��H,����СA�Y�D�<o����G�'����
��;��賐�t�*�-x����S�ozH��zr�i1�hbV���Si��՚0ӣ�
�+�_s�:�U�}Ƶ'�v���R�9Ҙq5��u�pL�� Q����Ub��:OȋN��"6���E$4AX���l��y]PtTI�=,�!��7^] $�&���D�_���ݫ������>��O�hLH3M�li
�[�K����5�Ѧ��	0�S�U��R�;Y�vӦMV����
���1����z�i~��x3�4!�:\�,%���Yx�LӞE���d�5Klj�J�0Ga�`o�3��{D�b��r%�+���c6&M��`0�� +U��_������"2,��*]먞�q=�&��0��ZƖp��C}`�y���Y�(�_�m��Y�К�q��B�eec� J���^d�?�>�yr}��(9n=̖K���O�ح�>�ɮ�Қ12��}��c
�֯2 ��G�,��Y��Vh�8��5���5fn�b霚�V����*%ot:���^r���M��>=۴������T���>[u��������(�7�RY ��%��p�A;I��G��5+$�өoO]O/g��<�I�O��-�,D�O�s�Y����y�G	-U\aHn��v�ko���]�SB�i�
mU�����޿׼
u��x��(��RG^�J�T��bMEi25�����-#�^�ۤ����ᡧ���-��h�?B�I^Y�&��k���0YnҸ$�n�Y����h[�畧aU���<E��}��Ʈ�ƄU+�'m4�����Ru�.��Y��?Q����W��z���z�,;\��hH���w���jO�H�� ��A`�,!s�bw 0ǩ6�!�EV�L�T9٘�9����cQ��"dyHZ���~Y���9}cì։��ԛv_��	��|((�a>�a%�u>���"t34aiuq�m��?�����m�5.������f�ׅ���*L���\�bO����,%g�q0Ry���
YS-QT�ؾ�LiLW�\m�0��{��c-��I�o��ڻ��U��a�{�=& �X��&NN1ǙF����}�{���\e6oTfԘ�s꿥���X�V?S
��m�f�[���٪�D���4�3b\�0.󝂅J+����ˎ�⾱�G�i��c8 �ՎP����5���q��Th���?xP�̈́tB\��[���re��g��e
�K�#��a��笥F������w*kmO�Q�|,%��A�Bb�=*e��Nw^���+Wo
���_+E^i�ej�ºl�R�bq�QezOR�3�a� h����>�|a1ǁC�۲l�Iw�i��;��8����,&���N�N�qn��%p�U�b{NvJ==]��ݠ0ح��jq�*ղs�W=!�Â�%+6OftA ��γ�H�/vH[����VNSG9�u��*v0�B�h�_PL�ea��D����R7�(��O�L�ڸ�T��0F�¸��`_�#$��� �B��b�ttJk�"���:�<�.��!N�D�E���p�������_ �N�<a�s C�jF1V�W�Z��hhRE�n	7�|�;2i|2y8�48��B�{���.H��&��T�>a?>��[����!,�2T���q�F�K�V��< �t
g���`Ȓ�e1�g��f[ݨ�7%˘��\�>i�p�8�z�Z��6U�����LQr@Λ�P�B-���B�dʄ��6������i���_ ,�6,iNY֘��f*�c�b/�f�o��H�ta�3�}b S� ����jx��0��@����;��c�L`��ޝ�k���ya�`�x��t,k>��x[:�g��{��)��8��y�'1��LZsd1�y��z���5UO��m��:�e����Z���	t*�ӔW�3��?��OOz��4��"��)ՠKH� ��2G�,E{8j ��p׸a�ꉍJ'h����.U����p��+�?}�?Þ�]�6�Q��C�5W�j��5�r;��S�m���w�Non���������8�Z`%�DT�ܯ�8}7eU8�yr%W�9�'�\O�N��y�����b�"�E(��'����R{�RT�����k�AZx�G������ک�8(dF��
��g�Lm)�5^PB�8���Ǳ��>&-���>,ɀ�&�8Y,��$87����� 3�]6�Z�j��Tpl`l��Ο�EJ7UU�J[�y���} =
�����k(.��|}�̈� �����&���E�y��X�턔��g		�������cP�� ���غ � �� ����.վq Xb�e�B��\EP�j礔~�����g,�*�Q��|�X��㥦�	�azd% �~��= �ZckU��1�vP�$
��O���`bj~�����yy���,���Ǆy6),g� �̠��6�H�B؀9zqYX���5�盐S�o<'�HxU�����Z��b�3)��@QbL�`"=�b�\�a�#�7@�_�M��[z��S���̰1�P����kO�a/�Y���`����ÊN+�y�� 9p^��J��3mU|��=�浘�5@,F��Zix�u��>��G��j�ڶt�B����	m߼6��٠$�Xd}��
����A7TR�Uޫ����{D)���f�K��![?j`x�KW_n��P��2�!f��ZC���x/�o�u���[�w�7u�[�_�E�XAK5-�4ĳ�,�{*vI��.,f�.��c���X���.�3�"� �`q"L�:�yȪ��:�حӡDb�d-�4,$d�R�Q��Ѥ��)�sBd�>ȓHQ�Gk>�zP �h��筁'���X�V�A3#m4|�
�����u\�.Bl�Z� Mr���!4�^����hw��Km_D��0s���pOW�
-�T�P�L
���xS��	-�� r��p��R��Pd�w��F&��6'�k�Щ�c���9y�S� �rz"qO�z��K��"�lb����.^5�����{������h;�r*�w�
X�H��I��6�\a�O  ��3e��t[�@�݋�e���-��9ՔM��;�s>~oLU �p�Ř*H]� w�"-��6��0cccAz�q�Tp��޳h_�<$�	���XQ�BČ�%�b�*L�����q��92 !��5^��⁉����U�6�y���N��r��A���4R���Щ
	�A�q���=S�A���ФƊ2�nL�kгCr�=�4��o�xX=��q|���Y�M#Ú�B�C�'�R� ^����Eǂ6vT`fh���Oh�j��w�yW8�ÛCI��i+����1S����5>!F����eZ�bX96��*�h��-��@!Xt�m�+Ú�N��W
��BlϘ����R��B���H�@AKm�^-&���a%��1?�1&<�u�t�'��5���O�cL��CN�Ķ��7�&|�+��~;GC� ғU�+�	PЩ��P��@+U1�Qqz�"�+,��\��m��?v�83����. �-b29�D���5�S�K�Q�;:v�d���4=���w�Q�Q���^�	Ǐ;Z�g7�d�=����8Zf�y,���a+@f��^,R�χ&qq�mщ���I7�[�B���>vߑ���5�oK��}��y��7��&6g1h�'c✝��yR[cȘ��Q"(�eH�2�vW[��A��:6 �r��2 �u�0WN���|���SQ���Ƌqdl�����s<����W�M�#� ޏ#U+Uc3��L������yoe)�����9Q�P����
4�ƨ�FU.�_׏��@��n��t\� �\���ay`���J`&�͚��g�y��-3&y8��f�������y�`i�Vx��@��B���)�����;��+�d��٘iz1���e���#���{������.��xm���N�ْhχ����C��F1�e
��Z�\��NZG�drX�yM(4x5g2*}\׌�[O�1s��t��LϠ�V4"�Yh�s���
�I������MX�XNGs�M4�Uv���T��Kf�û8���Z ��%�;}��E�w�I�����T�O� ?���T3��K,P>����ź�k$\v���U,5RFBa�X'�e\)��zD5.Cǭ�-x��j8K�rQ������g�x�p
�p}Ik��O�<R��6��V�>��	���4Lp)�&�[��Sh���5\�!zv�쒓	���u���H�[�5���!��!�P�a�����rᑵ欂e8 N�b61�M@E�0���Y�L�da �*���ļD��Z1,:�o�����&\j�Fکs8���;�.@�l�(�5]�捥�+�Ac�T�29O�lM`�+�;;e9�̱Gc3��D��PQiF%������-��!�gc���³�����C��9�I�	�kd�6Sk�ڹ�Lԗ�����ۋ��Ľ|��Xڈ�f�)~>/>�l��d<\b��f����>~H���y����k�L����C�'�6y�D��J�O!s�.�-I��8v�Ҕچ�4N������͕3�e`�4wKsڠP�Q�w� �|���r�����tK���y����Ѫv=1E��XN�h�fB�F�+��!<%���
ڦ!S��ie���PѬH�R����@AKn ���&d�]��F����+�K���N
(�;��'��6��zBP���m�:wo۶#�t�-V�xÆM�[h�@�e�x��T�bU�%��ߧ�"���]~�(Mr�����ڽzuaB�r��{�Nӄ�Z�y!�MKB��>_c<��zM�`��T�����Cv��A�bIx29m���les���@�ĺz�����!���[@�Wh��"����DƒQL/�e�3^<͏U'ܥ����؝];��p�~���(H�i6��k"�@Hc�ӵh�l=� �Ξ�w�{c����8�t��u��a�)����l�����K9b;��Trމ�I��H�J!90�E �Sf��ya��c�%��J�i� �F���.$9 �Gۦp�}VV@����c���?kH )|EƝe2j�꘣�-��u�35����v���{[���J,��.n{�%��n��ɧ�b�=���O�Y�� ��o� �Tr ۧ��Tj<C���N�iKڌT��P��^��.��k�ǅg��9�߳D�>}��bk27�U}zLZ�	�?Kݻ�p�Ԇ�V�U��:���
1.WH��i*t�f�<cZVu���aeRm��䩭�Ą���gp:�-��V�BU�y�A�9�T�m.��&_���"����D�o'ydX ��%�3�0sr�(i�"SJ��h`�K��/�?�����yO�yh�Ʉ�d1ѫ�����b���J�S�y��y^�M7x4�q���?���Xh�Cc�����@O#a"Տ��ۢAB8pZm�
Uid����mtM�Ky;�6D��Fw�i��8��Y�q ���R��Ս���SB���i4�3�1�U�C=��֠����r�E��:䎒�^��
����Y��2G
��9ǥ��t<��7����|�SB��?���l��{aƔ���U-��ǜ`���ԯʝ���[o.9۽���:Yh3�^�c��6��J)�t&'T�!9H}�F��k���R��f��7�l"�DN���k�9s�~��R`�z5s0��;�j)��MX+���+��9%�ם��� E�DH��D�`i#]��f�lS��������XR0�j���f��ZS[a-W(�ȵ{�x��b �����b�A����� ��Y�����0^�@�?faY�LbMB�]>�;Qǅ�l�s�9�?؁2z��8}�TLP6�c[\I] 
ࢗB�Y��b�[aOke��Q�;�6!��w�czʘ��>)��
��ԉ��6v %B�����)g#d�727gTyZE �1ZZ~c���C�e��<T��t=e}c�̳6+��(p���S������tZ)O_��~o�K2�C���?�[�,2�}\��*5kEG
}����fa{hk�O,���p� h�C&'Y��s��&IG�2���py�X��?�c=�����C| ����Z*���&Y_��[�O-p,v��Y�Z�Ȩ����^��%'�T	���
�J�3V�����Z-6jv*@DL~B�V�̜�ZX�ݠj�̠܍��:1�!����B�.1Z�}��#��4EֿK��t��� �(�6��}^u�uUB���]�s���(�������vE<d�[��<����,��)p,�c��6�)��a�Ү��;��4�d����-�1%�
���s��5@(�Ȇs��S�I(��� ����y��X�ބ�f�,6�e�X�j}�\���Ӛ::L�'C�@��V)]��v�R���!�n\-�-��A0�{���=��3�9�8I��R�?m)|.��plv�8G�[��F�Bx0܋l�9ψL�S lm��,�rR&�EG4A�"�� ~NO8��@6���w�c�%h���Ɣ��զ�N�Wm(�Z��~̇�d�
���3}����SĀ�X��LKgE%��q�Ԑ��z~�<�0�����&"1�)��Н5�as��F!!��R#x1{q�z�3�2�1y0h�>��\��q��L'��8
�y�?B`*�<�k	k׫@�>�bE{�l���kDUC��3��k�)���.��y�Jk��h>w?����z.F���Z:���I���(����
vڦ�;s��Y�m�Ȑ��S����d���'���-��VN��"KZ1��(�Wf��,�S����O��H���Y	SYgi���VT�����"b���G�EbpD��Ic�(k-�c�:蹤�#��7�	�y8�_Rc'a��XM�+^|3��_���'�����ݩe9�˴� �\���:�&��v��<%6�
�y� �D���P;O�P"$��x,����{[ T�gO�Ŵ$�w�'���!N�6�9�h�>�ut|�\x�Ha�8�E;�a7��v��e�%ǏӤT�iY(��R���qL@P�;+G&Z�nL��Ff<���bEa��ϑÇÀD�h˘#n�/��X����Y�]#u^��\��T���#����
S�{r��1��)���4.q,>���_�yĴ`�ʅP�]����=ލ������ d�bj2�(���"*O�!z�U� B ���R��'�Y<�@���S�,L��}��!x���yd��+|m�Zx`�`I9�d�{��Ajݢ�M���p���;��9�9atH�7�*Nb�z/6#TxN��-��9_�b�{�5��bC]/�ؾ\}��<���������t?Sb+��T��C��{(�X���e8��>qn[i6p����2U��V1�C\�l������"΍E��w>���_��Y �����e�ͪ����t,���9�yp�p����?���|2�JZ �����(��z[����Κ�a�������Da�� L�zB�Sa7ճa12��T�l]���q�,z���ݸ�C�[���	�n���K�Z0
�>p2�p8�"CםD��>������)��Hz���iD�]��T��}�_�������*�j�;�_Q��Z
1[ۍ�f6'��i
�Y���r�پ: �2�gi�l��h+�ꌢ��k '��A2U���ݪ��9C�VJ���Z�ZJ���h��+��a���L���c�����k��O���ggb8_bK�%�����&�/6��v)���g؆Q�?�<dU�܉�_<�bsjߛ��q�������!�2�4�&��K�^�#�<��t��	���"|�O�\�c�F�O-I\�7al��&t�:�*zz@E	�l��jz>����f�����,4g� �7��2��'}� ��=&`��R[�poF�s�{���7g� ����'�����w�*��fݪp�m*�I�#5MUx�Fb4]ua�ºzfi��6�_�?[IP?->d� &��7�gA���X`U�ft�I�K����8�悼N�f3Ǳ�=��O^�|�o.�A���=���%�V�Wu_��\ȴb#jYC8#���ÁTjW9<�k,QK�4�v�刔Y���7�q��N3�H�a-��	Q=�s\��N�+����׀ӈp�bW��s�-��M��xT����ض��S8��xB8^�e��x��B_b}��ME��oN =���H��'2L��ς.�ݴ�zD���xD�� �!mwЄ��5���U�uE|ĳ���bz?mF
Ѧ�Ҭ%FG?�g��ɝB�bk @���#��l��N1���38!�����ҽ���1��0��Rkn ������%A��	���iZ���
4 ʱZ��jDI��_Pۇ0���a찏�nG[F����r��=����Ү��j��+  ��?����~M��wc�q��b}R)��A���C��h]�<HvЖj�-����}���4������v���w�zF���+\j� ��F^�M�҂D�R�x�S�����a�$8Osݴ�Uř�+��s��	k�Ú��P�K�]*�A�U����"���B�#�/���V�숊����t~/l��^,��i��z�.�xZ!�.�����}ž����g �x*>"�� h��쏸�f��փ��nYˈ2�	p���,���{�� #�#(YX�ٱAp/�/�({�V��k���1-bc�Y��aR��D8�l�E'!U�E�Ђ�i��Y�'��y���!��qH��4 >@����c�wM�9&�ʹ�Q���bт;��@r2��)�s���S�������<�I{�:4�F[�cw�w�鞽 �����l9�@hA�4q�<? �&�Lwoc����G d 1
dM�p���b>�����U>N��(
Gdl��1�ϓ�!�ᤍH/X;�~1#$a-I;X͝ �����AC��Xd�(Ð�#.w���<~�S�u�-�yikBh� W_����D���c,noS�y���X�L؋�Q�����#a: ��#�Q26����BPr�tN�>~�]�96��i��E&A8@�����]��ەЊdp�K�|MNP���<  �QIDAT����S���;q=p`�l�ݷ��g�{S��Z��D��k�������5Aw٠67�����;���]�����D1��#BK�T���]>L��k��~����>��F�H����L��[NSe�U{�-��RbbyJL��d�M�n��o�_#C�1��z�̍R��� �`�m��-��siZy�>�ZZ�3�_Y�d���փX���z�z�ƞ*�x�-����h~��':�%��?fv��b���0��/���Xf[�%b�#r��ZڲP�*��UW�����a\�[��|��J�E	��
\�;�K�W{r�؉DPV�OM�����(�?�c!�M��0�ʛZ����٥�:)�"F�M��D� -��`��V
��n�r�B��n�������Y&�93�#f��qn�8�Z�=$��އ檌��8@��,~��B�Aڴ��C�EC6O���N.�pR�y�j����J�휓(ݮ����{I"�W�8���W�;D)�ź��rCדBmV����<����#c�J%$@�8de�/4^�NfG��@+D(օ���!��P�s3�/��� ��^�VSd�&�a�8������.��v#��R;3_���� ��B�X	;�դ/r��6H�"5C����z��qc��c@��Y�l�,ܨ�_&\�qM�l���Т���	��;��Xh\��I�gDL)Lt�
`�l��� 6!�K�.�����NaD��k�BJ'�Q��C�:�[6�s�;GÂmUEZ�J�[U�i�1E����Jr*�JK2����6@+�c��e��蔛V*f��Y �]�-�ތJA �5��4�-�;��f�/��� h�cl���ؖ��3u�rl�I�CB�N>��N{L�Ĭw����X�ww <���*��u6�=��MW�֮�V4��?��Jv}�BN���V����$6(�M��$����7c�"��!˚��ݼ3ש5lE��5Pod�p;x?WI����/ӭ\��t�R��yZͯ��Ѝ�Y5^�C�E����4�>�g����2V �{eo��,U^Z+��؀��D`����~F%@V�l�-�8�$�A�P!��Wc@t����������bl�s�{1A��D�I���8l e��H׏�S�Ϝ�ۡ���#��<ܳe��H���V���&��>ll8?����p���3�ź�� �o����Mi�;�is�怋�S�yҌ%͜u����h@���vʘm���.������3N����UșK0cn�q锬J7 V���W�e\ʜ�t���ݴ� @Ș�]��O���"�SK�nѩ��أ^	��r�~�硒򤮕����32Kc�`�V)[��n�:+_���'M��Y(��Bm��A3���=�]ʨ۰~�B�{C��1��Y����è2� ^T��Lu�l��Cp��m�0�f˞��������0tlR�~��e���2l&��kQ��1} ��e��~�ᶅ5:�X\h�3�"Uka[쌀������E��eZ~O�<��֌�k�]��ND��[��Z4O',�S�`��\�pӍ7�Zo��Z��M��,��_�bͭ��k �u�צo��#�a!�F�*Nƅ�/��9�G�<s&i��-ю�z,�ӟo�I�����,�bm�ba,�)h!��n�@��PV���G�G��)��}.�R����M"tc`��|a�iV7{x+�:\��>Q(��A?����9�� d���� |��g��r Y8����7�U��75�8�g��,�ëÜ�@pN�H�9��q�~���C6�sG0c�$�&��YB˄#5]=���H/)��q(��ҢX�F���s�R�;ƒ
�V����@�i���:D��6z��� ���(�%������K`J�o���B�rʤ�{c�q���2��`>U*%�����j�9_	[� ��'d��u���l��`�	����]����`�O�8����Ш�6�� ���`%�� [�P4��0J�4�A���*e�L{)+L(v0���?�;ƛ�^�p�\�R��!c�Rsc�����:�z��G:�5�K�B`K�U���U��9�Ը��ޙ.�D����g�a�,/�j���@v#�xذJ�����ki�`���[������!��z�o�9�@A?���`w�Gm�׌�&�|Bl�A��c�"7�'�;5E����g���g�,{V^��lQ����� �>%Z�U��ږ)�L����H� �3y�������+�x�q����F�H:~w�v��K��S}cq�6�c%P�D�8+q�nF�nD�1u! j�P��"���Uh�?K�2O�aG*��6��NL���VցM�����<�ԑu��������0P�R�q��4 �3�]��1M�<���p{-F��gX ���?s�B!�"�gS+��3���sT��Cu_�����@(}�,��NZ*����*�04��΍��׌5�t�g_"p��&dc�gؗ�U�#4
�R�NF�A�K��ZN��,]��~,�^<�tE�Km³V|1�u�����`�(������З���n�#4N ��W����٫�;K�}�<4�s��K!2�?U}��5�S�i��e�}�LG�G�B��%7�j,;K��2�����Q*�#t�Z)�Y����1��[&1r�Bu�	�Dpl�?E��--9�doH���--�{�l!כZy����h�5�9j���1�k��U�m��P��ιj�
�@kvK�y
�������CG=*��Fj|f�C����S��0�?o�\��]Z+R����y��
�p!��ò�Y�2g<��FW���ߵ8��X�n,�A��<8��J;p���?�i�ҹ�G,lw~,��������p8S��:iE��Agה�6J�N�@͡^�T�U��De��QN�8m	��cD���ءm��"��_zo��S�ARdX,d�\#�!w���P�;i������:�F�XY`�Z��t]Մ��0�U��J�<۝ǝ8H(�ZسYv��:,��$�S"��\o���Y@)
G��l�I��������� �D����v�r4VO�ГbP��;+��D �k`^�%��.�N���c̈́]J+�ؔ[��|<���Z]�U)�ɔ��F�W��zp���o)�1۪l¢.Pij�3l�g��qK���1�H`dʰ7:�d=lF�kf�k�8G����	6�V���F ��Q�)�c�(�1F1�.�0aI��0��s����H
�p��I#Ľ�,�M=�`S���k�{�\����V�-ia|m�fJ�e�����?�{hnn���g�a�V��k�w�
�mٲ%<�1���
�}��{A<�F��8�J��0T�
�ͭ(���¥ R�"g�[�3�3k����������=�ݡIM�a�����+�g�s�`X�fe���������<��P}c+RT�K	 ��C:�dr����0�"V؞)�w���Dz�h�b!V[�";m����-4~�H=��6����-q�y�� �
�}�~i��X=�P�=� ia��8��pG*&�&~�%\_���l'Td�;����v�����;)}k�D�֎҄��Fr$���[Q4�ݺ%����i����ޝ���'T���8|֜���K±,�B�J0s��#�h܀��䜽f!�&��L����.��S,��-A�'��ZX��F"�gfḭ&.�����J�~P���ǰ*��3/�6����.&:&_|u}�Dৌ�����c�#n.���85�4�J���-rL,J��W輴,��/��v�&t��0��s�J�� ��؂6
���>+2*\D��CC���U����������R�Ī>sM�i9dKڜ <Q�,/�Z�;�I�XB��^��u`0:^jN�E�jĪ�q�Cr�5zOE���?�F�b��Π�%�a#��u �E�c�ߺ�j�'���:vT��1;"aJ���(<5*��3A��	�E�?%�P�F	@�XL[�����\���s�0$1m���ha;�/�1X`�*�lP�cY4 9�� 4O���<?z\L���[���v���Թ٠4��5ջ$+�B;��q����y�*K3N�q����@�F�{(�Ƚ�*nj�^c�uo��L��7�>ۣ�����p�S���/�;���#�C�ګ4�4Z�����o�!�ض-\r�B'M�0�~M�w����9�uJ�02@�n�Nئf�"xZ.Y*R�Q��_��������p�:�i� h�#N�<m��P��;M'-�=N�
}��z��G�q�WSN)�\�9P��dd?�l����J�^�0�#M��bѮ��l�L'��%�0�^Rx�=B� ����W-5���s_X��M�������خV��"x,�r���1%��z9&���%���~k/��݂37h����k����d�2�%����;����Y ��G@�'ڒ��� o��uv�ޡ�-4�ԫ�Ƞq�@0�.&鴨�bE�\x�IE%Y1r� کN�����`'l�KYU,�w�_�(ҽ�����] �(�F�0rh���&jt);2'uOh �c�����g+ ���u��gt��'����
�zd�M��5U
}(;�>b3��k|Z����po�um
�H'ҧ��5�Q�l `RN����2hl�u�d�x���0L-�=ٳFA�R��s@)�g�q4��pưڜ��a^��d#8�!U6�5�]�au�t_�H�̙)��
]-�la$�O����y[-䞻��c��a��Uw��������z���'?��p�c��B����K���a�f47p��nR�e�YE�3����fUP�P�xxX̡�dL)��_��	`�p��0^�I�X��z�YB��[:.�@ē���e`�֐�����s",H8p\:�	�|�BJ��:�������駟�ݾ-��8da�;�C_�Æ�kB�f�����2}X}]��w��>@e1V��\�o�>�o�����ϵW��|�������U
L�]'4�6l^jUe�J��<s�
#n7l�g�]��L��, M��z�)�����E�jZ� �G*Х{�>f	c�Tܑ��e�=��j��2�$��J�z��<ОD���e�(��HѴ6X	-�'��~,���a�L�jU��r���^dMw�N��r�H���lh�ĭ�|�C�!�_�1�t��@��P	9K�Q<�
,a�/�8yI������J��{m��P�:>kqoZ��:�[�sm_�,��/�b�-�'2l"�B���Ǚ#J��0�4��=t�D���√����c`����N�3@�}�����ўj�W�^	,��P-c�X&-��9������u�Q�m!L�BY7�;t0Nz�tbӡ�{Ld��ޮ~[a�5�œq�����-Cԁ��gt(?2VSad&u|��͍��;&�0(`�N�YΎ�B��%��d'shC �����tu��n�����2�-��Am�9�k��E�10�D�=��k� a\�8xĘ����N�j��#ǻ����尽�znM���ռ���	mI����nhQ}����}�u⮬�]��(U	��֕X�6����I1���i��ח1W*�  ��hp	ȢAę�/�����1�
�ls�J�h���>r���iYx�s�kl�{�Y�8�֛o
7n�{Nأ��O;=��e/�\~E��G�Z��;wZ�Z���0��")�� v�8���	BM� �E� �ROw��%�_̫V������d@`��z�C�Τ�����ݪ(s���L��S���V{
�J`I�ؖ�����U�t�2��n�N?����jB��{��.{ԣB���Ĭ��5�h|�ll�<�5�]ڗ��v��J,йp�!��{�N�b�"�Ê���5�Ņ
��[o4�����������7�M�P�PW�mf���>)�60x4,�0�Jv"����A�P��C;c�ד��ň�'S�s�����A؄S�S�l��zی������zkk��]��3x������ h�#��S*M*� ��Y����iu&���%�%йq��v ���D��ɗy22��_�����YD�c�"�Z�{^Xl��	Q $���^��A�`ט��p��k��^/}��ڥ���=+,kn	�ݷS�d��;C�~����D�sSr�bW�\k�IV.G���L��Z�r9�Z�1X�~���r�e �����b��W�P��9��|.�Y�z9�>s�k֮7��Z��ش;n�=4�n��8d��7`#X ��=a�}������!sj�C�@ȧ_�cY�L9@�p�T�"�͐�9q� ��a��p��]a@��g�6�_Z�c�n�~[0G�3:��̇��V	l��1��\�#v�c`��/�y 8��Ͽ��O��['��P�0�{F�J���V�����z�5�87�@�m�i2����k`�L:���
g�yv8���6	��۷?|�[�2f�� \z�e� ����ڷo��{��u��E�u�)ï��˃�8&43 ��Ί�0�&h�B*| AXj�j�lܸ�X�Σ��[�V���+��~�/9a͏�;�5�Ҏ]{Cs������B<G�3(=v�[��*5��wBk���燹Ch!��̢�Ȱ@��1Y�ZU�Hk�*�J��V�Bs��H!5l��{��\tX��6Tg^�y�Q"�29��^����� (���=��_ ����>�|�֍ھ��a��ճ��uKT4��(�2@�� ɨ
�b�P&@�F6���G[v`� 3����y�7��C�l/�-���Kuyz�Q���Aa���֬g��9�!�8�£��nиU��3�5b}&�u� �1(;"����0�τ�Q+Ć�͖e�R���bk3�g6���:),��h�� ��#u@�p
�-�-�O��Y ��������0[LC��V2c�g�2�,���F��!4�Xp����%Zt���qR���Hdp���5��)|V1���rv,���\9J���b�ίX"E��#���ж����E���aSxֳ�θo��0��a��[E�2�c�9Ugm�v�0
}N���ؘ�Qe�Q����U|NU����5��iѐ���Ң8A�Ah ��:��a���叺/�^�JZ�M��ۥ]�!���0���8���[o�3hT����u��I�=(m;��?�R�W�[V����^cU�3��u�&BY�6����5�''�3^�c����ȹM[��ik-�����hԅlݺU�`Y��λM\�y�^�,�m�7�:�?��#1���u�Ղ�:.���a�!99&��`��:��
�ӡ����30���E�9.��/�R�FM��2]���r�b
zĜ��|=��~�٦aa�V�6���q\��o�յ6��쐍���}y����cp�IK�ҥ9#�)���½;w�~̯<�Ҿ|�J�>j�A���jc.N:���K�3"�@И5k�.�䒰R��w�����ͷ�e�C؊�9}��v�Ç��l8"�퐀?��"�7����4i�	� 8�ň�ٻ���u�C �F�|Ps��$��n�!��U�����8?JB�5���2�����k�9#pq��C^�\���f.��� �s&02�k���{47~`s�Ea��v�Rg{��}����ٽ�F�ݶ����ф6#e:*w���ԆP�*PI&Yq��p�4Kuu56���L������������G�.t��A���^��&ˤ�?z�Ϙ*6FS#�@/�(����FZ�1���'���8E<K��@��e��$Y��?�5��@��2 �s�̀���\[!TA:A%-�/�O��Y ���O�$���x�2 īA$��,�Ǟ+�L�{ �A�ty@�����SՄ��(��<�k$�C�����������a�������#̕�%D���
����s�Ia]�3�
���6�[�m�j��B�h��Ύ��a	/�8�|���w�1��i��V	����TG�A���F
���D�����g�BA�%²F��19�m�w	���t��"�g�c�(
�>��n��l\���{��9�s�1��o�a,Y5Mqo8�;�u�0A����z��N1D�4�4Ї �H��3�OG1i�t�>���ڑ�����L����ζ�σC dCV=Ԁ�"dw����+׆}���b_Tf��MM]b[z
&íw�c �]��C���B��u�&�(��<hE�(m`)̀ ����lظ>��b��ᬷ)�r�C"��&}8�s����[íw�m��y�i{�ۨ�� �ǝw�i"�U�V���k�B�\cY��Y�ؐ�U�4xͯ��~	x<��QX�0��m>�.�ǥ�u�B�A@�5n�޺�l2�*4� �U�/0dwI�1+pU*���ez�jX ��
����O�~Ŋ�V��@P���a��<x$А��@IG:�E9,V�R�ϙ�n������@bߪ�h��YGŚm�h����%��t��F�%CxL�=(�TS�dL��X���ν��L;�߫����_~�1W��֖Ч�61[Gu�!�X�
���	�ػ���l����(�٭���"��Ex>>�g� �s�گ9ߠ�₋.6�pT��:t��z�}Nj������w&
��1a��ZK�W�Lcݦk]�r�i���s�%��O{��E��r=V���t=�ދ�d�9(�/�S�ke���qڛ�C���bz>�����g[F� ]��{����m-}4��a�Ma'�*-V�-����I.Y<^%�S� E^����bZ�H;���̨��x������V��m}��@�_,�߆��Ц��C,���n��a[\"#�W
�!���_��S�v�=֭�S�PU8��_��R�C9��fD�:3kW]� ]AAuP��̕I��'��,��_-�1��#=á��6l�zn�+�6kml3&e��_��QNF�Q��
?�Z��gF����k�n��.���yv�?��bg�sA�f�s-[*rƥ{�����5�KWQ�p�2|�����D�še��PT�kv9�X�r��1E�3���x�s�㘚B���93eSv�(�s�5�u�ݲ{}x�3�v���OX�v�-�b0��/7�A9��.=˜���L���=���G�K��&��.4}Ǩ�.�,�|Ӎ�5(F�Q�	��u�~݆aL�q�ڵ�
�QШV��Z�P+�F*:E��G=�W��;w)ԣB�
��
v�(<'`�qD r� L��@�L��a�ˠ��bպ�apX��耴-8Sl�?�6 �]����Q1OL��v�ut� �c�f\�k����<e�Be����n^�ѓ	5��� �BF�&P�60��uP�I����U �` �O]͍5������^�98[��Q�z� �v���-l�X�0c����I%psXO�4a\FuM+��5�$� �y*�{׬Xv�Mk�Wi��),x���|-����L��W k����;u�}�b�N]�]�kÖ�N���
3�ܹ�jք\6vR����#�[���\��ZM}u8��L=_�K���!o�!+o�vO,a?ƈ�@2��4��7������y�gP�X����!@���<�ﴍ��F�}��Ko$پ�n��J�-�b��D
�`�K��kB=�� ,JI/�h%#��I^V��e���K�r +����d���8�)��}�c���'�,�`I�_�;�o���]�����+yew�p�V���QQ:' �Bg�X��m@y�@-h� ���p��,a�JEY%VA�= ��uon�!Auv5��e�c1wv��١�ѭ �4*ؘ(�Q��!R�zՑ+q���`h���dVYE	�s�Y���{vW�*iք��7�>�{��fEi�?Zl�J&�܎�k��A�g۽���:���g>M���QN���hPԊM�v��Yao��>���8�so�P��mA�
��
�ᘆ到(�>�����l���"�`��g(y�e�͢l.�A�Y��u�a9�uo��4 �bd*��i�V�S�ʕX��jh��0l,Y|5�0d�Q�yR�Z�Oc��VI܋��n�<B�)[jla��b����@��4�,��u떛&�۶��]�1
�+�k8�a�3c����'A�M�V[+��D�u
gM�v�"m���3o�%�\	a�a4  ��M
Z#X�*� ����PK]�rik�J������_�����-��F �MN��
����55օF����RGH��&���1=�d����)�W�{���y����~�u\@��B�C6?4����Z�	�<����_�П��q@SE��!"̝6�l-�O�.:$ا�Ė�j�o�5�"�Ս��X��p��T]��TM�~M8����ߨ�넴V�z� ����
w���֊+�aE6mۨgz��=��	1˹Wjİ5�铮��4Rht�+��Ƭ�9��iY�|�m�����1��`�i���׹�z��x�6=�6�d�pֱZ��B$�� � +0�l�֋%f^�����j��+�k��vG ��}�����a͖���B禬'^��.׭�Q9MI/DԴ��4W5��U�]�	��L��I����V7K`��Y� �~�F���P6^9��/~�K���U�]���#����	Z�`d�"F�=[�Q6[U���Y�e}��%�r�d�L(�_B�&z,Q�M��Y�I�R�7��Ϙ!��S�b��ۙ���К/|8R�Z�9�q])�U�V!?-^V�_ ����'P�0EA�W;Qj� �����/~�j���(^s���a��i��5�R�N���Z�6¨2���T6,�*�/P�����Ĺ���A�\X?��	�
��M�eF��E�[A����'Mx@@�ki�&��7��bB���ł���Y�&IN}hd�v�V�F�#�u�N!��=��� Ŧ���9Sf��i��ک�>��m,��N�����ڲ����fA׆���9���M�Ӱs�{B��ې B�B;��\v����Dͯ��\d�a�&|���R�� ��WJ��ܱs���+6OʹZ�\�p�"��ׯ�)��p�㺗f�j�n��|V3V�����j��3Ч�V������8&V�g�^����9G�i���Ҁ/��>���{����Wz�54	 H�D���z�ă�֛^}Ku�J���Y<�y�@U]���E5�v��T� SY�`��E�i��J����A��Z� �B���̍m��;�B4M��U��e�j$.�}�����Z�V��~���O���kW��O���x8c�&�Ȇ4Lϵa�ڰR�M�"I��l�� @v\u���Vi,���*�u��5�F����ᱣ�h���=LE���	�h�M� �oVL�%)��Р�?�x����ՑB�s�������=�b�
��y��5�X� Ԛ�����5qwu�t]u5��S���TRA󦦱Ul�6{:�u��T�\�ta��k\�Ț!8Z�^�[�ƒ6(6{����36����\G���v��g��b]�q��Ϣ�%z�_܏e�Ա�s:��z���m�JՔs�|;;�Y>zo��^�a�2MU��r�*��#bK j.(�`x`�i�tw'�g��m�i��%�yq0������L ��e�-
ͱ�.���'TPS�@��Ӡ&�,6u���� �2�B�iRvI��r����!k�X����T�`�hn�U�jG� �Q�'ۤ�M�9Mٝwt�#�#��������'Ѥ��*�!�`P\P�*��8�0 @C�1.`ĊWi�g��,�3T��i��eUZ�u]�1$hDN����V)[H�#2C�D�k;V�� 'ÂM�L�0c�uV��6��s�y٭j�//w@�n�ś���Ε�5Nm%��+�}�{��#�Y���}��^��A?Á����� ����j�j^��ҁu�|P���ѪR"$�g �؄�<$���!2�f4wתHz�={�+�"p'�F��Uh���>���Z<���Zjl���,�0���u$LN�0!��i�FK�E�����H1�U���mPsKU�Ѯ()�Z�!~	XA/�m��C(���
0�ku���0q�	�Jr֑�P܏������|�:�w#b�
z�*cm�.	�3�P�!�^�{wޫ�bT���ׯh����_x�����������}��� 힎I�v��J6ќB�~@�a�&��ö<3#��+Վ���k{��(i�������W���N�  ��DZx � ��!�J�����2�؅�/�jk�Ko��󁭻��t���ʧ<%􉄜��l��xJ�~�JH�V\Y/�'�10�}�2Ϭ_���}������l]@��y5���.�&Ⱦ��q���{^R������]K�=Q{�T��?�c���8T����p��r{ ��?n�o��HhG�+�G�F�w����e�e�=S�\��xI����u��U�
�&XXܭ"6��SoV\[dy��'��%- �0'�����E��Iٶɏ_)�P:ESE����QΛz �R�Z#4J�s"7V,UV�uV�Nj����p��<Te��tl+D'�A�oJ����w�)���r����"�%*�{Wv���� ��XT�kgQ$���d��O���f�P"5�k�{9?NG�Z?���a���#�(ݚ��L$��O�]2�`%��AR��G��<f�J��q@׀�H�`�
 lX�I�B'oB�f���tK3����%���~Z�f��)O�n鼰H�^� p`��(���I�nh�-�u�����wT�r8 �L;�J��?������Ph��<){&+�d��#�
�ɆU�,Ҽ�s���b�	˫T�y38.G���b��R>��%��'���4�G�*��3�e�c��T#�����C�!�N��R�	�CS����z(1D���h4j�_�'=S��l�0��4�$n�@�+�5m�='�5���jn� 1o�^����qB��i\'Z<&��I1����m>' W�y �̧?-�ᖻC�j����u�ݖ��K]�k���c�N��j���� �ֽ���?�� ��j�6#T'W�����zF��}�z�/��n��blm��m��
mP�H���p��������~�-��}��![�ɥ�O1G>;55jʣ�r_W���bw4����Ш�$���!��K�XW�֮ߪ5CϦ�%
��>Q��8�M<�܄	%�LJ;	#&��ǵ����JI�C4�lMæ��Xu��R��V�	�]��֎n�.!��-u�@���	;�
�J�"��bI���^�OG��90>2�qΦU?ش��v���%R`rQI��R�0Y�{���M_��ܾYq�6Ux.�]����/��ɟ�"�e��"b�����Y8��[t��P�E%ڝs�T1�!ЊH����P�X+I���Cr�X\��lrH�q��!���ӄ�X�tl2�X��#��1�yL�"��U�J���Y��W�mi�qܞE�NSM� Nfwk��C�2/�F2��- h����G�HX
�E�Q�d;J9D�t�~��$���B�7YNUrB47-*��,�b��NDǮQ=�)�!�v��$~ެ̰�sq�>MM����N r�.�$A�Ϝ*@�XE�ESQ����K��
�9��z�{�w�)�:W��
z��.���µ���v`�I�19	 ֐�8��u�J9E�T��"�;TPAGR���<+��������0����7���z1d��l�սh�Z�B$��'��1):�J�Ep��
͐�gnIcf�`�d�i
jR�ܗ��F�P=lR2�q.�~C����8�3ij�=�����E�悾����� ,�����o0�:���<��݉,l ˓��ނ��M`�*Y뺭O��kա*d�
9�����n���w@�Ds	�Zk�}˄�g�_��5��CK��0��G�cD gR�B�#z_sKUhY�Y��B��W��ZB&�F�&��V��a/���J�̭cS��J	��xm� u<o,+hgh�f�|�ќAW�f�N�ذ^�v�6DX�&��q*��MU�*��-4��ڍ�	(���g,uz(�)FsF��t1����=�7�7�Ċ��k�l{h����2�jb�YI7��_�K���f�M~�탘�T�׼� h�>��s-q��H-1��Es�,�z��mV@�j�XW(U��ÃS?loj���s�n���>��o\�姉�������ǿ���m;�ٴ|͕e5Z��L �E�(y��iaqA�@t.�RMML���"@Z���vr�_�>;s-,4�{f�0Y���J-rr���ɍ[�i-A���-H�2����)�c�v��+~�K�y�`q�9�ݡ�l�53���f��U�f��Dt^Bl�׊8j�c���9���*cD�$�K�[(H�RݏhM�A=kH��^��҉t��#twxի^^������S��E����ƵXO�!6����ƨScV�=:�.:��g�u��0+S�0�����{��������D�K���Kd�XA(�p���Ӻ� b����e`K��Å���t�ւ6
hr�o�ճ��U��9�Њ�6+,R-�S �Ze�ؘV�8%�K'R�g��)Cԫ��ӷl
�}�U��k�PTqL!۱���w��бgWh_}��-6T�G�ޥ�K�X*����@۴'_�,\��a佧ަ���85i@h�`U��(Qv��h�&���7�ڛ������;?�jOBr���E�;����M�F�C{�RQ_el�lEI�j~r݄�d<J
4J�Bo��PDhXl�ب��lP���$��K�Q�����5�=�Lْ#W*oO����y�y�H��F���	�qғ�8���u��H�
0ʔ#���S�1���NN�R��Q!WD�*�sT	
Uu*� ����I�I�C������3I ��}C��������F'�͖
C*D��m8�|�R؂��f3�Q��PU�jE�oC�u�ze�q٫B���m%�U�1)�6miVv���e S=�T����"K��	�I$nl����MIC{4'������HF�%�V	 �ia��Ȅ���c ��S��:i�3�"mh}��#�-q���U�(���`B=�fT�g�E��x`����sc�u�c/��Ӯ|��_=����>�s=岭���c������W��cfr��u-�[��F�@� � vs �a����@��M��M�^DΆ;;����yfi�����C�����)ձ�-�d�@����xUW��3����(�L���0��݇�!4��ò\�?v�4�� ��1���$f�EP�2\�8�Tk��(t�29*~��w�$�	NNN^[?�`���X(��P�A�����B�����w�����Rײ��*Ԗi���n��J��,0l�n�*o�H�M��p�%熿����xs<�����W�/}ɳ�{�����w�9F�/z��Z]�j�()U8B砇�Ha�RR���5�]��%͇X�:	b�vT��������+X���H���K� �H���{��<�R�ݴ����r�aHN��da`% Δ셃�ƦgT��3������g^&��nQ�ot*�/_��+��e��-���b�z��;L�������e�H�=@�FNw��`-�A��8�R�$(�ac��$�U+���k�B�:=+�1+A�c�?=<����L+ž��o�j��� a@���q��Yh6:кh��&�JJE*��{ի҆�zN�Ū���U��V�a�Rl9��%b�F��Ј�B�z1A%
oRJ ���M�YԼ������.����A��x�l%�����%�O}��#�_�R4z�~i��`6��o��+M���i�
�XSY' 0��-S ߦ����-�P.�1�9�f�@O�0jU��,�8e{�T��\- 3(���Bx�����J������|���ZD=bY9����!�]�9��ӞeD�s
��
4�c�
E[�ѓO��4�c�=U3S���JU̚J���3�:F���pkQESc���PD�?=�\���l&YGK�U�R6�I�4�+Y~=r,�A���+�*�BHG����;�ƪ
�3e#�{�?���=�?~�O����<�����/�����>���V��u����qcqiy�АsJ�@(�"�>�yr�qk]�&���܃|P�v(eCXj�I̯'�y�#�9�BVR���N�[�$��ΒF	0d9f,���̑�?޵�K�������[~�Μv'���C v����5c�p,�
�}���6\G�"E�S�e��]��ء��w�#���O�ݥ�|�$_��ځOJ�FOW��� �i�(t�0��s�>K������3���
&�ʲ�	}��xCx��n��a�V}�j��U��M4l �Ke�v�
5��t�eM�+�k|M���u�BG3�N��&��rD
��\5u-v�8hvχ:K�T���ׇo]��p�_�u��n�fk�4%�4G(��x!Ҧn�2�LY�d �}��_�w�T ת�������7�ax�K^������v�Cb����e��)ۨI���Q#6�D�nlb0tv�W�N8C�)1#ԁjV`���!����0�K�/XIfϘ޻R)��׭Rqʃ�����^���W?W"p�ilJ��T�`ɍf��w��$"G�"�3�kc�
շY	b�W0!��ݡ]"�J��L���1?}mh����J��B �q�́tib����Ⱶ7�Vb{䔩��Nh�[!e���J6+誘�0qbfaa���my8,�${�H�^��/���H�ޞ"1.</��-�T�[��9���`=�R�S�Y��=b?�:P,ۗY�:K���ժk׈)�D,=��,�^� ��3�%J�� <�P�-7�d�A����V�}g�*�K@��U��:ZH[�3�?������#���^1�%#��h�l}���!���`�Mճ"F{��۵W{;�n�����<}Ǻ�+ƚ�jg
�`j�thd��Б�u��x륷o������Zժk��Îl�h����tI%V���W���_dd���#��A�&�G�@���Ukg��Xul�o�+�� @K=<�{�+~�����'�����ӷ�{A�J��i>�ř�rP�-�ژU�<���@�B��5[}g��8@��~9SC/�Ң�o�Zp�ny�ߊ�R|ֲ�&��6��9�nN������S<�Bv[��On� =���뷮�1��Q��l,�� �5&@h�� ��rml�7���S{���p��������K_������:>p4��e/��_���Kj���#ݾM��cd���n}T�I�X�(�N�bAtlٻC�f�s���tw�{�zo���}��t"�{�S���,5�����M�W�P�ޘ�12�{�(�?�q�j��L��.9�^9��pM���k���5��}t��{0|���+ܽ�#,_����;���y�+�o>�2}>�׮T�Φ����-pTר�r�%���O�BS�:wk�,�I@c�t�e��F�~�����o}�{��/YX�^[����s^x�ܧ����`'%����d���#*�)=�e�����Fɡ�Aŉ�.k7�v�U���K�^�r�j�	� ,i\���õ?�>l<�B�v�?��Ԧ���<�4�yv��*2��wy[m�����z1����{Ͻ�н��j[�\�Ju�UȞK1��6�}�c�)H�ݩv���K$EQ��|\�d�K-�FFƄ\��&�� Lw�ҟ������ĳ�۰ hD�ٳC+p3��	�W� e�)L*�/@SZ�vb&���bCS�1%oH�!BD��Ӂ�#A�-.�(��Q���E[�9�?�i@��2z�}?��@{C��6���Ѓ�6ǀ���y(a!HA�bk��ƈs�����Ԩi�*�R���\��ª�ƙ�#���ɡk���K>w��gw\v�9��j��W�x����7�������O߹wە�U�6����3M"IK6��^���hc���=�Uy�A������*rTZB`RMcU��*�`��o<�O8��%{��^�����������γ���G&��I��CFTK�ɢ9Xd-ƄOLc�e���2?L0��ϩ����=h �H��j-�P�T�M7�EU��E d`v�H����r�A�[=��x��p �� ���4u�jت�b�l
�pa�қ����
+�|��v�j�g�Q��y������^�!�\�.�;��r寊��	��?K�'o�hz�D�[Z7BNBK��������S.]�/�5M�>��)�Q���}�#����=?<�I��=đ�E1�hj��o5rd�x���o<���;W�(�q��_�!\����Z�p��ݱ-\pچ��J�^�7��p��#�S�F+��څ��g5G�f�^���A���w�X[x�h)LDd��l��غ�#���Ĝ�fmKh^��å}��d	a�F�O�{��Úֲ��n	o矉u��9�{�bx���+��u_h���)W�⎳r�����Ӟ���<Ӵ&�r2���uN�K�s��yW(]%݇2�i!����רΕ����CaŦ5�}o}ChR�>�@���p������a�u�	�^���7�!�s������GՒcm�R] �^�ꗨ��y�O��Ca�ڻ��٤4n�kjL� 9!_!@sF�����`�I �}h�56�,%c,)��K0�*(��ΨH`��ܻ�Sn��s5�T�.��W�iVɊ�4}b+��dJ�A2���Ђ�����ssT*�E�-�+A��K�ä���d�lލ ͮ���vRT���2�f2���:JC�ź⏰}��<�������t^��h=�ةJBj���P�6�?�v|a������v~�U/~�?�����`���u�����#���S�zǵ7������W��h�|�-@+�r�K�Jg���DN�>����B[ ���qs��b��)Lq�*��F���wΖ=�[�p��PNy�i�&?���^�����_Zװ^���5�N�e�K�-H,Ld���n9�](,p�U��C��ve�ŀ�;`�'<B�2(~���"�P�|�˜��`9v��G>��9��O1c�5���O�\�:͋,�.[4�BH�L:1i��'禦�hg��R8��&��Ii3�شY᫆�Û�rL�r�ii�� "�ٰ�4���fhZ;��=�B���%DĈ�gX�R9���_?��bk�@�-�0+A���m��a�G�Z�,�v������?+���M��кБ^a�����ó�����B��~��jG��w^>���T�G�f��?��й�@����
e5�z4��*�������+_	{o�!|���~���7��]a�ڍ��mM�PhQ zv��E�VC$_, �c,�V��B�����g�|�\}G����n�>��+_��/ޯ��2��,���3����?{G�O��^���
{��1`R&�̊u��WVK]cآjҽ݃�O�����fU��6/��������uo�sc�fH>��&��pX�U03T�T���H��W���rI���g�^�����w�W���I�t(��Ya8��"]oB]2:���V6oj�X�j��@����Ⱦ�&Ҥ�Y�M���#q��-�䖨@v�\�	���l��704h�J4?a��q	ݩ9T$FnRmHJ�a7;�J�G�
<jnQ��Q�7��A����S�1m�B�ZS��u�QE�z�}U)HE	��u��!�R�B���e �A�?�@#��A5%��U��R�r+H�͖aR�Չ�!����r�K� ��ځ�/��/��<���m������877!�^}���s��}۾��?�����W��P�M�{��+��u���_�F��z�LmE啥��zq>�\�j��@�h�z�:)�Y0��e���8��R1�.�׈�i�3G7l�r륗�G���z�c/���?��������u��P�ش:�4�r��Ce�^���T�5jk�CK��(؊d�%"4����x�hPh�rJ�؉l��C��y�9L��(������8�]������d1��Rp�5�MƋ�[�U)@��QW'7�jv(ح�e҆)������r2�^���4_xv���1|�s_
��5-mZ����~�V���C�Eg����Ec@�Hv�@�R�9��d;��ü�j�N��fF���i�bYښ�;��D@��h/.U��ȑ��O^��v5�<+\{��f�"��Ғ�>��S�WJ[���I�&&��k��?5%��]�+��T)YBmX�a�|V06�H��ck��a+|é5*xX"',�	�'����c.`����]�#1C�}��-E!�߽K镵���RS�4O��ϐ�'V�t�Y/�K��"8��S���@'�R���v�]�t15n����v����F8c��p� ]�J�ֈ��߹��T���������7���sT�5�?��7Æ5��%/}Q8����WL���px�!��t?ý�]W�.���S4@pB C�X) 6Ť�+�f��5]��U �u���,$jb�N��`d{�����������������	-��հB-?��j_x�c��s~��7��$گ��y�L?��o�Z�4�:������e�O��X����Wÿ}�;��M��J��:�ڀ8Q���ރ0�<Idt����:) co+H����R���=�&�R���x|�a���!CO�C�V�-ٚa��jp;7>|d�}7��ן�/K@i)Y�Z7u�w������~���i�RQg���峉cSS\4��ʰ����z�X ��%�Xq1ץ�5�%T_�ҎQm��W�Yu`Yk��{ʏ�7U�}�_���o���TQV(�)�<��11���G1�^��91��a�J/4z���!=X?ö�H{u^���([�f���\�cD7�H_����lV��W���#s��}�b��!}OE��(ѝ�BI ��_֗�����FJ-� �5,��Mq���}�I�AS�d@!���u�y�I��Y�Il����%�zZq��n�M� ��S�� ��E��0�.�Nm8��aSb�p*M �V��febV�D�pX;2��VP�D_��T��	���� �`Ũ�\����e:����B���H�oQ-�Q�
��+h+ֲ��M�X9s��,lC�i;�h��; �c��E�d"L��I2�>_5a�}/1.x29D��*�?e�����~�]n��Z���?��M1�%��mo���4f��*�z�����Z�P�դ��
�'i�z�=���}���&�J�2��N�uP��uj�Ю�k�u�Pxޯ>9����V�RƔ�A��3�S��x��qr:vk��m�d��jt=:K�M��@�D�d�Uڒ@���(��H�6�g"+B˦����)�<)��WTo����/{�uJKT�l����ܾM�������Nx��_�'K�Q��^��g��3GGC������hoy�o�']~a8���孍�O�������*,[���Ԍi�'toT����jn[Ɯ�uϱ��^�\�MKD;���<E�����+UpN�:�ȴ�_�Y����P��H-;�$P��Ա}����e�7^��������	�4��l;�w���|}wg�	�וh@�z\戴iM��ދ��tCsC��ʯG�2Z�PKkR�Ƿ0�o&� M��TZ<�m~Nu��5#���t�LU5.� <Q��=�-:D|��ҮN�4&����,	��D�������UY��.O
9���M5"��Z[$��ϧ�M)�FF������a�i�3�@|Y��ź�������:/���*1?v��~c��-&�,���c��Bנ�'�)�R�n\Up�
�Y��@yJ��
iy�%P%��J�E�[Wj2ߨ�LM�&�AT�nN��*9��/�<������β�.P���~�$�8{U���������:E��:z�'\t�i��xr���?�.���]7�RCQe")ck@,@��#껥�Sa��}aBmZOo
=�#�y��VZsuX�j�	iv(<�b�����!�0ƢT�kt����͊�������0pxO�~O�j��+p�c�3�x}��KU"�����sW]$2�&n���oSH�����o�|�+_����1��*e�U��BgBJ�D�N��
��ѥ��-ר�K��\�
~LvV=�9k�Fh�E��9፯xv(��K_�O�lԉ��5�ۤ{W����zj���=�r ���<)��T%cx9��N`uN�ŀ�u�91�cbR���y���۸Vۙ 0�*�N�P��(ܥ��9)���~�������d�}��Xs�"<�O�G;��V�ii g��p-/RE,U��e����j�Eg�_��p�~'���.�������/}~��u�B�X��7u���a��A�c�&�ia��,���,]�&���5��� ^܊��w�	qK�}Z�i�&�زT�Hr��@0h5U�Q�9~��_���Z��33~��Yk�>��������ǏN��Ըk�@aXm&um�V.?��+.:��Z�i��e���8�J#(U�E�]ԸjXXk	=�!��]��c�V�]�lY���љr�j��C���8$j
Y�eb���0:z�0�ؙ��E���%�U#g�y�f��v�Ľ�j�PbV
u��3�@
k��=�x��2Y6��f��˳P]�t�����ؖi���b}RA'_�-��E��m^��b *-OKS2��p\N����XTH�J���P�Be�P`pF5Z&�f�Ճ���s�*9�������.����W�vز�p��'�[�.\q�����P+��yn��I�R-�9��Ë^��p�Ĺ4�,x��g>��Y!���J��]L�\/����u�>d!��=����+����S�|�z2u�.v�j�9L���fi�:�W������<=��տ�ᣟEu�T�*�}9��B�2sEL��g��۴L�������F�Gì�R[����/�M��� �&����Z��OSGt�G�~�O�nTO29ezDU�v�W׹=��c��5k��K?�9O�T}��U��oڨ"��l:<�O]~I��ݲߐ�q�T� Z"�u֨��a�lQ;	F���U���O����7�Is}<��^����	�x�3��V�Ԥu��c�X;'�w�Yᆛn4�UӠZ:�}TF�Buu���I�D��i���U#���c�i��<&;6r8[�,��hH8���j��>$�3�;���/c������"����(|�k���P֊����@�\
�JCF����>��de:mE�Q���d��^ce�V-%�@f>Br�� ����db		��7�m��&�|N��"��֍91S0@V�ܞcv;�A�n]dU�았c��2sMdYJI֖�p���G/:s�w�ҋ=���c.;��w~���޽��%�EEm4��� ��fKssg}]Aij��H�@AKq��:�׆ʦ�*k�gkj�TA��/�^__=��ֺ�P�a:V9|���+�zm��� ��r_��:�	J��I;i����fd^Y�j��H��qzIb�x2��-zY8 ���\L�1L��"ĂZX/�q��9i,���߳xG�X� ��¥6L��3Rd��RS�0D�e�z�����/�~�^1
5U�{���a���hWh@�jU�E���\EMK�~������-��ȩ�y�
��1_�}�=�{w�{�_�W�.�<<�����G���uk%�}ax���rd�O������?�����������i��i���֨�29���%�	�� �t�}��36�7���w�o�0!�J�ݏ)3��r��ן�k�z�w�R��kTQ m�M�cs���������~�	Լ��oox�)%ۦz���o}�����Mi��¯��s����*�o\6m����o}o���[�*�*}���5/��ҹ%hWqD�ղ�5����#��'�#v+�uŪ��'>�I9e��+<R#v�4R��G�7���p�B<o{���.:;4()�C���}%|�_ ��(��������+@��p�c.�"��fX�b�U�P=�Ç�����û�����������f��w�&Ӕ£z����JV�#Z}�F����ׁC���j�F�11B	�������R��Gm�:�K�\����|�����ד��87\#���g_iMc�}����];Á��l�B�z�+��c����k�K+�*��z���$Q���дl��Fa1<�^�o�.zؘ�獴���@&(��F�'W�¨ .�iJ���H&��f���6��6��
���%�?�v�*��ѳ�I�qb|lv���г��巜���a%������?{Ƕ=�zj
�mi�g~b|�\eH�ͯG�2Z���ӍfbJ[.�?* 6Ewg�?�/d-ZY��4='�ش�m��T��vw�ۍq�А�aZh�u�R��X @I� Z�s�vr���s����i�`vX�-x�ύY%�>�=\P��q��t<�Sd��n�ɝ6?�5�=c%~o���YϺ�B�rk�x���FAԺ�d��@CtM��M�x��_��K8[���(�Bw��51���v�h�CGyRn�!T������{{�����B*^XQg���9	W5�^r�.�,|��__���TO�'�/[.�"��z�5��f�@�ֳΑ�����7��@E�ո����O�2��/��Cuk���g�-|���}�ƥFm�����װҬ��()����f��C�?a��K���/;��� �؃��1�
+��j��榛n�ÁЮ����ub+����w�{��^ۤ�}(|�[����&ց�-b�zU�X B�c۶{�U�4�z�/�N[;������תN�5WY��J�`j��À����WT{K��	��v�����ưf��[K�^�a��Χ;l�z���(V���e�[n�5����^��ɑ�*��ad�/���1<U֟y^��W��z��ޫ_.{Dz9Mx�<����QG�X��	w�)�TL�OM�A��A[�A�Rޟ�7�ĳ+?�,,�9�~����\�r;�3��_$|�o	�y�;�Y�~t���[��Q6؜�	��7����>�#ij���G�}����\����*��y_�k������� �Z�*����Z*�@;ڕ��xf�g}�.R���H� �����Ș/��� �_�|��A�H��^�O�o���Os�z�����g�����i텖����usϷ����#`�($������=(�7�i� h�#^_Y6�P]=֧�j�4����?;6��C4�B��K`�|dx����a�����j�5��,K �̞��)���Śth-T�}�Α�d8�q�\�`� cb`}e�(�u<��[w�R�?�;��$/ X�^��7�C�p�m�*��Oz��X?C�nBl�?�]-�ֳ��S�J�+`��&g	E�-��fw��h�-�L�/-9*��D�U��$Ǒ�_���:
v�����W8�P۴v���[׋��Bp#�1O��TEW�;]Yd�]3����&�+U��5�\�i�P��ມu���u��LZ�~U��g>Y����W]���:.��:��]�*�)LԤ�mZ��� ���kC��c�����H h(	4 �%�2��q�{��Δ���c��l��F���.�ތ���OA6Y�v��:��ڿ?��O>��9�P�@�r����YL�@�!������8�f;e�0-ب�Ya��Ȝ�T��C�����}Bb�~b���J�g+ugH@\������9��Q�#TӤ��B{:�*��CJ��;��3'�9!���	4�gk�ig���������m�jR�����������ܘ�}��5�	���i.��>�*Ǥ��0��I��'�M����\`K��z�)�b"h�2.�U�bm����b�fҥ�{���~�b{���5�ݰ�ĭ�Y��|�[
�Մ���{�%gn�����}�>e�	$��	�o:csht�
�\mz
'��5F3��ఴ@�J��Hi�8BN�a�_�!a_�"��6ր��=v|��+�'B�V�Й^��jc3�(V�.Ku�`KƫѵL�ό�jm�XV���"Pnjh����?:��hlvV�
���R"�o��U�w���89�#�j��/�2Z��{�����]�����OL��JX"fw��>�ǎuu������*�7B��19��ʡ��f%r��j��,
���*U�&������B��y����|�Co���K���Vq���L�$�0k�
�-�u݇W��wa2�����r��?^�� �|wy@�tG4t�b�u\�����3�SU��2`9:w�����Mz9��)P����b9�֊P�{FbVB��Q��ڵk����b��u�	��Q����я	�VA�M�k�-�	��7�7ܭ�����7�R�z5-j�9-�M�&^���_�e�!Ԫ���Aiu����0�~i?2)@7��u�)lԶA�a��l=���2S��{z-�R�h���S�mB�U�]��B= ���IP�]&��q���A�]��E��� p�a�:����B741%ӬG"�Ze�+���5b��S�eU�VH7T+�U�̪�e�Y�������F]v�槴�5T�h�
�]r�a��X�\v��Om����@Wݭ���-��ebT�x 
�~d(��e�~�A�"x0?��Ig���-m��B�5�},��W����!�z���[nW�_}x�^~빏����^��pݏo��f�AuuJ�Ƶ�ĭ��Wx�߿6|�K熧]����k���G��_c����pDU�ר��<������0����0���b�0C44�`:�ɂ���d���'2�_f�4�b���9�$���ª�MP�G���*+����Rgmъb�j-��*��..���d�b=Uך�����q���;���?_� h��1�4������̩u3�h��f�;g�O�`�4��%����������-k�X�)pg�yZ_�p��5|R�Ҥ���#���"���3I��=�~��,�'���v1�J:��?�Z#'��������I/�O6�e�&�FJ;M��=��`�F0�X"w�)��	 �杄	[_D�����|X��!��<�rR���c�G ��bu(�V.&�pwo���l}��tPՋ��qf觞���5ᴆ�IZ�T���%�ՙ���������Ђq,�c?,��m��L���c
����*^8"�  @��ƃ"��_,!D�Ǜʌ�9�^����ɏ�����r��-�s��A��cM�����l�J/�I�\Lsa���9$D:&@j"~9�r�O?�YӤ���@)IP&��/a���u���7�.���ŧ�'���4/�J� [��L���8�#��dr�r0 ��T�����b�?�"�m���T'�m���Z���+Tʡ)|熛��2�KNZ���*���r����½;�)��U�\�	��R��w���6�����m�����Vv�&1�0Q ��U��s��	6&����#,)��n�$�oP~�!�O��7��jZW�=�m�NC�R=�|�aD�Ҳ͔V��A����!�z:�yŒ=�*BMq
5%��in(����B���,�A�M=>;W������kZ�������C��8;3�y��ܾ�ˊz�x�>��xO���O�v�UujJ���!&����`!'[,^Ls&hx������S�=M�T��ɿ[����N�����µ�x�RRi�V'I�9+�e�͌=�E��3��F
���Gl1�p' ��8������c�135M�LYO�	�=hƨ�;*q0L�+�[[�=9Us&if�>�H4TXq����F)�sb>*q,mT�8%�M㚀��Z��ċ"r�`�y'�{aX�JoCe컶�-�3�j�
� tt߈��F+��a_B�T}!�����k&gJ���՘7ԥ����Ұ�`}�K_R��!�[e��{���+V�2�5OX�"L��]*�^��XE]~J΍끅�0�gO�J���{kT'��#��^�����C���7@�N�k��Z�cǔq'mz)��FCECU���Y�~���4mj���e�m��}Ki�-a�g ��;Ø�$���y����6��������-�F����Z���wu��I[5��,7
r��o�jV۫4���	���H�5�����Zs��\�7_��,n�E��L��m�aЫ�F@�Q��x��lC����y�٠c=}�Uu%��UE���T�@��U�$�O?��p,����� h��FNB��Ւ)��sF���]yþ�g_�o����羽�TJʟ�u�ۗ����D�Ji��/�~�ŗ�g��O����S/8E���I;���D�H{عO���N~�I���JN�����{9ձy�-�ѩP��0z}c�B�\�'����Y5�S\{Z��w�Ƨ��O,-�M�9�� Jhd(#�D� �D�-䆎I�!����U6�K�ȸu�:oڪ�̣c�ڦT�FO��Ƌ]:@�m �z-�e)����z���CZ��/��ԣf
p�3�c�G�"����f/@�gU��
/�*n�h7�K��JúH��c�Qա�\Sbp VU
CK�V�l2����8��a�� 3�E�sF�� ��S�j��_St��(5���EF�!��Zi�Д���j�s\�ڦ~��견�e�9�"��T�Iu��yƔv^By�$BX��c���kv�p�A��O'3�ㄝե~�y��b�1�_�6T�,7 ��$z��n�i���l�O�~e�U�5�Q�a�ƇB�ŲM����^���	��1/��Q��^,��� o����7|s�QN_O~��F����c�R�Ê&�����ޡ1��{y���utb��S_�޲���ͭ�i
�������U��|����t�0?X$�������+2��j�Wh1�~Ȅ�9���xު��g�d���_qW����v���y��5]���+˦�"쾽����%�"��؍��8EQ������ ����-��z��!�Ŕ�)��@wF�A��94�{KXQ�;�d��|�4���D��X�v�iG뇏 r��Oz2[�:��5.�����c�|o�MD-��-���� �S�@A��I~�u+.@Ct:%%ʞ�f\�WZhKT�b��nl����6�6��BK�r2���8�H8B>˸9rD=�v�:1M�UDGp�b�h��`�UPś{�5,d�����(�g�ki.�P��:T��>[� F*���%P�U�RU����(@���g(�c���|�ۤ�V1���C�C-,X���je��@H{%��q����' կ^Z��ej)�>�ܰY��2���J�6*D�^�T�A���r+�i�<[��T��
f$@m!��ܙ�J�����d�J(iA����տO_G����&��2�(���B5�J5��B��b���T��A��zp���ҿHMdQeD�ٰʘhr���fƟ֕A�+�ܘS�������σE���_Z7��
@�,��3YI )�*�ٹ�ؿ-��F����i�w��G�O�+������+!N�-�A�k���#�-q��r��xV��5<�����X�W�����?�_}��A�AK~]s��o�뾗�T�n*��.�⏓4-�8��R[N6�"Rж�Y2�RKo���=��uq+�T15>\̈$�b��Fqg7��pqX+��	h��%��x�@N;2��]C{X��E�� ����ig`�b�0�\�#7*��J�5?.,̮�Y|��}\/� �[rZ�C>�צ�p�t�^���ߌC*^�
F�B����� X!�kTA�2�H��:pM�ƪ9[m}�R�@�tw2�`pRaJ�pd���Q1t�g�3Tn����tn/iOĖ�M|�Z�H��s<�u�b�J�6��� ��8~��p<g�$p����i��븴1@�C1D�
� )�<o��V�a6�}E��;��V���YZ�G��5.Qp��r�J��r0zV�*+�3)��E�_'���
A���F5���J��lJ����?��Q+e�����r���!��l1^�emK��2��:�J-0��>�k�R6yo�C��R�q��&�gzt����W�a����xhs6!�rZ�gT�V$}��q��B�\.�Jy3����\HC�:�3mVb�.=���� �������E������JuU�3ݧ��$�[(�*��M����+����S��Cݶm��C=��O��t+9�X� uX���Ɇ�ꮆB�Úв�?���$��⟓�������DeY�$�4��b5�bv��-a��3��9�������7���]�e�ڻ�\s�ͯ8�?�����eԤAӀob���!ʴ�܂C?yN;�ű�����Ď?��ݹz���!Z6�}�69�t]���y����
5,_�w�:pց�V�-�
]��\Ӕ �|Hm�v]j��;֟�}���Y�'Υ���]k��|8H�
��~v0�},�g��y��hg���iG@9���M�wB�pjF��ӵ���~;yמ �b����n�B�;��tTa�RlK-�*�8�EH�ȗ�V,@B��¿x�Ƅ�V�/�e�8;'GSQ�����2�o�H:�)\F�M�=��<�7����n-,�{F[�Yo0�:!Qv���>I�!0X�z��dz5��U�M�I�Ka.�Dr�֞B܁k͘��;���a,QdM�AHs|�\3���X,,�Wu�|-�.S;�+f2Y�7����;e�%�MFk�ߌ��|�ar=_��B�+��T�̘=Ӎ�c,��`���){�o���F�0h鹧����ʶ�zN۹������=������{�145�Ue�L�%@�Ҩ�ǌ���������r��zY k��8حu���E3ݣE��M3څV�V��בɀJ��[ղa�����򚳮��ES]�����_���_��\�����K��x��׮PCL�+��gFxh~��>1y�b��>'�P'�5�o���'̲(�~���Y[f����CA'����̼��y^W��b���{4��k�`,�1U�D� �	 �uk��t��g!�>]�O��"0IvJ��9���^i�.FE�LG���X̒�p*骑Up~�0��'�K�!ZoDw�?�N��M/�e�gEd ��S[l�yh׶p��lҌY�Z��b�B�@��V#��j�n[;増�� :���.lLX}'}���(7�V�3���^�Z3{1�gi���EGz�v�@� ô�ƗIS5)V�O�g���x!'��<��&�h�QUSzLN�z�Emw��	�`��h�Q��a�k�u�����J����y�9�����|�,}:eFZF �$��6�`1���,;^6>���2��g(6�5���1d-<sșw\[�>��X՟��q��8�L��æ�ã�&�/.)k��~��;���3�n�rP~�ׁљ��~��'޳�೫�V��S�ƼBe�T@�ácG�7/�o�M�3\z����2Z������X��G���ytY��9��,�J�],]�K�J�^|���g�5U���������M��SG�u�����54�M55��ssǏw�t�l���笽{�?������w�l@vgM���H���h/,;)��Ӓ{�4go��W�����ŋvJ�~(L�bg��XŬ���s<�hXp�񓛵�t��Y��9�3ӑD���ȼ������o�-Td�X����T,E�8N��� �A�t�'j~ _�1�/c�����7{*�Y��Tw�.���5���޿�� Qr�&D��*�}�0^z�J��UV���5c�5�k�� �]+���X'�������?k M�VvarıכP��Ҳ����R�{
eΉ���9����P ���P��k?Q~�F���ʂ�E��ήcV!��vu�`y�4:z��A/Ay0N{�c���I{����%���Wl� �;$�n�FJ��r�%���TBB�SXbY�X��DB:�$����}~ߞO�aΙ3sf�+E�D.����^U���b�h0j�E�K}�H�dW~��Dz)� V��&�W�i�%W���D	X�����8�j'����n5Or���W��em=�l��#HD�����`��Z§�)cs����L4Ϳ�>�33zݝ�F�z�?z��^q��'��YX9��~�<�+���g��+����g-�7�?n5�յj���ZV�z���&4n	(e�.�/f46�P���;������:Z+�`�O��}���5j�a��͍���8��c�,)����=����yj��2Z�6�٫��	�S,�I��N#�`���?�Cc�k޷���c
��%5�?�)#Qy6�y%��1��ʼ��+�]�|hE���s��07r̀�v:��v�Z��Y�~M�{c�X����Q%�}��T��o�$rrs�L#"�<B�49Y[Sa�[a�J{�̾��tܖ?j�B�����v��w�4WLb���-B�ؠ��Z���8[B��7�+�W)y�O♇vE�?=x��u�SQ���wLS�����ڥ|��kK��C25���1��V�x�}$�>>��&�Y��� ���>%�t�䩪�����Bz���W?/�.U7c5�y�ꁶ����^*�Ӱ ��'�R��8%�ت`D�A4�c���jQ W)�l6V���O�=|J3mbH��J������n��}U<>����y�W��)����6�2ʃ'���K�d�'��y��y�iH��-�J�e�^K���DK���[��v����m�mAJ�jb�\����Wb�_*z�8/�/:#�C��J�>f����e��"Ҿ��4LKy��?��i���I���l�9!�q��u/�g�}����x�7�I&����w�KKjƟɴ�A��_�Ǒd?-B��BT�W�0�b�s���\=S���2dh��"�?c�ޓ���w�Ŋ�u�7k��1>�+�=�0�w�x)�g~`��Ӊ^3h@ ��#�­C(ͭN����E����p@�V�҂/�����d%�|x���Qՠ;�M��V���ff���1Nǆϐ	��L��mEѮ�}�#����s2�񿞲���X8����h�"*l��UcݽN�T~���ZwدS�柤H+���4<�4ܶ%xG�V�ݙ�9k���>�0ҙ�\���B�pS8?��3Vh��*�G&,iL���C��!��Ɉªҙ�|H���K���t�74���*�b�{2��$�&��e����[ǳ�1G�8ô9�� ϔ0F���]9��q"l��ʍ�mZ��ԥ�ta��C��3��1r����*T�Ÿ�T��3��ۮW�q�Ue��J*@�L��u@a���?�?�/�rj���y����i{>�/ڮ���q~_۠�'b칀|�-��:��v��-&��ۂ�-�'��R�4U�u�U�Y�݈�SАbI2m.��)~B3~��̰v��f~���0}��in3l��C8^�Ig����j ��
���`���7x�d��&NHdR9p��C}J'<U��4�_�O�ŴO�)����"���y�4j�P���3B="�;^�����Z}��-�г���t9�j*�@6P5$�lkrx ��e0ԡe�v0���.ݶ.��8}�&�>�k(�~u�03�=��h����e>w�����_�������L�>�8�q������k�F�G�]je/w�u���W��:����]�S�>�:�;��՝L�^\�m��'�"��E��c��Ɋ�D����UH�h���k��FGKw����$8w0޷� K��n�f���wR�*����!���M�\��o��Y�+y�=C���}����l<g�F�p2"�k )s(���ɠ'��?G����I6��O�7��*֠�3�bo����rJm����@kr ��M�-���9����jW�`��āT����.�d��UD ���Ф*�_�uW���9�3����ΒP����4�%���/7Љ���Zܤ.��C�Wk�[����TC|˥���:�6�њc�͍]����u#\c�$,��ت_�ϸ��r�����;���*������ ���cs�U�[Y1%oO1�4�� U�5n�6΄A ���Q�^�f����;U4)�y݁�\@#c�B�8�z$�H���:F6BX����#3]�/�m�A����Z{�M~j¥�|g7�߼�qqfC`[N6��}]�f_��}�$��g�\Q��n�T�d	9����&�����6z�b�V�_l���fJ���E	��ӑ9d����l���M�s�;�|���9���MY;4�-]Uo|��t���@���<��ĭr�op-�_4���1����-�ű1P
�5 ��(�\�j�W�n�>��������ۅ�eJ���2�����[cg�_��
�L^n?<�xY���� ���{�ۍb�k .�>MZ�����\:]��z:�X�%�B~fwX�
:\6���M~���m��H�������suC2j!�����`������vf�6��+��b�ū�=%J�ˑ�2DDR�����|5�㸐^Y|x��VܟL���~�&/�ˋi�����@� گ�{����K�
Vh��bDG��Ƥ�<�H��%G<*:i�Ax�0L�K��̊��_����x59�������N�?1�Z��1�$��M���{�P�x���E����RGJ��;����*{�M��lh,�ᙅA����`��)����c���1lD9q�'�+1F)�Lou$|Ø�	(s�N.�_���,�v������oh�MPT_�W
C� �oUǭ�k�Jڤ翵�ɾ�ƫ!���F��G���Dsهsc��J��Ĭ�F�!֫�L��?��Xvw�z��d�$2J�s�#4�Mc�˸g���H1�����=U��|���Ϩ�g��g��]f��=����5�!�f�FD��"M��&��_�������)�E��%��G�RO^���7p}ǽ���*���w�A���\ķr��G�Z�u�<kz3@�TjS�<�K��}�Zj��v��^�2H�Y�"٪hg��n�|�&I��^�OF������$dd���,S(q�W�f0�f����Ӗ���U����9�6Iw4vW>`�c*J�f_�g��{&��t_���]z��q���|����/��Fv�٘�r�v��9�ڄ��S8��-����y�*VV�+��f�6ᕮ��M�l��	JB�t,|Et,��Lu���$�&�}-�r��M��6 P=�G�ԏ��X]��^U��	��c�+�C!P�r��Zs�ċ!��̫ -�9�}��-�m�[�PT:cM�z��UnV%��Vs�j\$06��V�M��}��Ķ%��!�5������<
��K	�c7t������������̤�ͫ(����''�T� _P����\Ca��Y�,N�*jU�L4{��Du�Yw�'����|y�o;�`�?�,,��_ʌ�RHWb�',���֢g��=����2������34���p��'�s����F��²�'>y�ա��f�7���,.��B�����0�]�zM@��It�w�iM�u�l2ι۹����WM{H�S��Ÿɹ"��[0-׊7;}�9*|q
��y����	�|����ͤ,41��P~��z���il_�њ?u�Q���ף�9��5׼' �%p1�\��`t�����%�W���D����H���Vs#���2����dJ]���޸j{6�Y֟�ӱ�38�N�J�,�$���٩5���q5�������5 9d�I�Z~A}�m�<7v^=&���F�f-���(kMuS�O��>�yW�Eb�i��ix��W��kL�*�$`�x�ko����V��㴑����l�J�"
�X�����9B�����{o��;���b�m0��s16���+5[K��r��]�0�Y�/h,����I�q�H��-[5l_iQ;C5�����2��o/�_	`>�'o;e���|k KX����[KiB%�/���V^qX>O@.W���A~"�x� �k�4"]����N�$\������Y���<;f���^)�vh?�OΙ�0�((�O����&���*�H�=��Nw�}F�_��%���İJ�,��шw۬|3���g.�/g`9(��&&���sB��OK�q��G�k�U$A�-����ь��X�Ix�V=�cNq!���� /���gt���E0���]Ll�k���AO �R&'MyvG�Y��������ӅnR:97�o:�\�+7J�d����.���������%ϩ���sf�ԗ/��Ņ]����>I%N5z;�p��g�^#�"����dl4�C�2���[]6?Ȑ�/M"��;���!����ǉ�']hK-&@��d�V�Zt��x_K\��lΊ�%��'��m���o���8�K%��<���]���O΃��O�ϯa:�Dr����О�� ��3.�u��R��}j���	t
��^�gSD���||����c�Pi ��-E������MDF������)#Щ��'��e�ֻ3E�K�o{~� 敜TU��]�?����&<��1��g����NW%<g5��.4J��rx eX��pB̮�cl,{2j�}�6��q�b�'��n�a��� �Hc��� ��"y��>I�(�=4,i����>�>��;�&^��B�I�]����IKt �:B-�b�Q�F�@�\�Nm^�3�2�v�\��ⲵ�r�bY��L���"Ĉbc��1���a�0�J�iP��[��Y52q��
"	~��F�1fNk��v~lI�)Vc���^�~G�����3�*ԝ���&B��3���O��}��-�����"W���Ե��Sxc�d�X��X?J�my[������L���@,�_�V����QZ�Ca�n<�EM�A���1�p�k�f��� {�h*/uٲ-���v�����Y�㷫�	���ʟ������J)�s(�v1��1�8��}G�7�cs<ǎW���u4����9CC��ᓷFji��$�i	D^T�o�mx�}��٦7�-���99#�ΤN��z5�Y�D����4�E~�F�獓S������۩�#F
��.��;v�:ԓW=H7��Yç�Z���|�l���4�l�a;2���m3��tcɗ 5��I��HHE(S���eγY���Z����ji��RV�m�ZezY\��k$� �];�#z-����!!%���_���<��g4=U���<���E����;�D+F-~[��t4��u�b�0\��amַ̀���tS�2TJ�U�uehٵ�(�Kj�J'g�vlQ�}]��U�#��x��N��d,��G>�y̡(��㰞p ��4���!�2��AA������(kp2��	���ک�е�
�X��F�6Ū�_"M�
�91!�h�)�Q�hb��ph��6 !!~�Go�i��p�/�@����>�A�n�=�u:�8��pK�0W�4�n�K����q`e	wW�;��?ET�c���q���6��a,d�.CZq�/tX� ��ϼ�%J������O�Kͷ��/�Wx] j��,�MUjB���ZtV� �SLo o��11�P����fO�D6���h�i�3�b��I'	f'f���ct���������R�������N��6/O\\<nI<q����&�Xh%G�グ��z7ҁYyS<���hbcE�jû�[)i�ގ�+tusc��4	

j�+�GP��@x��a��|��eֆ)Х[oS�k~��;0j?�T�c��iy�u����xe;{��j?Z���B�-='�ɟ�!󷓯�\��ke�
er�������:յ�ňm���p� �0���i�#ڱ6��6qO�����(�X�5���C{	�n��)V���A+�Wɛ6��!D�)�u)��Y�E��/�	҉)�������a2������V�Id���5zvV:�c�.��ݵ���@��27����XK�&$m���_��/�Z�����?����[����,sN�ti�J%�OSUO�^���� PK   �cW<�� � /   images/d3b60164-5006-402c-a3a5-273a0eda4daa.png��[T_��I)��锎�[�sQ�kh�F��[z�!鐎���a�����_�繯γϋ}��������MKC	�_EY^���ſ7۹�U((�U�rrZ*rrZ�lQP|s�3��t�)CN��p
�q:U\Q�"&�X��^3��b��[�}��:�����J!=�ڬ��a�>�n��u�9���~���,�3~3.~�8����C!c�dR�*G��Q��
]h�}�BB}��J�沊��D�/�Z�	��A8W�=?=v��H�B���N����8c��A�j'n�ؤiy�!�	�	�~|(UB`�i�R@�M����D� 
?��wC�4�½�֡�quVqqP{�����^�I 8��E��c�Em1s���ݐ۪M��=Olݮ�$sg��Ơ�&��)�O~WyiP'�Ec�,��4�	/.�:H�%(SbͲv%ʨ���b�}s��M���cJ���Q�~����/[{m܀���hp&	��~HᾨnN.���o��z7�'�/!WmO1��?� ���Y���~��z>���}�b��w]bQ��:׮bV!ԽśF'�>�a��h�e5&�us��yX�bP�>�y~TF%�`p��lcgnǹF����3�n�.*G��0�[�7�:��r��A�JE��W�����f�{Č�y#�z�1M�|���E��/Q�u���O��3xC��Pi���-�GC��ƻi}ѥ�0de�F�����|{�o)j�#Ͷ��������+�����Fg�6߭�F)��>IhfuF'K�J�?q�`3HRe�Ĳ�)��E���,g���+jN�X�J�8�0��:鷏;���_ ��E����;��]�hآ/OH��!w��or7�@l�������u4A8��(1��W��1�
�?S�tfT�p*h����
ŴZ��g�I�cK
~�q4���F��l����L�G��)�j���{�Z`�ȗ�J�%%i���?dV�|M�I��~o�4�I1ҝem^� ���M�M���L@�y�;a�MD=�y�2fk��M���U���մ5�$�S�2p��un�
�	&
~�'BϬ��CX�UF�HuAzAɎ�pE���]^��/廪�z�	=�Z��[�{n�a���$�T�`�G<�(	0�Z�S�5��b-�wd���Q�y:Ji?ٻ2y�z�Mv�46}6A���ZB�8x��u�%�r~Ѫ�YZ�zt^�M1�)��b����tq􇴌Kݵvb�=�s*�U�+����j1g�1���&oA���Ab.�{S��W��4�uYY?M�H�؛��_�X���OQ�~�D�7q(v��U���?Ʌ �~/�!A�LO�#p�|��r��:ۍ͚T5���&_"_�P=P1�O���w4��r�^���+�H+6�'q�͛
��ĞP��Hf��)�ƮwR~|��c�ʲ�}�	���E\�#��?���}I�O������Wӗ�/���>���������������'Kk�����mH�W�y���իd���Α�?G	�s9�y���%�N���m��&i�l&3>i<����@LW��Ӯ$G=�2�|�j�|���������w��RգƄMY�=�Ä́�z�aG�G&ǫ��ǕG�"Z4���"ލ�db'�G_
EǼM�3�W���Ƈ�u�}�����;t��6�6������w����"��q�2�����k<��˜��j �
Ś�I����X�,���_V��:�s�� �,�t�j�@E �@�L�Cd/P�
e��Ui�i>�?�>���s�20s��0^`��v�n\@�`���2�=�����륌�SIs�gG��ٟ��l$�$JE�"�儣 ��Gpｸ�]`������(�I&
�8_�R�U�qg������Uԫ������ԏb��|)l��5�t~���3�CL�d�B�j8gL�CϮ�v:Hxq�p�H�g�~���.�	}V����g�u��Wd��#�*t*�*��)�,�%��i�/������t�����O����z���
����bS�K@��n�(���"e�	���,AN���Or�x�����6������e�����r�i����it���{ ��:129r;���vv�`��O��;W�4$�9� ���jsF�b6c�b���U�sͰ���3�G!�����v6�8V�?�"5,�������,O]L��o�5Oot�5m�s>.n�u�o���ܼ�U���F
M��#!�Gګc�-�|8kWa���b��-�4���y���}*+�}�NYWϭJ-���W۩+�*�*�N)�OI�J����x���~�/��zEBj*���A�Aw�g��^�^^XM�.eQp[Dx�.}���Z���<EE�b7y��~�.Oz|��w�W�F��9-��jV~I���1����֌�T�e�S��G��.��B�2w��o����bGÛ��{_�Y����3�g�G�����</��C�S���#t���_��/����{���5�۱����\ua3�F�g��`%|���t��~����"�����-�d����J���a�$����K�(p>��\������v΃%@�wJ��@$X;/�pF�%8�a2�l7֏	T�H  ,��K0�T���8��X�x����q��l��joN�Kf9}���zWvw��2W�0��R����:<5!L�Z�l�llH�҄���'��0��}�BIA�Fe�>*e��z���p����#��r����O��RA,$cD�q��:���� �o�^��`+L���;�&5��Y��A�]����S�-m�)D��:j�x�����"/��kq܉�*������'��DY�����2?ȴ�0��Qk�k���H�h�l�+`kq��燅0���`�UV�%Q���ܕ{�ܱ�����s���N�����VW j����g�b�򙴈˰�0���C��}鬴��̳n���8l���rz���Hl�O��NGZ��r�[.U�M�k����r����%�{��;��} U�S�7qƱ���c�Z��D��:Ub�6ʌ�b�M.S]�~Pe:s�RR�:Kw~����b9��5�����u��ke���r�?�d"㞼� >H�y�K�Z���p�o��w%����Ծ�׏[�����%����7�Sґ�{P�lmPM��U���3��f�ɾf2��~�)87�L��mZ���v��Q��Av����9�7JY��|��/��omV��Br���`�&�ZJ/�Y�kAJ1l����G�7wYO$^C��ޫ����+l�D� ���5y�;��%�ԛ�%԰�)'�1��=�}hjXgp�F�eH�wP��A��&?�z5�,5O@f�����P�� Y��\���-��c�7��Tz)�@t�'�떩�������#������䵷�J�c����� D-/Z����Σ�qk�F��ʠ<��y,�a���z��l���\�����Χ�Ώ�ص�]���eח�ח��{`&���8w2�D�x;���KdUJ�H�oȦۗ���c�0��U���@�q:#vì���I�y�a����������?��?S�jZ�IvQo|.R#�Pj��ytO�׼BLE������4)"��t-���Yg�>����l�t*���qX?8;x:r|���v�Z��;_���^`!�z8��A��x�D�X�`?>.�د�k�_�;�|����l"�fi�]�*|�(y�jS�=�=.��'q�ci��Kk�Ĉ��M0�wZ���X�p�(��(�4�6��g�D�&�!{�.�uD]S�w��i׫���	�M�Ǹ�|���7����Z���a��b���������ɒ�RB�]��?|�7ˍk�vϵ�O�KO�rj���2��SYuLu����б��'���ʔ.���{ݩr&ڿ���A��*�ff2���A��M�H��z�\^!w�z�8�������P��	�uL��v�2c���n"�i�:�2ֹn$�%�q���<�i��'=h�E��ۊ�,$�=kW�L�SR�,��g̭�;�y�D�.�)7��)�+�7���9"��[G��/8f(��0�s��U��y\�s����@�*��vC���Q�ŝ^��O�!�+~�?3`��/��K���"��1޽!�g�`�WF�Jk�>��؊�.����B1j�?���~�b���G{�"V���#�1�Tц��X~Mg�z��,}�l�do��.tx��\�V���y�޼E���X[+�Q��87ꔢ��!�"���ƞ�l�݅M#�090���fS3�UsRC��?9J�����CuOy#�\j 6��h� �ܵ��[���y��-��Q��Zn�il�#?tl���U��qO�����Y95Ec���i�͔�z�ʵ�<��{�Z�������U6iK��sf�#ZC�Z�vC��mq����B�9�_�&]�� �k�g�I�z��f�(CRޭ����L]E��ٖM���ػ�h�[�mS�m�<<:���@H:Kf��3���
9_��!Z�A�?N'����~a����"Ղt����	b��G�g}�P`=�Ď։]�8�9�F�ϿA��&ly?��+�b9�U�-fi�w����_B�)��YO�t�-U�\��B{�m��_;�)oD�-�9
�
��H���j`$uŧ�T���K�_��+�%bT�Ǝ����JH��;�]"�kIq�E�?�F�~$hqu���ᆨ���;d���;��b�M9�U�%c�+arCA�D�S!�	����� �x�����X��AiZ���x8���-e!�zͫvl�g�*���)dN�z-�����5˲«,�S8�r{��S���x��Fú�k�'��{[�]O
!�g�kIC�@?7<4t%[d�Y>&߱^�5	��nz�EE��*dk���������n�r��g��˴��[�(�{���;�捻
I+��:s@=���Ҷ�?�v�`N �Z$����ǽ��V��H��{/z_�ډ���I���j��P��S����Ǿ�,v[!���_�6��6�?�z��S�8�{�u��
�.uv�����]Ep�����!ʹ`�F��$p�V@��:�LU0;�����j���A�N���l��	����u�vFl/���=�V��8�\vT
�����E�k������+ϯe����.	iB�Sx�՟t�EPB�w��,�UPvw������X..E���
S֋{�z�)�3�fU&�.��~�~�=�q�p��|,�W)ֆ���WZ�2gf��C]��Ɇ&w�%�Mm]�Ѥ��M���n�87��B��Z<X$?�-�@����>ԥ'�Wgq����W���+;�&��Z��$L&�M�v��t�4����>mq7B!%c�끦��,Rvh:\�ܤ.��d\#i��{v���p��H>в��"��Ǩ��p|ܴnn��et�B�h�̞΄FAtn��4���n�b�[�ߤ����ǘ¼��|�:F�+�>2�H�j?��/x-p���Q7���pO/I#�P'�4��h��V�d��{�xg
�Ee�gU����w }��n��(H7�+�e���H����E(S�%M."�k��F�Ip�P�p�q%a�M���U'��^OD}"�ϧX�T$�8@L�,�%����\�c�2������iM}l"���5�i��O:�d���k�G\�;
*��ӿ�D'�h�0b��j1�>A��@W­���j�W��픠7Km�=�|P��Շ_>����]>=��]�7���r���:�˩��%lx�Q�AT�*:C��&������*���u��њ��LRơ��H�X�bQ�Ni�������P����/�>�����9}��j�L0�a2�?��c�NG(;�u��+m��';<�|z�淨_�`��Հ�Bw[��rF0vN����3k�9]Ge�~g"��a���6l�t{T�6�`CKk�_*c�U"�����[C�j�x((f���>�������_.h3d��$��\���Z��*�e�>�\��Cپ<�(��]�ޏ����;Wu;Ќ�5�J��w��������T�vLH�<�J��Y/�C��.Cܣ��AJ:VV���}�_b+J2'ɆI#fX�mB�E�A
B����B���Yj�m˄�L|,D���4�a-��d��N�_�Ňi$j;p���с��rhg	��`�5*֔�vuP}܏�o�}��B���@U�VVƷ��4���6d�%��Nfvn\�oR��(6*��nU�ʠ��D��k�T`#]]�Jj(�����Dt��`+��˱�%��~<n{����y��j]-�y�-E��<m���wY-��)�:s�{��;�L%ի�$.t0���? t@w"�v�p��NM��V��t��JLst�h�\�5�hfԧ���O�%
��C��8�����T ��Μ�g�Kw8��x���,��x�V��s�G�=�[D�G�EN[��� �qM����th�>��y��������ah�`�HHJK�(֛F�l'N<��%��re(x���eA�ez�9økUb��5S�޶N��.Mvǉy�&a��e��˝O�/mr���3Q��M����ڨ܆8�_z 嵃g���/7��~���cd��f���3�\�F�I7�5�Ic�����#kr���;Ҝ} ����!���_}g��� _2��f+������ 
��&U�/l2V5ဋ��s�`{q��N�����@��u���kBs<{��2g4�d���tH�M�U@W**6�j#�؅;���Fv�B��z�ճ�
N����믧��o��ZF�o�FՈ�Ѩ��l��TdO��c�l�{�5�DO�>[�%g�""�%x� \�DAY#s�-�%d��Cl��/B�>�L�2go/�u��3,A-�Q �(��:6��<~t--�C�!�W�ÿ�]�Y�(>Xr3d9o	�<��ur��<��_�� �
�W���=|���������Y�&$Ϝ�u8��b델Ri�;6=�]����=#mѳ��C�,>���	��%���2Ͳ���y�{�jV��֢ONkVV☭�/B�ڋ�7��p� �VS��1w��d�~�)Kp�?�&��c".N���4)WY{oM��n<����1��k\1&,�x=9�u*��x�Ȋs�I�2( @&�}	g��w����Ӳm���)6�p�IoGn��+[��Qv�i�S��QC۩6Z���Qm��Ǡ�>��j��Dp�X�S-K�_w�g�&�l���W}w�1ԻX��SXm4-�ģ�t&�;����;1�	�;��*v{ٮ2��S�(A�]"y3�sq�D�x���u4Z /���Ǆ���2KW�c8Ȉ�~G�澲x۽(����;�;b7��"�ƓgS���L���D���Yu.D�o��OH̳o�r*����ֻ]��U(��k�6�[Ǐz��	���$��{��?�,1���(/G4繖��ю��xnh�yL�<�� �[�8=���j5�OJYGd�ٮ��������f/�!�5��,_^J��U����Iv%��:�E�F�+[f��Q�M��or�9�Qb�s�2�T2�T���խ�w~%�/�{#���Z���0��J�����Jo~O[׺�E�;JB?�P*����	�U���:49҄tk�G�rb%�껰��S#2�l�_�����ǴV�<:l�c�}��W2����i�H�x[H^��Z��%%ܤG��G�?��Mb �K\�+�����Q�rȠQ�lX� �>����)%k:~.jb�Avu�3���HS�b�i�Ig4`��r�44��#��#L���O��H8'C+��H_.�u��x���"Hc~=YE����d�X��,PZ�IDWS6+sGkߪ� �à/��Wx�,�0]?e7����SD���JJ����:�X��UIQ�jC�DI�\ٯ�z�[�_ݪX{��
R.�%�h.
Pӓ��`vd�y���᪀c2ιYv5ʃ�bM�k܈v�BZNwe�ٴ�Ns�w9�������b�㑽�hd:L*M���K�?q���-4iI����=Kf�֕#Ԃ�5G2����K�!�IP�����t�_Hz�d̏l
����rqY����hF6*�;�_��A[מ\�-t�����6:&�W�6��v͇#p��	a\�[E��X�����k=1�ƇЅ�`]�ȉok��F�!hJ���n����7�k>�w����#�<[g�^�]s�HFO�e�՚�%�;Q\�S��)Č��QAM��Pi;���Mí[�YWU�@��c����OP�10x%w�ll��𧁸�ebq�|�G���Nږa��K-T���~��P�����y���%��凥��b���E�h"m"p3x�b縷�PX������P�Ή�S��l?M�_i�-#k�/o<	��a���8�� ~�J�8iPAP uZ$}�Zl�X��Ǧ�Mj��� ͍�f��FOZ��$0Mp��K��FO�Aus�n��8f�,��C��j&C�/�on��>�wcc�[&R{:��0��`�ĉpS�a���'MI��%�z�g<-߆#��昘(<3��{���0�˅�u�������N�og���:�z�x�=�3^�n�/�r�Öު>��/N�?�NJ�0���b�<��kn,y;f��=$�%�ۀ^ٲxՎw �|��|��X��1������� a�x�I���O���Λ��<���i�p��X&Ik�@ǰ5�؄�;Zh�X�>�^ w�d��Iz�،�M/���=g��H�V��Ɯ�ٟ�K�#,�l�����?+��_���)���$p�q�Оɏ9'��(�1P+�~�Q�nF���|��q�3ԓ��N�*,Yh-��Vs'Ylsbz�;$� ���G�q����|$e�7��0�+���N��尳cL��%O`�U�#�8F��-{=��F��r���I����:~a��UL!�$-��̩�L-	PF�ߦc�\�ʁ�	,?H�tӜr`Ч���
u���B#�ۻ (�m} ��F�#G��kًr�#�e�ޙh
a݌�בǽ@�&�O�U�y
�O^JW����N��M(�oR�.�&D�6�K����\f����a>&���1tNq��b��Жǀ��'�H�6���y��OS8T8�<6^7���1�P	{���EjB�S��?�i8!^Xpl����@�+�,>r*bC��z���_�)2]e�y������O�B'�e?CQ/�9�֦4���00\��^Z7�Ò�8���̙�l�(�@�_�`��/O����e6^(ɜ�w��ѮD�J#^�Xe}"���.������]�u/)��)+���Z��R��<0�r>wp���A~����sx���ߍ�Kco�v��6r�]~L�o�M���*��z~��m��x�/�T��~�<U}� g{D8t�o&�=��y$�嵹�t�^~ܘ}�qw���&)�@�OD�Am�1k�z��M+��_\;r���s��$�&z�q�[Xon,j��0?P5�^����@�S{�����z�^�2G.�y�X����� �����Uw�=d7�i�yq��ݜل���Kw���${e��W��v�f������N��]<��u��m_�$�Kk���c�8���7[Iv���\�qѱڧ�Z����v�o(5A��Dt�)�Ԩ߻L�S�B�~��L L���U1�"�{֋�{�?K7��P~�'����堳�d�jld�F$��qM�ʢ����������v#����(U[���uڡc�n�)�X�;�����B2��R��>���P�ɗ��3�֌޼yK���>�ĄN#�j��j�����GN������a=�2��+�(�{�E��R�������4.\s+`���ԭ�Љ l�]*�FE�o�0�WC�\F�>��«e��#]0rf��d_j�m���'L�����������?��m���CL ���a�������KZ�Uv %��M��+���WĖOsV=�)NZ@9����+��Ʒɤɀ�����8����Kbŭ���n�V�* #�6�-@��ФF��٤FNv�h�tUfQh����L�b崜��-nG�{dmaSDIB6>��o��^{�?.���K�g	>?���w}��|�NoN�k4�'i���_�^��E+�%���`����#�\���+��wn�D������^h�K��I���v3]�H5�03���'%�z_�]�D�KR�sRZ�;�y�M�/��ϺZەSrMR~�Q"}'��ދ�w�G݉��T�87qɖ��yN0�D�Ge�^�����k 6[?}Ύ�<��y��&��o��� ��k�x���#מ~��I(�;�R`���9��u�T�~A�!N�^�r6>��=�wo��?l���9�R���=L��}�&&#�t�| ~:�m	�o�x'<�gq��_��s�>��a�����饄x]뽎��:�7G�BGU^�N%1Y��"�@QS���#�{���6~�+Jl�C���� W��gn���w`v���[a?�i?����~d���IrPCs���=;
�w��#-�TY��_����<�d�U�6�Tn�:j��.��ʹ߫d/`5���Xߩ�D����جv��BU����;���S��A�V5�u-��x���A�����cψ8�U��vk�PN|��3h�j%οi)'y�ٳ�x���\� �r��ȡ~�Zȹ��Vw��7� Q��b��k���4��@IJ�Th��L�u1BLA$g��>�,]Mɦ��৽��gx�c�n�3�6{+Q*H!PWpGϯd7��Zϧ{i�3�e��$��bb�*1��I���}��j�݀�H�;�����/WI�F!�������u��B�o��R�����_�Z"d���uH�/�XC��Q�vK��f��p�6JV��Ό�`�פht��R��0�S=�p��Ӏ�{!�nn�������-��[�^�9�^{�W�Ų���"��?+��t�E{d�b������0N�i��H�/u��#+-����XR�~�o���u���ZX�Y$�QX!���7�&=��&:#�H2Da���3ܫ*�ƣC�c�4����t)\1;��n	�e[�[}��x�\� ��r,pj��f����T�r8�H�4^�����H+8}����'�	n�ݴ�FU�N�vs���\�D������a�O�`W(�Z�M�6�ۥ�_Wm��F�Y)=���<��i�	��`�q黽Ma�Ӭ ������|�b�?�%�Py�ZV1<w�H$�T͚�����.��f��B�K-�5�xU�O����>��m ��2%�ӓ��Ԣ'e�tC���ٲ�.�����4LH�Bb��;&�ːßK.C���~C�
%���i���zW��w3o���������v_z�=��/���]:&���\p,�9�F+��V��	�����2�M�nz�|�����n�� gJ�4G�V�����I�xkHN�G~��W��)Տz}I��ɽѕ���KN� �LW/2V>a�dɛ��Ǡ4��!리��ۭΗ*IV��6a(V�.1MÙS�+���ȱ��������[#˪�S�Q(8�,�i���w�ln��}7y7�g���D���UD֞Ğ��ʉwK����H�O��	[K�_�Q�~�M�.��]N(�-�5��O #��M6l��J�=�SX�
�H��(2�&4����(k]{�	W^����/{�MU��9���[ĩ9F�>���.;/��]��*�$}���a�9T\$�$���r�x���@�W4r�c�	�
ϧ���k�n����A�#G@��*�Ws*0������R�u�+6ʲ�F"G��t�R6�����g�ܐNGL�/b_o��ƿp�;�g��"a��]�:���栀b9�� �q�,�<Ի~L���ϩ5A�?��
��4��U6ܮ>?��P�wo5Dw�fK�@h�8c?<b�|��&~e�o��������$"�j�'J���X��K�b�*��1(�̶���Y��D�����JkX��ɗD=�C<$9P`��Nchq�i�:��sW�e�{G�}��O�[�o~v���'w%���t���AΚ%��6	�%~�i0T���2k�.ka�X	�cxq�pF�aЁ(�oG����{,�XSX�]:�.�F��0|�X�uR����B
[k�Qj'j��[�0V;r���֐+��gei���7�X&\�W5��I�B����&�����h�E�bոv�676�f&��:,Xe�I����@;�@�D�0�qE�����$&�A���'|.z�rzR����H+rSY��^��;�0��Y�c�E
�["90{����e껂Fgkv�!'��͊�<�Y|�Tynq�6_�8���m�3��~$dM����d����ޚ����8�k�edr��l�l��muX�i�5�	���1Qu��� ���(ْ���Q����r� ���om�&���~��n�B��fj8�ݔU,����� �:�~K5��ص5��H�Gx�������	Y�L�@ x�#����E�c���Pl��$~���D�sxE�X
��� ��z�P���m�=t�W��B$ܑ��y�up�ɋp�u4��`|e�8���i��8S�=u�h�쫰�%/������*�Ox��{:��+�@�'`��T�7��u�6���x�������ՓI����5�����;��"*�+]�7�e�y �c[k���p����ޅiB�o6J�>gD�n���u3#y8S�y�ax8��2`+�}[|��^�˚��R�Q3g3�Vn�@V��3���������<�onW��^ة^R����G]6�@0���ǜ�����W�^��D�+p1��̫G>����XuC���6xs;�6���z>*F��::���p�¡�cŢ��K������
�@�[T�.
���di"qZ����5�"���IO<��/V�m�sn⸧��R�W���,lnһ(��t ����M����f6}r_�Y9�����:<��.n����~9�3g��������e��t�A��!Z��5�Iڗĕ�|���/;K�P�0z�[����n+}~�4d<���C���z�hB��O���J�B_]����Ai��E�e]T~i/��b���~`�����ã��V�	_"t-�)q�P�x����$Ft�J�+}�|����Pn{\.��W�$�W��;�4O�r�)@�P��@�
��p��|�XO�f�pi⭪��ߜ��D��V��W"���~y-����1D�-��c��
5��*X������rR	�a:{⦞߮D6�	X�Ҥv���C���V�5iO���|4�T�G�Oa
����1��Q�T�ϯI:9%��{�靚>���'�6Ղ�[vO��s��+5xq�e��m��t�G�3�\���F}N���V�%cn��8m�M�;��$�Yӓ ����?S't8��}5~8[�`����[�\"vH�D��Q�����Gq�2w��$Kx�oN#Y����o�HC�M�;)��p��w����(�6�Ux D����%��C����w��9���@H�=\#Ue�c��ܔ\
C�+�l�`գ�x���v��o�=V���N�U�܇*%�A�=����Uv�V�ޝ�^�N��'i/}��b��U���r�3g�>�Ub�HXM�Κ[:��+/��/��{864�T�ܣ����-����q�e��Um�E�ĭ����/M�ʗ�y�E�8���ӗu�y�M��E��g����o7�`2 _�ԭ�����}���� �j��=0�kR%��p��~�^�Ŷ�!F���ƽ� ��	���?{�;�u�;���}Q��,�q6��������ٮ��Q>������n�&ȁҌ�go#�*�gwP�`F}��UI)���e?mE�)Tbﶏ�Ԭ���E���v�t�cs�k=����!�2-*�J�A��yy�NNO2qI�"��	{�Z����r�Ȅ�P����G\�\���܅-O���Ki��=l���!/uLJ�Q�����A\�-L	�q�^��_��(�@�����$s}����k00d���&��~���O��a�i�~4�Φ*q>��P2�׳���9� ҃�~2�"]�AE�����;y�d�~Qg��N�����H��W�J#�F<��� ��l��d�6�䛛+:�z1����ϻ;���5���!*���}��(Ŭ�|��J�N�����L��b���b�������$&��	�~��s�EwcGw�Ue|"��/�7g2��ٳȡ�yb�lR�1�*9I�H=R�«���*ǳ�ǽj<P�t��{��f��L�Pԣ��2
�������Ep�@��_�@��ɉ��h��S?+�-���XZ1��.��u?�˥E�_��w�;���9<LR8�<�_bzd�di�r�?{�1-�ͣ��r|��U�e���Q'6�jn�}�2}m�f�`,��#��mk�ξ�v�̶[�i�\�/?�o~{���P��d�{4�Ԓ����x5w��B�����S`�+��탧�vI�?��P�ʼ�n�Mĝ���w��LJ�I�����9/���Zܰj�9u�{:{�*D�U��/��q܊����o�#�N�����a��pޛyT�����⻳��כ�p8���A���cGPyJ��Y�r�_��V�ӡ%�5��ՎE�Vz1����c��Q��M�����J�J�,�>hќyV��=�!e��hi6
���s�d�k���MBR���\<�A�jd�ŏ��.�X�1O�P�%b��M+`o;�g��������JH�YQY�%� ^	Dr9�&�r�h�a��f~l>�<���Z1�.�??] ��0�1�E'J��P��*�<[�J� 6��A#b��,��S�
yS�3-"a�I�"��BB��^_7�I�c�6W�|�I�G�0ǎ�#�-N��uM`�r�q#���T�K7��EߧP�b̹��%n��<=G��Į*�*��Q�a0I�H92+��O�A.�Y���IZX���E��=��_;%H^/�8���6���E�N�(t����Ƽ9$X�7V� a��	᩸6�J"�+SƤ�or�}N{��f�8��bɸ-g�s��9�t�>�qz=���2���u�o�^ 
�n� ���,���b'������;l����Ba��u���BX�eC6����3һ�;��]�μ�@R� �tT�̺��|q��^�>`�R�X�o��d��l_�*�b���#�=d*�W��gbe"������r�^�ڞ�ϑ�$�K�w��Rg�RuK���o}��Љ�������q�;�+p�n5�;c�O^b���r�k�7�"�����e�����s��5z����T����X-0~G�i�3����L���&kz�g�b	VtN!úoh6F�i�xYJi�����i������,j�n�7��a?�t����5{xx��Բ47I����'���%����=�����:���	��۴�?����e��8��F!U��9�G�=f�oZ��,qť�Z�̎΢�A�JZ��"@�F�P�}q,��.�K�{*vN��7�eI^�C9ѥ���X*�a�-j��w���#�q��e����&��@�\>�a�x��;��L��=��zڒ:1�5A/�`�����Ks�RPK�?�BRՓ���A7
��P3�	�q1�{f��tl�o�z�/�k3�3��Z������S����rN��XQTx�'_@�(1Rn�$���WB�ɑ)�CosJ����e�nE6��#<�yW����5����k[J�~7����ߡdb���=�$1_���k��`�>#��nI�u�?�`+�W��8P�<��R��䘬���Ǵj�rS�	�����il3�����/C��:�=0oX��p���3w��p���8 @��)�}(�V� G-tZ��S�I��%߱����V��y�{���+L_w�IW��с�W����!��F0V5�vc��v���`�?8������uĤds<�c���� �g�#L'Ô=�;�g�4��v��N��E(�[�1��Ŗn�v��$K�ہ������I�w�L�8e~=xu�B�W=l;FJK̈́'8w�	m�o&�����bgv��i�����B�]K�H�,\m�bR5�v��L�)����M�X6H@,g!���� �s*�3'�0����P���8�4����Uzp=�O&l^Ӊ��4�Pd�.`��e����vѐD̤�
��������e9%��ӹc*UHp�g����#��ϩJ�a�Z�������R��+sq���9�'ӧ�~����W��ke^?3:��1��Q�o=����-��u1'�3X������[ſ]\擷<���ZI$��ò��IW���F)�I�c�h�����)� ���.��A$Fw3j�FbĨ~�?���}�{�s��sg��@Kh"�JNx|�Ͳ �)Y��v =(�+)&{�;��Iwijp>r��J����]���37�A�9�,j`$2����}��{�!�r�ʝ��=G?7��T�� �=�\�����eև�wY煉س���+�_�[��f8$�f�@�^���*�-r:�& t�ol�<������GO,�>�L(��fD��,vn*?Ǚ/ �P�95��1�Y�>����36�!n5�.�nF����`C$�b��P����B�Q@ȨʅҖ́B6�*�$�[e0r�w?��4��&�Ju�T
`-�q�M�a�N|Yl�j����2�E�s��|u.�+��>������=��b%]?��
��N7���H|�W�q)g�3x��2J�HL�30��_)�����z���~�r�`����j��a����heX�3�aU�Ը�n���l�N�ǌ�>=l*��)�EC��ɻ
����i/g��7�x�c��g.��gi������ˌ�Ī*m�[��Ja*�evhʹ]mю������Te�ٛ�F����>s&��@`L���@��4;75�[�>�?l��^���\�My�=tӘ ���-�S.�����0T��H#�qՙ�$��E��d�K���)#[�F�c�6�vs�GQی0V(~WY��x�� �
���߂{&&�č<l/{95G�d��әA,�Iǽv0��#�hg����V_�_��n�U��"��]��_s ��]��yX������=�N2Y�S��Ax�D`6���0�!�Ų"V�/]�&�Pc���ˬ�qO_e}�th�U�9��E׊�診�s�/�p��,�ݟ%��w��b�ֻ���]������=��v,B��*�o !���M�Ő��y۹�+�H|����\��UH�N� D�JB����K-�pH�!Kpb��\�E���=q-�^(��S颅M���k��N�I����n�v��n�W��s ��hc��3������ǥf%���R
9����Y~�U� 1��+	��T"GC?�_>�k��1������Q�C&t!�(�s���i�m�q'_��~c�{�]癏�T��P\!���~>�!�0���X+����9�G��n��4��ݥΊ��4��<�L�O��GS�e��l��3G �K#ԃT^��<��uS��0;��
}��t���S��@��>�F��G��k}K���8��_X��L��`t.(K��d�d3j����.C?,��kz@�aw'˧�s��s���a����Q�kf�_��wU.���Hn֥,���9���	@�D���S�(�?�z�la1V@W F@f�e��@Ǣ{�����sc���>��ު$����>-Ag(��WP������=��+_'���L+���s�(~,?�ݖ�R.P�y����.7��}e��``�Ql�"��%�EeB���Pq����?%���f���>.��Nl���V��]oږZ?�5���a��E������}evZ$�Zgz,{-��៷��9Ԋ�v4}�ż+Q|�u��źT6�T�a�o����e�S����qtJw�@�C%W��f��G?��z����_�7@����(�Hd��g�`�W/�|�݌��`��Q�y*�"�.������W��fx+�\͂�Ia"��Ac�zV(���eS.?�9�C_IB~@qRI�w=�~#��C=��e�Vt���T���o�AN�M0�I�5����g�{���uV�a%�)�����lL$����N�V����}Ӿe7��6
�7��辛FŇ?�zj�TX-���ZsU��2�V쳐�S�h=��ћ�>GWG�xO�޽ت{�b�"Tݯ��ھ�����t��ށ�К�qMV5����B����4Iװ��<�򋧟	=U�|���wM�e��� ��H�m�eH@X���M�qӼҩ��u1
�K6�􋅱�(�K�H��|F,U nI�}�k�����a�Ր)����)1��7�K�����������K\N�U7V�E���ԙ_�����ֿ<��:�*�f��֛}GG���'�E����u�A��\d���@|�;Q��ӵ��Iq���Kצ��Q1����O�q�'�(���XS��-xqE��X�s�.�-�@;w� ��y�$�w��a�=�a)�?^ɹa�Ĝ�(�sb��HU��kg�C��M�'t��pv��%��Kn���P�W2��ϸ��\c'^l&,'~;�����PK�<E~> A;*����>a���8ʦw�s���f����o�@#�a�0��7����x��Ӭ�*j��_�.#� L�rR�Q}�DMC��k�$���6z��R�������N��\�^
`�D>\��0y�f�Z|��I�wB�p���'�����)A2�l5f��4�.�2�u���n��2��(F����q�Υ���Lv�ZeLw��Y�x�Y�_<6�N���1�k����9�W`�شb��ndt��hL���G�������15�]�"ů�9^M4�l�>?�*UDp��+��Y.��+P�P���x[���g��:�������/UMwD� �׼2JK��
^�����˧���~��g^voG�W��9hd~��&Q(��+2����=��Y�,qM��6R�Ά7��Z3怍||q�@��j�Zڊ.�����ލ1sHXs� +\�̺<����=�\3�1�V	ʜ���1�4q��)w#��no
G��|��G];L2v@�L���L4�@�#������d�����
������M��j֥3t��at�����x�/���Uc�b�������O��Z|Vr'�w(d��oӀ�L8=`�6��Ts�W���ޫ�t��+�~E�Q5c��a"�˶:]�XF�)���C�R�^Y���M���f�V�O4Ӹ��M&�e+X:��E8��Hp��5b���'�ʲ�?��×da�'��t*L���;p{�!����e�Y����X3���0 |��K�<*[|��H�����^y���#b"��:�y.ws��^�}&2�O(�ͪ�����O�d-�R���k!;�Ȁuj=�e>�* ���A%X��0��fG��xaJo�3k{db��� �ow"��m؎�Ծ���/zR�C����9�2���N������2z��ʗ����آ;���������rB�x!�B�f���X��P��Z�����Z��{Xѩ�be��ӱ��@�.H�����Dy�^�~s�TnGڗ�Gv����HV|YQ,�U5LaD��=�-�Ksd�V4j�����:@��PN� ��4��w'cnQ�"�OUc�N�j������,(fKa.�aW��qT]�:ꥇgz(�md�� ]�#�=�LMcW���D� Ūn�A�K�%�@��oц� ��(sj�8������Nm0����h96�j�����8�yR�k������z4e�%�a���N�j?w��/��C��v}S�,��I�mZ�k�^�G��!N)B�R�+�Q�-��|�����Q�CN�!���&���z�ߎs��D��A4�a�bTI�6AZ����C�gF�G:m����G�)��[�sA|PYӫ]��V�������naw��%W�l��K��[�;(2KԆ2I��?��g�;#8n�)E���w�Ҏ�������a`=����}4��J�pR���>p]�*�*���6-��ʕ��m;аc����0�N{��I���Ey��R��l����9|�/H�/E�%q�9�}v��:5#q$�sG�#|�+z��T�OcĦ%��d����'�O�� I�X[+�.�t{ og^qD�ak�S]�8
��������0	�D:0����מA�M��M�WY�Ue�1��!u 1��a(���e�I��lw�曳Z���7���D�����P�Y	�ã�[�JM�����t��u-:Пi����&qLh���>|zeL��iǢp#c�
J��i@v&c� N�9#���H:�HL]vה����p+�,�(��Y���(�)�.
�\��4����(�s�����<�<};t9f%�g��a �%��BM���$���	�i�������p �p���,N�����c�3\B"Z~��g�n2��e	�}��=, .�\B��xxÓ�kRKG2s�5�GAFf�O=L��Fr3�i]��#���$(Zq; k��
�芈�-�'&ʿX ��_�7��f
�,[�'B����-ZpIZ1d��͙ʥ7�3)��P�W��z���[��!���W�e�b��c�A�I�ٴ�6X*+^�(����4@����%Mո����4��_��z_��hI��ZK�Z�#	�5s{D�DO_��`��MĮik�2�6~'���o�aG��@�2�`,y��F��L�B*�0���l����c,�MhH�
�5Ku	V{l�rRE�q��eʹ�txەaD�S��/�>�l�*�i,�wM(�
��ĵ�mO9��Qk��m%��/�����fN��}h���4��#���ѯN�b�6'sTy���`:�`/	?�\T�&�&���dL2�U���W�g���.
���;w�m�< �߷��S9�͖�	��	.�v$�*{4��Ϲ<�Rb��ӬQ:�p����%,��CnS�6C0��3<5��󟪛�A���>���|��F��n�q�O�(_�o�"�9A��w�|K�*��Ǵ�����Ob��A�Mʝ8�F���k|Nx��2A]y��zCĕ5Z6�E�T�Ma���*p�i�Z�3ஆ�a�[�%�A!��3/i�yT���jo�wIEP`���F��M2������ٺ�w"��L;Qm��/Z�Y�E��y��,fߍ�z����.��L���o��8M�듵�>��e�+��f�h2�H���h.GP=o���?�`�
9jy�T5@�#�����2 1^.3����IB#�p�4vt��i�IF�s`("G,�����Ȣ|�/��n1(�w�@`YPn^{���I�<ҕ��]0s���c��ߧgK��!o�T�M��*4"V���E 9���/�MT�MY�x�c)w���&R4��[���m�e.衠���D0f,K=W������n�����_g� AV��A3{І��&�ي0�Z���.;}��a˻�zj�ݬ' ���_���m��z�#&������}�p�J�쀑��P�݂�I���}��z���)9f`T�"_�%��Q�7����Hc+SB^�!��W�aF=+�v���$��s��T�ss`�-[_X��dlz��\�iѸy�^�C�7>��{�
�%.~��6�����Ywk�m��ι����@�_9���u�U?7ou;�hn��<�Ĳi1E�/�_n�Q�:+�<��nkaL�ɭ�l���RCƩ|���y]��,,� ��c� lI�;���բ�/<���[h�>��ن�<F����J��ۧ����vB��|�Y᭲_h@b�w�m�&.@F��B+��G�嵇�҉��U�|����0Wm�\��C���|@2����s��Xey��5ȵA�����i��$#I}�@6�OxD�HJ�GVոk']���{�ݞg�]\�B��+?X�2�������Ԟ�������6=t��*�$>�|4�	�2��-
�*�E	�#����1~@eʪ��,�O��lc t�{_@�@#}�W���8��߉�G�0��053�$�缚�v
�"!o��Sa�H�A"[g(W����Z�Iw"Y!'��Ku&!��Q��#�Z�
��yԮz7�%%x܍Е����h?�[;�I=30�L�:��Г9�V��z-�����Ke%N���h��na�k�ů��G�|�^Ԟ*��i�-��� /�d��m(�ߕ��� ?�L��×?O�:��
[�aF���N0�������ti'!f!�klz}"��%�rp�6��B���L���7a)6e���X �$�.B盉�E�^J1�O�(=�4�[&A<�<B\�1V{~L��?	���5MZ���Z�a;�WVׄgЛF���S3B�U��q~�c1������6��`��|->IȆ�oYe:�(��G�p�<)R�M��F�6�f�\�(���S�A�-͵��F��Y!NP������� �2���?�ںk�(��h��:�e�qP"0?S�52T��X|^����2�tZ���0�a&kl�x
by!Z��7�U%־	o9}��v)?��R9}Q��N���T�t����������$"�J�P5�P+�>���ά�|Z`0���KM�|��;��
��݉�Pjmˍ�Z�I:dq�x� �H�H���jiŒ7�҉�m�!�7.�Ǉdg�?\G��`}	�e-��A�2���\ְ�F�ߝ���vJ�+C�ϓ�ȸ+�
yI�
���ը�]�):�Z���+}��3����N�#uڭ2�?��� }	'�4��A��s�����B�[��=/h?^�y)՟*�`�b��0^�p{�ޗ����I�0Nӵ���r�N;��x^��rգ%&�`��7ȯ�$Ng��N�Lr���L�J�ϔD8���Ս��0�BkV�Jz<���d��gX��2M	��v�̻�6���
q�;���Û��QM�.��*Zz���@�i��^��Q��jBzY7��HJ���J@D��H��'�*���ƫ(P�v�t��g�������'�O^��g�d���+c9�Ҏw����X�!���V����N�U�6������,_�S.@l�??Z�ru��f.�#�W��X����2@���A�$��-I�*c��6�R�n���<ڔV��/��qm	p�����,į�ۂ�kf�Gآ���+�[N��GEb�������tha�y�r�6���	L(�%r�ϲ�-��nz>�2�����X��#�CZ�62b�l���P?]-8�u�Y9���|�
lm��H��j-��3��o!��}�3�>��%�}Ͻ��Xu��3��E��1���ٛ���|�v[�Q�(��Ac�J�~��� �Ѩk�8�_�����o����8��k����䤿�R�"Y�'u�v��<��i s�di�0b�[Ҟ�c�����"&*�c�m�����7�c|" �_�3LU3G�ɒ]ߙ�v�_��\tz�=�*a��a���7�
 e.I*ӵ�N�{0`�Y�Lc�h��];Jbԣ�����L�`��N��9+z�`&��������Mf0���$��ꔔF�Z7w���e[x�PI6��O�%6�`6l��x�Y�ߐ�nKV8s��'3� ��AP��4mwhu��
���|2��)H��$F�U�M�;N	�����ܱĝ���_�����QN�'�J�d�BI�ɉ��*���h���h�4SeC����z���A+�	�������s�^&�%�k6U��~i�oA��P�}�vb�}iNtw�	qB9������rt����d6�"�Gƞ�~{.y���\e�*l�{�A�) k�WD�أ�L|�v�)��g�7����>��K�q�����i��@���Ŀ�pt�*��@��T���ͥT�o�����ߤX"t^?(B�Va��*��y�D�*�k�L3Fv8T����l�M��I���e"���ϗ,�����>�q-N9�-�֕�1���5e�v��R}�q���g���_K��x�U�I�K��1{AOX��FU����^\��`�j�z{;3�k k��ɨ`J������x�Qn�ԇ�Ѡ�(̨Ď./ Z�Ա�����J�9��>JD!��("��G㷮_P���I0E>B-1>�vf*u�-��Ixu��\�x�2��{�ō��ȗ�Q��:b��i��l�/=�n�ӫ�ׂ
�3ܦ3e~	�u��/T����Y>�\�)��it;�<���!�/�e9T9�� ��<����?Bg�鱾{�E��/�8�o�i��d^)�f��F|~[���E.U�S���ƒ%/�ub�h�Ma��b,׺��4c�~�P!ѣ�r�.ٙ:�m�h��7��fS��|5��+�m�"b��u�ñ8�9�Bh�w�j$�F�e.߯+�ov=`�E��v=��}[���&E�.�wR�}�ck�`aH8N�����W��l��3�~2�6ū��a ��:�GI�B/��N���A��#d������Py�m�(���*W�`�]�b �}C�_��P6���Y��ǈ�r:;9FV��u��̀��$���_8�ٵ����ţ�m��5�CP䃶��R9	p��?�ʁ;a�-O�F���e/HIbE�}c;[�&�4�_�Uy���Sҁ��>X~V��dFg\A�-�IM�v�;�����7=n;�i5u8�(o3��ޫ�0�����I���M��
=Y�e1u�����8��㏨�6�����Y���q;��N�M����f��#2�W��4�V3���C���<x�C&혗����d�y��7m�(eKr��D;Mn�MY�U�h��<;m�� ʄ?\�q��6nu�^?�j���QS��s����G`�.o�	(?�� (�YD��y4��a����OS��X��څ3�/�	9IQ�n&��u��9p6�jSK?�v�2d;u�e�]=x�8؃���\�	y��l�H����i��X��8��G$�)�İ�>���0�^
��p��pH���n�V�?+y�y�px~CG`�*��V=�%t.�r�����щ���3tbabPc����t�{�l��ⰨȎ9��]�GHW�?|����Њ!� X�qQ��	ܖ��m ����a�!�g]�c���r��<n1��E�3~̚�d�x�L�9�_Ւ���A��};:N�FJ�&�<��(_kU]���"�X����EG��؝�Pχa���Y���tM���u�
�IR�?���X��B)�@�M�\�-s�!�&/���PϤ����b��d�P%M;�h��� 5����pڦ�=hF��}����4�O�Nypð����ԻR�� A0��V
�JX�_�٥��9X���1\>�ߡ0�f�t2��}�91��.r�(�Κ>�9��_(���B� ڃ���W�;z�Ń�� �Ù� �@��-��*qH��2��I�P��� ���,�y/3>m����I4��O������o�
��W`���j?~��ѫc���L5����u��p̸8L���r�xU�������M{��ݎ��4E9n8�\�t������f�T) T1NX\��v}Q+{juzxQ��o��%�^�s	b���4H���>�6t�D��`���v�H�`�)l�Od�qk�	p��X��%m�l1�"���Z��N}����:�㞵,�_Q�f1� Y��{{,�����3t�� j1�.:�C	�^�Ӽo��v�w�z�cr�Z'���u2�킟i̱b��3�)�Ae������O߉n�kI+���=�i9�A���O��dت=����)'Y(�Sd5�U��y��֧��k�S�?[.�\�A��xy�˒��&�4\�A��u"89���LG<�L[�z�D��:Av������	�sE��"B��MK�3��g��[�ʠO�r�Շ�9C̍��^�Sn�D��R���p��,)����j�����<�q�dn��s�7�-2�����$��Ձ�4e3W�
�ן����FfT�Eov��D�gP{~�8��v�C�?|	j�51ºT��2/I./�?�ˣ�E�o�[�m���͚��2�D��;ŜZ��.��t�b$9�5$��ń��C��AЅ`͞��Z���H�J�l��g�%��RN��"U�~��MA�����d���0r�q��0''rZҌ���1���sܶ����7 
Y�ߞ�K5��h �?T��w�"^ð�I3�xi��t�37�־��=�I�����t���|*��$�iT�qacJ�?�z��W��Meg���wTBOJ���G��,;
�,�r���2��m �o������k�f9����j�:+��O�8�wʬe?����(2Iܐ\i��_�!�eQ���V���ǆ;;&�1�3�!�i�GM&N��L_���T8��NId�Й3n�9��l둊ķ/�R��k���"劋���+A�[��m!NK��5w���$�gM����%�B��mԟ���=�Z�d]��A�2 ���d&���z��m��El��	�Qt:�`��R�U��7���{��{� [��∠��,נſڇ��/��]YT�/��L��"�dv%��q�Ι���k�t4��4q�qyL��C����־3�̍�KF�����Om#6�s�b�"4P�fY�����	������03ι_Ă�Y�m�P58X�+�DnQ�7ˏ�o��Y����kYP��RY����N>NW�E�ؼJ��p�Y���isD���5��V[lˡ��~�o����*x&���v?X��U�?�n�Qy���v�� �-<,�O��^���~�l�@�<��w�:�^�v��Db|l>`BM�c��_�d�p���ط?5(Z����J�ըc��� �G�m~H꽺�� ]/��7�7�>���'���PP��q|0JxP\xy�h��;w�,]O<��[������D
��B�����=w�0�V�����I3�Z���R�T��3��S}O��=�!T�����<��P�0�e�?�x�ӓ>���E�1|誔��"O�m|,���m�J7�Q�)�ԫ ��9Lw���:���D÷�Y	*t�O�e�<��0��m>�tAwW�v��]���	�l�q�p���7��'e�C�~ f��lw����t��,���=񰡍5����s��R"CW6]����t�ة��j�4����s�h��ŀ��5l�E����ޛ��[�r+�{�����l}�J���*���/:6�c�m	�ζ�PWO~��g��Z�U4>{���{B�o��wM�"e��ͳtBI�	��'�o���y`��g���Hw<���g��^�1�*��I
S`�1V-�[?�t1S���\&�K4�F����;N�:�W�Q��W��b�R��	}nMǘt�˾<��|�%�X���ؓ 9��:�H��!����i��g29Q}4�؈���A39	4��<�U܃��/��Mv�
�@��^?ϓBߴw�gm筎H���vtY1`��3�DZGo�h����{nV"_�����6�=���ůگ����}��ƩW��qw���*��dJ]x�q���������7w���Ot��GJ��-;ю>�U/�D���ںu��8s�?�\�/,�5�3�[�SU��`�k�D�RrЯ�ô�ѓF���E\ũ�
���?�]xӽb���Zz�.Jh��vM�f��ש�suc.M)�خ��|�,��>E�S��
�l���y۹2t!�/x�S؆s3'1�(������| 8�8!!�!��ɋ1ko=J���	�Qt�˂�a7RFб�dl����7�C�f@��/|�#q�>�^��y�_�t�{�l�{��^����]�/��0�A]W�K���ftC�_Ɉa���w�`"1�u�G�����e�B�#���3���ifASsPQ�����k��~81�sDesC��w�2�-�`��i�����0#t(
�l�w6�d2�<xg�}m�o�]�u�����[˦�'.��u��1� \�=\���<�z⫇t�f[�>�m�+�#���ͺ�mH�x^���'#�D$!��M�Իt�f�4B�4���'/ߌ'��A���1�FA����܍�.@�΃Kn� J��W�\ ��Hm�ږ�p���9kx��p@
���i��+�� F<�^ʡ����uCh��s1���	"-s�$�Е�_-{���f
�d�
Ӣ/���/����ng��N��DG��i`����b2 �x���JR�F��k���^�d����3P�f��u"K�kݟ�`�����<�c��զ�O���O�ī8�dy�e_.�l,֯N�٩D,�����ޥ��J�@ޑp�E�pS>R�jT�ធfխ�>�$E��U���5��`������_���S׍�Y�K�4	�����VU�"d�"����ܽب}�ccv5?��ea=w*h�����{b#>�����'`��j�U�+���j.>���	=��Qœ�b��2�:�'�ϛ�7���c�g�\2����2��s&`a�z胤��d=���_��ݑ����:=:K�/�;��K��)�!��&�5x�L�8ꎑQq�y�[3�3��g����ǔG����]���rwo�(|�k�sg�h�5�I�����Ծ�҇�����_�5~��E�1a8.�C��hY�M�f�����5�NxV�����-�0&*�H	�e���(ٸ$��<-����}�W9�~7�3q :_�1�h���(M�]n�硅n�Z��#������w�j	}�;�
���S����7w&�y�X�e7��X|v�mX�9���M��y�{Oc�KaL�Uq��מ,.C0�>q�z��4�ޱ�n��yRa���_���㷰�ɟ�I�F!���	%�a��D��\�����kƞ�.U�O���QKl�O�'}��)z|2���wy�?�b�P.�sHJf��{�W9�#�����3ݍ(WK "��Oli���߽ �&�V��y��었>F®^A��*�x�U=�7�I0n#cYtf�W�,�84�!��(*��,�d`���ʜ|�1�|Y-�	ғW U+q�kJ&�Q���
�;��%��z�ti�ߞ��ة����_b��'��)/��S��wj\�{G�&�e"�Pπv�V"�*$B�N�_T���
�m�1O���m�q�O-�'�+�H�%;�"9B��Y�V���+dX�N�3}��O������������GM�Ʃ�����,.<�ɮ�c��%�c�.�_����D�~ ���ba�C+��	v	�`����eڿT�h҆l�h�nh�u��Sm�}.y����%�(_��Vw��\���Y�{$�/i*78��oL���%�o����xeڡ�������;FEm�����;��9�1�'-��k}20⊯Q���L7��Pl�ň��Ymr����������v��_�)�{`2����ԣ�bp�������{67�:��)�Ҹ;���/Qq���Ex��Lw�1Z.�2V�uvl��o�-�c�7�?�:W�\d^�E�*���̷���Od8���8G&x�|;t�l/8𾙳�^]E)B�C�u��^���Y�r+�;2��6<o=VR��׬ק��YV3>�M��m`z[.�*��H�Cd���g	��z��N\/Ԓ������V.���_�Il��]���V\ͫM�c���ٴiX�ɀ醜&_��B����Re�3�2K#+���_������j�p٧�çs,�뷐ŷ!t���g�~��a�rM'�-W@�D�j��$�vN-$� �����~!3:9�S���>L��}n���@���̑"�h7d��A�@U�դ�z.�r��PnZ3��=~H�k^�بf��+�:M;4�%ɽ��)��I�����?ksj���e]z?�EN�3���*��W�t_q�I�X��^����/�cM����L������Z�%2�O��~�����b��c���y��A5n��4�U��^��J������M�{��jE��������]�_*"�i����9PR�QFVI�SX�^1�f�Yyu`Ӎ�SZ���/gZ���򇙥1oPP~+��N�3�k��n?��+5��ؿ���+Z��9�������nF�	�D�!3y��w�+��杁z��#%���i["�4Cm-���?Pő�MX7|T9K��Nn҆K^t	�s���=��uA���G���|W���H�>"�mHD�����uK9P�Xb+ǒV�[,[�q�«��v�j!V
�.c_���%�㦿F��k������!�rS�k�?�i����:������ov���C�M#��u�������uO9K �6}^B��0fZ_��Lf����w�'h|l���2�P����� �����E�AuM~Ev�Z��v_@���6;o»�CNFc Re˔FF���(7}e�4#f|!��>���z����oMc���o��S�#̝�.�Y.�|��1�tS{ f�\An{�V����b>I���������!P���x�p(?��D3j�_�6����2_���ё۽�$�jZSd��B̘~I:�������E$v'w	�S��Ixǒ��5�/eb�����H����<ɥ�?����՛�*'������,���i�D�۲$���f�j_z�hѠ��q?��ӊ�}�x}��(�q��Q�15;F"��2��|����/w�|;Qm�K�au��A��{ʚ��{ bH�ՏD'R�x���G�m��1��E<r�n�fn���d�W��L�!UT���!�T���[_5�B�_�kze�%[9��][G$~:�o�P�^�3���o8;� B�x�@i
^;r��%�]�;��� �nU�K;��y��:d�
��Ǣp���j�Д8����I��P��D�W�o�/UOZy�pt��ڊ��!)����D��T�3�c�O[z�Q�� \�Ʌ���L��(m<��xw<��O�.Τ�]��)/�j�k�Oơez�K�C���=J��ln�j�
����y�~yq����m3�
9���H�bCCu�~�n�v|i��y�
��T?���2~x�|越t�02�:�;oTP������h&��a3����V?<(��\>S�+��uU��e�����j��1���XL�?��8͵t\���oj����;��N{0I�a�O]"��i���� ȴ��o3x���K \���c�s;m5�'���h�=�܂� ˸gQ�E��w\!� ۃÇN�BP�?��ѡ�>��6
,wn:���*#�j��n�y#�{����گ�Qb+�H���""�,��r��Ի��@y4�@"���Ηr+wg�wH�}��'��.����E��ܳѨ��;����F��W��xx�P�zT���X�:wc��+[Y� N�I.}Ez�A �ՃZCa���>�x,C�e���{2���� q߳�:cs-�pD�n^C���_x���c�i�h˅�]��q��!�\�#���~E��{��ߣ��OJ{��r�.N[Eį(�aȗ�5�Z<C���^P�u[M��=�`��I/h�l6`�e����J4�M�{*GP,��E�(�*�>�y�����u_�,2�3�8{ɴ���'��~���z���f/fg/���-lm�&}��z��� �XR���}lc�WG�W��SCCVP����zR��˨��(�_�2���1N�'�8<�Dx.$��\���s�\�7��>�|OS�N���^Fs"��X�a��B+Ã���/Ȍ`9b�c�G�_��}����m�%�{��j�K�g���o�����&`�o���ǣ&�ߓ/�T������KQ�o<��7z'�P�}�Q��E��_���Sc�!ȟ���M�+j��0��E����vo����f�����M��ᩆ�YA�_��f��E+B�|+fv��_�#��[Q	St5]z*��wuoy��#$��#�����kɾԭ�"��F���Q�X�'�{��Ƞ6\`��2��$T��~����G��Y���&4���^�*�l�6���.���!�����ý��)�陰r�ͷ�6rӔ�&�Č�f�<��Eqy}j��m�t')���|N|c�
�S^�ق�SxW��>_U��v愘&ƌN�z�;?1�g�O�{NM[1*2S���g_+QV�Hr�Ff_Dn�Nhv�H�p��ܢ����:�=��[~uO}�yI=[��M�I��3y��L��ƌ\m��&v3D�I.O�3���V�K���wW���J�B�˭��	�~���L*c���vǷRY�����g��򝓬����8��J�Ț�O˼�_�e%��{�_��lU��/�Җ�j�ǎ����	��u>����-���;�a�`��D',G�U�(`�����Q������.X�S���[������kW���
1x ���?>�e���c�~�T�:/�;C^�O����pM<�s7��#�	t�9�7��P���ɚ������]�����u��o�l��Z�\N�g�n�Nd��S,�f��-�w)|�;ŕ�s�P��oAn�<e��EL�K�a�Z�v-Ą@��v}4�v�ؙ�_�)���?U\��z�=Ea��¤nh���5�	m�φ�����D9.��JR��D:҂?CwΑ����g��C�l���'��m�������x1h�'\�k;N7Iy�1��:��'�p�M�S�5��B�°8���L�#[�[y	���ݝ5�WR���oL&P�Ӑ�(/Zܪ��L_G|�Hn�VEϳ4 4���
	ÇKS������ܣ�� �� (`访��~�0�8��_���)v���Z�OW���)����FDD�[J�?��a %HHJ���1B��;F3i؈��^��e׮}z���>����EN7�rϳ�̅�8x���u�E�������g��������sgd�)��iQ��;hU*���񕞐�q�K�9�n�	���ԊC	|w	�T�]�U�5<���*�N����:�À,�����98������/W��]ی>=t<5�����Z#%>IJ���ɘ!MGl��XV~�D
%��*�Y���qlS���W��c�G��$V�½��Kuj��V�~j%��OKֳdåC�8m��NzR��(5��-}��O�=���f��<E)ִ�9�+�=�c�{��igk���jg��*���D��sz�*R����}����R�'���"�p(���f%͏��s�V��궮�2F�<����z@!�OT�"�Hr��K���ZF3�0ԲMuD��]���i��'8��&+F��[��sa�P��>֬���Z0>1�M;��]�1�*��}n��fH�GH��J��W�3��g�	��	DӮ�\�"�w�\N����V2������D*�l�V���Ll/���$�K�����א�p��6�rUN��|�qn=���H����1���}�"�5����( ��707���� ��d��AD>��U�`ƽ��w����㇅�j2oY��z���OU��]��&N�!�2M{�m��_VO��҂�0���Z9�?����74�0>ۓv??��!�H�"��xKC�db)`B]��n���K+-&�,�{���DF	U�8��8�<c�}��/#X��{���˶%�{��;0u�T�
�{�u'��ݜ�%|�;�S�:턦��Z)��5��%Ƌ�&��H��>,��X1̒���I���X56R�%=/ ��SJu�={e���a����6AR[q�������èR�u�q�l*G�C�uT�h*C4��Ż�=�	����Q��tÊ�	wy����~��P1�ټ��\�\l�����0�9)2�el�»2��LY�$f�7��wBW�Tn{A��m?�li �����S�=� �<��'�����:#�떍xƺ��|�)�u�9�\�3k@�����r����@��7.1����4R�H�3���g�~w�/��vf�F�|�
b� �+0jM�V����X�}��Z��?L�_"¶,��W�����Yq�مD���
ĵx^F�RB�%����[�<�#�L�@�C�gʏAB u��t���Ҳ��ӭ��:��J[Y�N*�����e�����`|�Ȝ��bR]U�Ga��x𗸾�gZ��p{�˺%%vl��qh��������(��l��*�Zy�'�#ǟ���s����a��6>��z|i�::���k��:�o��^>� ����4���SF���%*V4�B,�<xٿ�'��`��
��w�1�"c;3��wJ�]WӰ��p#�L␦�EI �� /w����J�>a����#c���ڍ� �l[i_�kLN�uEV�l�ϒ/w?sY�Ol]gvu맏6Rv���B�����}P��8Ee��$1B�����	s�$_d�8�}}͂"3�����P��5~�tƒ_�B�霿9�P3U%^�n�9�`a��O�P�J$������"���������Te�-=k��L�J`0�z�4:!��HaaeNs?{����?�m��p�<�����h��nO>e2T7�|������z]�4�!cu47"�}O����d���1��� �������'r�R�)1�w�u��%A�PͩZ:�W�w�t� ��a��O��B�9ʚ%j�/3T:�[�s;7���*���M9<Y:4N�:f���q�D$���m�:������-��ks'�����XA���ɲ��5-"��@P��Ց�3�Pw�{��>����_�B���p��1XESI}M����U��c@�z]�w��K�"��'q�ʎ��bUG���˗�{fOwUX�V�{�I�il�[g���ڣ�5�Ϟz%�G���μ����:�b�Vt��C��C�[�#*Q7��WqT�y*�YZ�y���(p�Ua��U�}���܋l�c���������*T`fg��!�9W�h�D���ne�˭���W������^��Ϟs�1v4������yA?�办��7��
�6�aYDN0cM�L� �bњ��/\�Z�5��w�N�ohA�7r:6_0���}�^wS͘���d�k��UV��Q*d�<��r�~D3��1��`��&d�.d�,����m��5r�%A��is��X��{3�._��	6^�4���ƫ�Mm�� .O�!E�#Z�ڋe*�?�Ty(^��Z���U��K8e��4���Ĭ���X%�+���e0�r�P�@}FHU�.窄�,>F{AH��{����A��-��~���Lf��V���߉�Y��q�W���Y��Z"�7u z+������JI_�p�W&LU��#�\�L
�7�io��~�/��V�2�+���S$:ȸX%�~^�M�%Y��`I�y��"����#���8��`״��L�yD� h���&(����G��N8��@��.e,ˋ�%&�pO�
�NN�-~.N1}���=o���n�p>�Y���E-F��6�VW�D]��C'm=�dx3	�M��G�n.vE앨�e�~*KtLRUF�5�Oõ��{�9Xp���������K��FlZ���B��Waה��aJ��O%��[�ʤ!�)��G�a�,��ƖZn�[@��5S�����s'����9� #��z���z��� bQ_����6�{�`�������X���+��\?��hÑ#��pb�w@uJkF�o�F��tz�G�d����^�L����nZ�$��m$���������*�JzUGW}i�'	sh�s����i{W��D�;��>��UN�&��j�x��4�&����t-��N���7�R#�����%))r�nx�?�޻�)`�j#��%�$ �̮���.}'���r�H��lt\=�D��ΙC$���Kd�8x�-�V��e�u?�M��#�7x>�=��?D0ΰ"^~47���+G10z����ɱ�EWb�t�0lf,n7���<Ac��եƢ?�|fw;V�_�>�/S��+K^��Q�[X��](�y�p�jr����L�;�J��N����m�����z��q��^���``}����U�X#���J����/6��U�)��iH�]ч������y߼Z�ԯI�I.�b{]�m�2&"�G,�k ��0��lQI�_��v�%%޸#�5�~䦥O�+���'��8��ז�\FY���/�Z^ilL�C��^��K�d7N�c��F>�;F3�ޤ	z:�i�"���cPT&����bi�/s�ޚx�%Id���c%<`���.�_!-���*���H�����@�nN���W ���1�^��kÛuⱽ��Ը�Ҩ1��;1���s��1�A�a�Y7M5#A�O���'�Dv�v�f�a8^AH_)�t���:�jG39�^��<�e�Q�8�F��K9e�_݉�����h�x&� ۺf���o��Gii���-K) ��լlPE��:�]���4R ���ek:{G���WZ�R�kݪ�ժ���N%+_��[�15�8�[�*i��`{M��P;���~�Hso�h=E�����d��<�����[Iύ@���E A�ie�:�vR�(�ҍvKݴ��)�E����a�Pl�z���fQ��Q�79��' �^��8�n�D�<�<�mC�R@3w�f�q��40�A&��kC,/G���ܨ]��l���`h2���@�h�m���F��]4Qa ������뻲��l,xSu�j'R`to���V��������!�u�S���c"��w�ٕ��i[�b)mW
�yhp��I�$X̏w����ͩ�8�B��g;�f򟾌����#�o0��V�6O�FR��}�����0�`@n��f�a^-#a�y),��0[W��q4/�#`j���P�if���o�� �܀E�6���T�*�雏��+`���~c{�"���6Ƨ�
a3_R�%�p�x�<T_�}��i���K{7 �?���cpSV�=���6�ie)��x�Df*��'Ƙ";�e�\�������Q�?��K��$ȓ{"�vN�K	�j#Ǵ؊P)����(��*�>��s6��࣍�gm�|��eQc�2":�䰕3�Q��o�8�G�L�#>��温�C�s.&]�i�ń-��H�AH�b~��ȿ��)^��\��frT�3bU��.��A5�T�t^3d�w���������Y���Z.��[��e��b���P�j-|����@����Lr��(E��d�w��!������$�|�Ξ�RrK�
��#"�sê~3���9��b�>Zv�{�����p�����6m��|b�Y3�B�dO?���0��늵��<�q�R������Yͧ�G^�<�p������]���5�9�x^�D����u�r�}���h:�P����㯏к+�M������MzP��x?�'E+�l��Y�J���Lis���!�\��a�̒��TA�C���O�\sZT��3�u�,�W�����J�ߪ���hq������Y̶�� �LV:�D+��TX2���T���)���[�˘uCn���<�wv%z�k�P�L'�e؍��\�	e�=��8�Y2�ݨ/�:��h���`Q=�1P5:�4c�X��f$I�nT}�r���M����[�����pz�6L���Zp��ݛ*;lw��M��m��;�W��*?�)���?a�95-��G(E�X�r\�j��߱hM�W2�CMM��M �И�`��9���7��)�F��a��$�	��RO\�R���o���c �C����q�#q�bDH��:�\��[�Sf"�}W�ߪ}>�İ�5�� m���[��86�%�(�
�]|���(��*@k��|^�y������qd��!o��vj���j��(�`wuzY1�_�R���f��^��$*!��[	(��|����u�=�a)��9��E�	�w10��)q����:�	a��(ܔ������ߝ<S��Y�o؃���@Ea��N���з��,Ͽ���}B��,s�2��#���#}����sW��Lز��5|��������
d�vN � �L�/4ٍ�g�1د]���[N�b�s�Srʊ�35q]��\�L��@� ?�KvM �W��P�C����8��� mJWy��b�A��_��p06��?\F��������N9ӞR�i66s� �I9rOi����9��#.<�W���ڴ.��^�ؼd�w>�[�O��(�QJ���=˰a�x�o�+MmS~#�*Ua�,�CU��8�W�ĊK�x�]g��	3�����8�t�o����b�E<@���sl@�*�hjXc���{8Ps�Fz��N@��4���cwu!���S��sNC[�~����J㴷���v�Ůf�2�7�N�%������2Ǯ�!Y��]��7x��*��d%~�	ڇ��O%� Dv�)2�����T=�r,HR�?�=2J�P�q7V �N�ۂ���P~���CcI9P���).��xw��,-�쎁�[k�>��/x���z7k�0EΚ/�&/��Qϳ������ܸ ������n{�ZZ���2�	U��b<����ٙ$�+���_@;�ww��;(RI�%�U��٪5�{ǞX��P�4۲'^���O�t��`���ܒ��z�M�m/�{$MP����� �'����2r�����H���1�R�}n�Np�ގ��I�)(�e_��k��A���J�^� ;m[=���O�5/�y�~ᔸ�셹N���/��K#MF[0a����~5�X ��CiK�֌~v�����r�	��tm	����Z�����Q������a� �]V�'���a�t�tN�w�����G�ݩ�SJD/1Y�g�W���_����$�E�	��b�p�id'a�`�7�Nt���N`9��i���Vq�2}�2u�����4���f ���*�-d�4����a����8v�X�R�3��;�46G��c:�:Jw�E��>��P
B�쥛ކ�ڊ�'��?!��`c~���1�Z0=&�"���o�[�©ʐv�ˎQ��5��]�'K�����w7 ��(R��c6������a��>����)�fk�_~Hܓ��pt~��3~6�x3�v����|���G����9%b��\��Y�ɈH��K�����K^�Li��G0������AN�wJ�P���!��r���*�ZY㶑�?H�F �:�� ���� 쉬���S;DG�î㕓2��o0� �EE~�����+b��]u��w ]�����'P9y�{0�`�8g*�{-2�v�"����Vmϓ�Cw�)	f� ��G������z�u��Z!����$-�����Kҍ��p��^S�8I!$�T2�8�2FZ(9�a����&Y�q��p���A��"��$(�)/՞<����g�v9M��?����c�W�c֛H�4�V��=#RC�t�91�K�jr�wI�ةeݵ���
��ּ��6g@$;�ҫ�L@ͧ�D85U!��]SZD���+'v��ࢯ|%�^�
�=��<4�U_�u���-��;	�^Ra7��K�~��~BA�V7�.&.������/�?L)��4��Ȥ(s�wXQoB��r|�>�
�Z=Z�O�,�'4~B��r|{��ISv���/Mù��M1t�����W�e��Pd�z��s8?��=�׮*�G��`b0_����z�����=�Ѕs�#���䷒C�ju�bм�1!�E���𪧖�#�\[�mj��ǋ��,/Ӑ7�ˀ��J�6�q��c����d[�~�J5���v��=��"(�zu��&X��G��>!�e��'�⏎,��K>�~�t��aψ�!ADEUcH��c����S��^�A[g�!H������
X��^{SX XZ�|�w^�81 �ڛQ������}��½�ij�<�kuf�݃�Z�G��u�}
�����ޮ��/[�Y!�r˟T��p�S���T[Bd�z9��!]�"��!o�,p�j�t��ĎX�2ZFCZG	�%�v%%0^���b�+BT{�[��rl����#��Ā����b1f�G��6��~�����j d���K\���D�h���"�?V����x���w,��ėۮP;A�m�I��|䲼�?���?O��{������.��_H�(	��qFbva^�r G�2T�p�Jd����L�]V<-I��}ufwн
���=q0m%1q���+9A����V�0P�g��?�`ohE��q�d91�_)l�i��S]"�m3���t�t�H>��RՃ��?o���n�ū3��vן׎^���zӽ��U�SS�Ll���nL��޹�앚ǌ��+ɀ�Z�W��Wb&��Vb՟��b�ׇ3�2���_k��PW�.����^ٳ�㎚�&d��МO�x@�u] :������N5��-�����qX�N���SK���YC{��&s2`Z�uc#�/�����f�����c�_�ǚ���h�^~!�<S	��(�[*���wY�fhr�:�\�W�C��E���?"i��5ל|=�矝�S��0�lEw�nz��Qx���=(�9�ݗۈ94�pzjv�\��y���U��˱摠±�����<�Ę�Ef��+;O���7s�Y�Ɠ;͕�vВW��Yw>���',S���h8o��~�jj��Ң��0L�^)�(E݆�TE׏a-)n����m���F-��X&4y���0�<�Lx�?���K�$y����Fˉ{��g�#]^�/����W���<���9����+. DO�������F���V������,�_��Vsf��3n
�1�	��B��b���p�K��;�w���R�-�)��X�.+N>_�2���	�
c��}�V2_����x!i�=����b��r��t����H�����O��M��5�Q�b^����)ߡ�iֽ�W`��c`�H�cO�0��˰I1�+_�o���'P�]�߶���� Fa��l?�	��q���v����TCu�b���Mm�~�zh�#e�٪����P�t���8�\Xd�=������Om�h�+��[�M1r3�!d��߲�
�	酟|Yi�dw[r���Ȃ#�<��7��g�u��)���[xM�Z�=�5�V�<��i6�"P8����l�/|5�#�q�bO� �����:��-�5�����3[ώ0��#[Rw�@�X4�q�~���&z�/o맼��	����5V8���p�?�5�j��؃L!��v%")ۭj�h���+��yjY��
�Ʃ��b%��l�Fc?n\&�8\�AKy-�r������;��������r6��&gڿ)�;d�����f�ޓ;]�SL����Q|�Ҙ�E1���`�!�����9�z�{H~���!��n�&S쇭� ���~$��tFh�	���w��\{��Q��9��"nw��}���݃�E�(�"+���	��8��t	D���zm���͞xjm  �J�	�̽��*��]����`Yl�9��4��4Q��qe�-�O$v�s��{iQ�%O*�11J�vF��KZc(��W���up�zN)���l��6���k��Σ�n�~���
IJkMĹ,����`�z��|�,p�I��c^l�P���weY;�B���۞d��.l(_3�a~��Eb'v��9z��vS�=XLfIx�"DϚ]���5��8G�g��5E߀�.�mV2F��ʇ�$�!�#�����[��+����*K�S�M�Vx�aR)9���v}�5�p.��֜��,�a	X�ae,���ɩ�
�~�.�W	�I^i�q�g�jl[�C�_�m徨恭�J#ֆ��7C��vb�W�޴���==�`媣���޶��xQ������*D���Oγv�Mcw�v�͢{�-�J�
��/��җ��y�9B;Y�e2G�b{X�No�(%|yI��C�n��~�C��!����wݨ?���.��h���D��(pDD�e��+�T��Um�����EY�e�ԓ^�_)��ݎ��o�Q���q�ȃ�O�+��탔U����>pޓ�}0���~l=�,>K@�A �V�?�t���x�Ǆ�i��m��-] �uo����o�5�; L��h"�!ݹW=yB�R���/��*�� ¢/%�F�� �|��2fx�孕���%Y��=�E� 	#	�`a�T\XV)y�������&{���g�H3�:���K��<w]���mf����~�S���m��4�$�,:G�?$�nmo $��U>+duk�aF�]��0�ӟ�~앷�PGf^2�w�2Rn��U|uɎ��w�>�ᵕ�[5)Z���:�?ā��u��L�>F1�a
��X�������p�;�f2ӏGm��@UF�G��Ew��,��XQ��f�.�&	�,,�����/o}��>q�Ej���Y���0ظH���
t�%�y������؆F�;�zh���I�G��
ͭAj��W�Q��MiO�"d�&oO�R�=?4�ܓ�������[��r�S����?�����1gt��1��-� ��7�羛cIe����W�/��B�#����n�b�X8�ub�̌�5&R�������������U�쩯��A�4��R�[n�<r��ʵ�X�߉N]�e��Ed#��ȃ&�+�,�[V�wR~l�Ç�%�8�>�3:�:�n&ԟ��0
���b��r��2]�z�K��3�K��C��^ƞ�Ɂ�2���n�W��+��YM����aӚ�u���ݗ8e�`wa�D�Jf|��s`̥�;I;#֟"��Z�&��ڮCiW�G
�e�l��|��j
�)Mm�������2�;�0���Wz�t���N�'����'��F�t������w���\_��u[+x_��{�ɱ����H���zClԶ���`��G��-�̼�<�!�Ng:FV��;�-����������r�׶�,)��y������ϭ�����%�㎮ì��'���\�Ed��t�~���&L�O0:�xOX�?���?������c���+u��%^�|y�H_m�cq2Ʒ�#G�9�`{��wM�jl���0~`��FO��3�+S. 8b^xAC\��"1f�W�_�1�y��UC7\���>�[s���詩��e0�[&HL�)�򺎏K+L�R�WR����p��� ��FA������4��N�3�"����#*���+���%���(�Db7[+�!�Q��ֿ+���N`��ٕ=�e��ʐ�{����3���%�7փ\h鿞�a���]d�3Te��9M�<�� e��"g.M���������m;��~�p�?�����!�Y�]˗3m�+`��� `��-G<�U��q��I��!�Z�A�	��՗oŠ�K���ڍC��o���ĺk�M�>Q9�PҲ�p�K��H�-��c H�>dWGl�ٳw���?�ʛ��?��6u�Hb������$_`��ؐ�1�I��b�T(&ڐ���b�I�*�bA�ؗ��E'$/8G��B����9	���#�U�+J+6#�S�qk��dy%=�.���O���]���~sG�Lx����ؔ�t�xR�M��ŕx�O�$=�e�,AO��l/����:����ѬK���\�hnw03_E�-�&˭2�%~�Mϱ*�X��B�ZI2k�;d�=��`N60]M�bu���wѹ'�xl��$i1IQuA��[����r��e.z�$5v����i��{Y�� ���jW
4��jY�řm;d��tn��,�SJ�yRZ����#8�-yܸ�X���2�5�@ïL�#��'�m4,6��qM��@�r֌� 7��1E��E���9}N�S6>{���5��z`�G���;�f�����K�^Q_�B��-���G �x�/��q@��j�@^�J�<�d�v.�,"�@������cc�	��k��j�并l2�a*sq��(i1q	���^#�X��`h��b�ET���Jl�M,(|���e�V�e�o�m1���15v,m�5��0��^u���6�>��K��B�ح����[*k��g�`�1#��
j�-�M�p��w�jK�J�u���[����m�ּG�qu:Q ��0� VҹQ�KB�9���U��?�}-�d6�Tg QO�u��f�	����F�V�ʆ��-l��a危Z��u�o"���/�>�s.��a+q/��?"T]#���8^<��"�ihR�"�*��i��I������OA,X�3��բ�w�.S]`Ɛ�rwE�cQC).�/-N8V5\y/������D��q$��9�W*Jn���DT!c������e$���CW3ES}GI����B\ʻpڰ>}��>l5
a�ŒZ�!O����t�x��M�ue�\���4>�t��*-�>")�����%��jPó@�,&Rx	i؜f[f�ɒ��K���E��kf�5�ȽW�+�#����Զ����4`O�[����� ��5Q1`\���M�k�\�0�ff�n
��1�u�`b��H]�W��\�U0Ӆ�Kw.d3C&N�VkX����|*��D�FVn�5���7�~P9'�՚��$�����
�Q_ñ/��G�৲�l�H�Y|u�C��W�tLK��|��tt@�L½v�*�h�l�}�8�s�B9l����xC��c�p�����o'(^��Te�Qka�����]l�/#:�2�*7��	�~���GS��y����4�ȶB�i����qw0�Ӽx[u�P#N����f䮠��YG����Ѻ;�w��s}�M�Q"�-�A��qv�w�% �Ų�ܹ����75p����n�#ii�h�!���+s�!�"pV�M�F�J�Z�Ŵ'��B�'ٝ"!�g_���2����i��c�vl��|����l��1��"����-q�����TK����E��U�Ǜ=��*�#�@nqpKN���s�}�%�QdJ��t�Je�+����j;G����(di��)ى��[ѧ%����������|�O�'�[��k��8��J�W�At����JBNX�g�}��`��>j�v��}4�����z�Rl�I�!<R��1�z��*U���3�ϧ�����j�R�
v>��z����[Aj�8_"���f1�U|}=Ԯ�{�ջ���<0�ƈ1M3"I}�R0U�\%>��Qˋ)�oi��1�0�!�m�a=��4�0������������3�3�}���a\�";jB<;�	��#��>T1�tR{�����"���;C}l��`0�z����04lb�i��a���J�ō~e��7�>+p|�!>lURm�K����/��zA�dC^��@�1e��,�hC�|��B���[p��w��<Ԫ\%�� s������4Tz|4a���󿣃�w��0�q�Xr��$��aG�?tmbMp����6���GazT0��G�?m����YB��BsC�����������C� v�W�i�����O��803�E\�.GFY�0$�t�p�
�f��}{�3xF���]Ԏ�����kmY����%�"�CM�iϛ/=�\G�|��E���Ng�;��J���b-�����R�`��<��z.�ŵs�6�Ż�xH)� �;7��͑C��x�	�]�����n�a�u����s�:2���i�I������&\R�G��^`L�4�E��Z=���F�ȲD��y�~/	���M��C��jI �������(\��r�|���.O��~�R���\������4��Dè˱�&X��3������ɨ����R���]W��Vf?��m<���C��ڝ����^��F4q����[�ΐ�T{�R|��-x�jDmۿf����{���!z��T���F�G��L�7��QB_$L�����&��tʌ�zM��U����5�e�ֳ���b��X84E�dϫ.@�Q���,�y��z"��xӎN�QX+�y��服P��:0E��r�]Y��h�u��#>S�>�*�$��S�*"1�d�k�[�k}Md[�:�2�z��gy�f
�=眩-	��2�y�)����wj/P��x@�����n�M�^M�"޵c�{�_o�M}=ѳ�59�L'��������F�OHZL޵��k��Y���*=�A;���;TU�?w����kz�4��s]�~�L�����ȩ�8	Ȥ����"���Q�&5�����ؘ�L�]�q�G�]��%E�rS�	n�gZN�/eJP*-�'�Q��S1�G��E���X_�m��4 �ȟ�r���/^���0j������s�+5�j���w��)��x#��B��+~��%ʁ
5��?|v�u:�����x*������XlJ������r-'��S�HoP�����v��D�T���R�Q�;i=2�-e�l}����k��8;���X2z�澔��n	�zp�*q������X��k!6Z'�C���8[�0����ӔYb�o�����@�3�
Wt��J��}�昆�,?e���Z(�FE�������7vP|7����f��̒�ރ�ko�7s�$�?kA�bv�3�q�R B]��#ڳ�x�ٴ��r���#�XL���X�*���-�e����o�G �/e.%r�Յ�D�h&�R��
������R9-�b�'l�r����f���s��ݟt�[׮*���T�Z;M�u��j@���(����I	ޗ�!"�O�ӣ�L�M���#�Vx<����GoKd�bm}�ܻ:5Xk������1@F�m���]x�)�Vӓ��޽��䏥o��=*����h��(��#Y����8ɯ��=+Y~OF�5�I/�|��W�u?<U�������/}�/��}D2wl1+�h����Hh��b�g��-�n�&]r�}��%#Q�Sl��l�M�L�6t._�b��wL�� ���*�g�W9�L��d%n �M�+��ƛ6�Er���Wշ�L;�`��-�7>��@��G���:*e������WJ�U�����m�U	N��2r/�
~.�/���0�,,�ғ0��m��=�T'.�R�S��w1"�U�������+��9��+�4 l�%���1�NΔ�Q�J_���]��rKwq �Ya���}ޝL�fk�ć�-LMܾ��������e{L)����o�?�c�%p訵d,بUUdYO5`7�۞\%11�� �ڮ����rx�x�ȆJ��9R}G�b�)cj�7=9/ϥ8�O�-�<l��B
V9`d���G�ozc��0��Mx���LZ4�G,3(�M�i��{i"�0�!�yX�7�cs�B���m�*�'�yP�6�'���M��Z�����;���,x>x�*ǜ�}����_�F����:D4��:�ڲ�!�8M�X�%*�d4��ƀ�V�)����ʨܧ�T��S���{�P�v��$�|��{S����抇�Ӽȭ�~����2__��vp$~�Z��������<���q��*�=-\����(G��Hg����0��p6C�ͱ.���.B��վ`q��@�[%o��]�W"������z���T0Қ��LMf�fAL.�У�3�̶6�x�ɺ(��B�L���=�^�8��Q��?���F}G�N\t���vХi9J�q�.��@ĶE�2��@�V(��I�i*ь� Jj�v*d�]o�Q_���ך�|��GZ����M��Ƣ'4V��"�s��|�n�[iZ�L���iU����X�t`�����eJ���QN�W>��;t����'՗�D���#Fê���.�o[O�\�g��y�5O)���r�����>e��ڀ�?�f/'�F&_˳i�Y�hyl�>:b�p�*��4+Xfg�yQ��ې*��?6�~x��}Z�R��i:᱀¾J�U"	�$Dl~���2�e���q8�W�~Dood�L��R�Z	��4��I�c�nɏ�-�L��}����%2>���'��}h[����g�}�`������K�M�������Jk�*�29�trD��e��+8iJ�J�Z\�R~	�if���mYܑ�j��̉�UE_'�у!�nu���\]��C�gO�,�(��"� �O�(��[4��7���T,0����	���a�3���V�W&޾)��F��s��3�2��rdX+�4N]��jKu4vݡ��o��h�\�� ����#���9\�G��E�*0�.��p	�Ff4��W����v���땝��T{��,����75���[D�3iۤ����L�d1�d���N;_8=�m�i.���F�{k��M@��?�����Qsa��媩�?�̃��>;��H�K(l����1 $cT�a~���e>��7P�I��ho��׏O�X��&n�{�{`�	~مh_�L�鼈�!_�83� ���ոJe:l��Ŗa���(��E�����C���T�V��*3U��P[���G�9�cy�;�s;q�Z�c�_.Px=~�e���F���=8V4m�,�ݙg��ޮ�_���Y�"^�%�V�)�A;{hz�I'�i�7 �U��kѻ�Y�7!����1��i��^^�@��7"�?vNY�4�,�/��|��!�"x]Y�S�Հ��>=s�Q�)�{8<�ԍ�{��G+�{����A�a��R/-����AĶ�ol�,��E�Fj��G	^��I��8@`�qN����-���z"����)�I�.!o��4y�j���B������}��JKJ�1J����j`f>�܋��^7Hq<�t-�P*/k7��R澉d\�:����v�dָ�6o��+��6������
�M#Y��B�G�6���&u�������ݟaR�������5$�X�i���P���.��f��%A�<P"�!���АQ'��p*�z?U{�����VfrUZƂo ��$�����O�d�VU���_-sn[�:N_ ��}�����R���S��-"���М��t�v�����.幈�85��H��=�ދG��7B�M-�ٖ�P��޼��5z��Z��*EyY�K��T�D�����M���-ۺ-�ͮ؜�X��~��a������Ƚ6�fUГ%���J��Θ	]��F�WT!�Y9�d�����q/ ��n��=aO��j�׌�^xgw�㜟U<ҜP.�y����ę��G9���NF���5�̭>_hG�o����}����C����������wjo�~�f�!�s���\����qjԌ_�Dg
�|�磟yЊ���O�����K�mf����l��	fjj���;�7��V�d6t�Q��CV6^h��n�Sy�s��Nl�+Tj�y ������狥^�*Go����z}��S�����%���������lW�p�i8��2���R���B��mhĵ�+�cP[b7��Kq��%:�+[Q���UF5K���Wf���`�	��N�̷ǹ�M�:�a4�~�H�hH�l�����t�M�mFBRZP:�т�tK��T�$GwJ��4HJ7#FH��t3`��c����?��������̃��#�m;
0e� ީ���c��a�T'R��TKU':�cYB����Q�~���5MY3��Fn��p�t11覍50eм8�'�t������u��hH�?�8���C���@��e,���$���`�W2�&q!	N�z_�r�mU&����Ǯ$A����r�{�m
�0�v�	R�H�V���#wΚqp��#%�_JQ\��S�����h�6T��tR��GJʉ1��I���;��n�{�|)o�21�n���k�ą�tT��Į�&=*Ʋ]�}����.���c��j����>���tEX�P>xĉC4L �:��>˹]���8�:#w4#݇�@�g*
���䝡��u7��1����mu=mN���&�	�|��X=,G�_Fͤ'm��C���N����}��u�綿�=����-�ֹ��=�����<���Ƥ��$D��5�i�s눝� ;W��{t_�~4y =_%L�&�ըR�����IH�C��Y \J�=����� {e�Ƌ�|�b�|�O�C�ϹW��:���_��`w�����-� !�d�N�H�ѹ����E%�+�e�}�����PDe�Ƀh��n0vHߝ�H�n(��G�l�p3�����|>�e��(��kj��=_EJ>Bܭlk��l��nG�N�KTet]�;�w�'�]�}L][R�S�n��(�9bI��=�ߢR��T������F��E>E�ϭ� ������՚�ct�ne.͟ֳ7ʖ��l�q��<ʧ��ɨv�w'�n�RE�oc;>[�BW&��C����sp����d�濜X����[����5���s�S����ޱ�DtiS�`9JP�8z�~��0��w7b��2��O"�~;{f3&dO�G���Ⱦ�(�g�^�@����4�'1J�@��$#3l����6���?��;jxX��$
�_��%�(��E<ꦴ�Q�ǼB�p�]�K�^�ۺ��б�B�#�(Pc1Ҷ��B	��ա8�jw�������j���+@�9}z��M޻�1� �,�ܧ�3%i}qP�*pL�0A9[5������8�I��Zi#��qWmaiy)'��u��*�jFS�g�`Ɠ&M�\x�|,�+�-E��$��n���-wr�n}���"c[e\���0֟��xb𐑨	��E�YOq9�k�s��$O)i�cg���j�N��N^{�ɯN� �t��.���V#Cn_k�b�/Њ����|6���(�Y��;f��o�	�=�گȸ+%@�~Xs�%�:�������C�;宝=dgOw���ʡv�X��|3���ay��q����L4������1PuMq�>�x`7�{^�.�E@\� z�YO�v]�څ�`Wih+ʽ��ׅ�mK��\*�yey�A�P���nlr�aM�KmF��F�x�IZ�'���25�����w
�1�KR�";�6�0�Я�Ksw��E��;� 1��KF�FD�6��s�:C��+X���Rrq�`�7� ��G�<����k�7��l�j�54X��d�NŨ?ݦ<� ��j7���k0^��t�^N� ӽw����e�w�fF���[5�߿��&6^Z���Z�!��dW�w�g���'L�? �q�[a�j(X��F���1��%P�K��(�>���_��PaaV�W_&�t����*��րA�|,B����GE��/W}�<8��;��8��҇@�4�ס��>��&��G�p£�0ʽ;�1�T��P8k�ɝe$��N�R�g5�(jw�:i�.��d�ߺr����L��c����߳UF>�y$��@�]_�b���������+��H��6�`a��;b��1� �T!��I��s�HxC�pT��'b$vF��9���4=��b�t�m�X�F��5��K?�p�� ��[������~]�F��1���tPг��'��M3�ݓ%����+Sk��Y6�_�∽��� ���rJi3
:�&��w�m�۸9F�J���ц61��E���q�Y �����g"S2YH�SBU�<�^��$Yd*{@���Z��� .
@��[����3�f�{�,�z����;����.	c�ˋ쓽�=�E��]�k�~.�(�Zx��͵�ҡR\ϙN�Yn�Hg�]�7G*7��߱CMY�5��E�2W�a�V����+{����ݲ�`��r	��r���_PG#@�o�+d|�'�(��Rw{���X�+RnE̼��%k�Sѐ�ȝ��rh��3��:�_wZޖ�Q+�-��W1;c?�O�ͱ�^F	Za�ۓV��E)@�!��Y_��ļ��ӯ2'ʃ�!Њ�Q���ܠ���5˝��S�SgD�!ug]��[�5��[��y=Z���=p����n��ʢ���}�xO��&�uH�X��!�2S��_뺶�g,�c(�}��d��:5u_�$x>��������:b�ف���6�)�Ɍ_�@��d�I1Z}Zs��YTa���Ն������8n�Ր'�����g0����#���@8i�-���9�	i_����oiLr����"e{i�\���{�$Y�IO��wY���J�S�􊓽��7Am-�ü�j(��-��<�J9���1�Y��N���X��G�~�ѠA=�GL�6��]C�q���|��O���9�̭�H����M���K�Z�ZF�U��/x/�J���[1�'�T09���]Fv�M����S����Q�8���6�#����x����[�b��c-�JDּ1�����R?��.!��$+{�y�zM��k�Ě�R����Q>��q�o?�La��� ��@�#[��ԃg�O��黲��2 O�����Gu���0<��Rv���슷v1���
����Y��I���"N��vD�!�1`�"�ԐP|���{l�oX�r"?tގV�CeQ퐎�y�z)UbL�lt��t������4�Fe7���ɍ�W���'f׉мU遚+���M�$m��O��@w�H?��0���k �;���#����4%�I��P���)pp+&�@����Ku��Wd�6��0�&rUI��	�l���N�mJ���4?+jF{[\�<� ̹�'�{Ɠ�rE���;'�x���&��_ޝ��ͺ聄�� �,wgs�j��.%U��>}�9��ʘ��[�d��1v(Zۋ�p��'+���U��I�����/��n��&�5��dM�g�>o�B,�F��vxvV?�Q)V$�}ׁ�~�'�e�?�%k��(�����L����f�.�T� M[?(��T�M�~֟F�ۂ��u��6/��	"'�{۴�X�.�����SX'�i�bFJ$���U�I0�JP��>�j�J =�K*#�&A'{"�嗷L�����<M���Y���ݩ��~V��' �/}F��?�wAz��x���5�
/9Q�:8��lďm�l�-0�U5<�Fٞ�~gjd(k�ϒ��	4���m��y��n�3�NmRf}�XdڥcjP��-m;��cy�"�R�L���~QB�D=�\E�/<�k��7���.D�#��1�Œ��G��E���ڠ���F�Nm��� *�$>�� ���R�f����]=}:qsX�Y�y����D�7=8��M*�R>'�n��I9}�!X"�N��w%�{���=���-� ���IH��DX��Ac���"�:"���8g��6�H��%����Q�@Ml��R�*)���Rϖ��o<�ǂ?�A�k�/�LB�M��ܖ}~#���-	� ������a����M��r%���_2���y� �[�7Y�����D�B?�Q-�q���A���
=�n��"��o*�`�lX��/��Y$�[���?�Fk�������P��;ع\v<o���!֮=��?�]ϊj���@9�85 �u4� ���k�OƊ�����hƽJ HZ�RTxN�[x�\�&��=,��NpZ���zƘD�ݯ@����ˁ��o�}�w**��Ndb�6�sD��h<��Z�h #�&�C��F���`�v;��۴=o���՘�#�R:��qV=�&i�1�Y۽��~���o%Q��x���W�ӸqRW\��yH���ke	N�����4ˬC��3��(x^�6�{]QePӶ�x�8nm�����4�F�����@-��
z����*Ã�� ׃�4}v��@@ [��(\�ڟ�J�t�߼���1��l�~QM�������F��dU�7wM�c�Y�e$����
2bE!Y?&S1��n8�;˙ڹ�39,� ��R���4Q�y�O���mף/~nf�NSE�B���&ޮ\��e� ��5�ϯa~�ByV�7���;$Or������9uE�����H�b�$xU���ڃ�_�L��ƥ�}'i<���x�_��DL��_���5��V��T'�����[�(�X\�*�N�~���W�81a(�������L��G�]z|<�U��YZ�f���ĺS��'����?=E]%�j�k�����J��9��1�U���*5�]���ɟ���L�̶q9�����9N�f\s�.H��c?k��aP������o��Mܪ+�t�֯�]�o�QgZ1���+~`+ʝ�o��$D���Z������#�Wz���_²�rՁM)�H�����_� V��v���w���NŃ�Ї��I�4�>�@�bX6*D���6��6�q��䭬7�uE���m�}�=�:����;�+�ǒ�|s��LWX��)́v�c�1����E����x��s-�%Ǿ�����[���\9�i��uκ����`����l���a� 8#�e?�}��g*�@3��]V9�r�ޤަ�\��=T4a���\�5�z���q�ϳD�����+7> ��m���J��q����)C=N��n[�{��$eD't�i�0��=�8�x�Ny���o����ʳ4�׆9Q��ֿ��� P|���k��5��-�Վ�7�����*��������֫�΂������?�ٞa�ͣ�v��}��vz91��1o��G�KD��o9�B�#��;3�����6�q�{��g��L&��_s\/:���^-�Fm��e�R�G+<���a��5�ݭ�)�o�Ǫw����z)����#5�Hu�M��)C�x5�_u�}v��_��DϷ�6O�[��O�o@/p]��t������Rܥ����U���:?�m���i��j���i�3����CYϕ4�����`������}�0��AF���׈�f�c��F�2ya���n;S���,g�����trĥ�� �Q
h$yٔ�md��꽬���k-���B�N�+�-\�>'/��t8�2��❗zhu�0�y����&a1��Ic�$Z��P�������A����7dM/��	�(�Q��/J�9z�	�x��g"�o��;}�46��Ӡ��j�]K�^�7�����Hy�E�~g`��pp,� 2>�&�\]<%��+��\ -�4[���)��+͝��v����T�g����ko��?W�1���e⾾:����W�#r2#�3�13��7����8~�W�ϩ8���G�}�!>qI�}�g�c��H�7^{�+u��M����_�=�j��׿���T���<.���fs���}Fv��1�^x�L���q������J;�K]!�v��ĝ��5�v���<��wS��M"1ȟ�y-9��7�dmR&�0��}\	�O'�<�Z4�HX��P�6H*��S(�V��d�!� !P��c�B(J��,�H�i�v���i�nŤ%�2�aP!!��Y����e�|�1w�l����Q�$v.�w��S�z'���RFMcmW*.7&�����4�Y������uʵ?_N�v5�c�.�-����E���Ms�o��B��L��02ks2���}r����G�~��ar���{oS����隫r��R�cM���n�����78�Rt�O|����.�i�W��H�������붅�LL�}�q$���=�1���#�!	l��j��P�`X����TQ��9l�C(E�]˿�ˑ]p�uZ*̨�0A�٦#1�(�q��"'B�n�u��oK����肟@�.?(�W�1_rh��z��t_��2,3��Fd"��q�in~�נ�p��fG���eM�$���AѰ���d��f/T!��E�A�մ��f�g�'$��G~hIQN4�]R|��xYc��f3\�#�jƳR��-�$<��jG) eΰ���bqw�	zN���`}��m�٢#d&�d����ΧJ��<��O^=>ջ<?TtpM���x�~�\Q��+�2	x�Bb���/l}'W3��6s=׼Ǒ�w�C2m��b�ծ���i�(��*MlO�8#'�g��
-v����;���Wl	���i��wU�KU�?qL�#|ɑ-�j��ƿU���$�~�»v�X�U2�~E�jW�}�_�!5S�m,��tX�
^it�,�B�Ɔ_�}��I�"�m���q�ˁǹC��[��H�v&���0��~xBx0����*��[�>~��=>�LWԾ%~����]x�IG�;�>;�Jq��R��O-.��9U���-�YO�[��o|_���5�XC%E��m��e��ܱ{���ke�� ��w��Ȑy����h�Nj�����^Ӂ��XTK7z�н����bt����"V���ߋ���ƙ��F�Z�s�kU"�/Yб�F�y�E�*#�O�6�;��1�-?���D�a���"H����	b�Z�Ŗ�l�ӢK�9��2��yO�l������˿���"�O�p�mH�v$��;�j9Q��y�� �hZt�I+��&��Õ39Z�N��d���vtc9b��%G��i8.f�ܨ~{|y�¹���v'�#�m�67v`�	pVg���Xym?ք�qaQ�Q��K@�.�(`��x=�쟥N�v�0۠��;8;��G������x�O�b���_����+y��q%��X�����wb����)?	\L}M�_;��V�Dt�2�(�l��-�d�mxat2Nޱ�'������ߦB̼,��ӂ���j�<i0"���'���%�������+X�
�`�P+b	:��n��O�ȰV	�"4�.ۅb=�pRNA)���`4CN�����'0��t�/�/A�!���J��g�=�ĤHM���M�[�8���%(��:%Q2�$Lk���}Q��-��}}��܁FO�Mh�'-�@'m�i.+f��+��'k�F	x���wi��x�q>3����"�:cj>�b���,�����ljԻ.j�M�ŋ%/,�	YC�mo��_)���ְ����.���G��L��.8j�̠l�D��9q5r�Wl"ۧ"׹�{����F*c�g�<�q��������Fa�G�iI��<;[i�@x ��^'XB��h�&��[�.�bWJAc8����;j ��C��YA̘��U��榝B�˶1��:qQ�ҿ������ب�%���I�̘���Q1�`G �9��q�b'��bBh��<�{di],fœ�����7b�w��Κ��0;=�1��䜴w����9�O��
S��ʆ���Ϟ�rx����=-�-��t���8��t��h���a��V�\-]QK�L��/�#ǔ	�85�t����^q�Iװ�ƍ����&���%�^�K ^l�<zEjh=wS�b�d�	<�w��m�b��ݜz^�Jk��
�(�|�jpm���H�,+_���]��\��=_�/��ynH���3��5n+�g�G�O�d�����B[��b�/-�i��g�5BH��K���?��y7�8z6�)����WP�܏��;�0*�>Gm�0
(\�����	k��I�&��O~_��1^��R�+L|������US����`�Ӵ���k�C�<�)�~O^i�S�D��6�K�7k�J�@U[	�rc����5�銖���у��#��������3��EUf�űqv�b��
L�,����]@L0�=��������L���*�E�P�,�w��_h���7X4��CI�#�yL�x0�G���t.��L�#v�&ϗ͕fŏ��#��U�jp1�&�"y�:�th��L\��������7�e��H�;v&���f'��݌z͓�l�$tP��p:����k���?jN�FW��@���0r����T��r��L,h��[��.�d�����ўkU�g̷P��(l���oW�r�M�R[�ci`����n��@-�m�\�J��ѣ!˽\����-28a��t{~Y=G�[��L���I�8��m� ��xI��WB�9gg���K<Lie�a߹3�1s*%���u���͚�`��^A��2ğ�������a�o�?�4��Z�	 ��浖+Mӳ��<M���r�6Ťac�'֩	��O�������]}�MI``Z�+�/P�[�W;�qq��;JOW��1>�8(���qM����a���d����(#-���a��O�`d���%��"���e�D���/�K_�,��$6�?e�Ϋ�oT�C
�:J����l=�gh� ��ػE��'a%�Pp�W�Ŗp�0�(~���w7��CS�3�B�������Wչ�]����r<��p���Xf@�zfU$yL�HI�3��{��fx	{o�;�@&y7M�C7B��Լ���([rE��K���L:��'A�e�0�wU���� �©(&��R���ԃ��x��̀��}�ݵ�g�i��<�g?�.�%�GZ�����̥�����ηAP{�c�no�Ī��D���"=�"��(@x@��U�;��CH��@yJ�C��#�3���s/�5�_}��إ�띊CE3vO�g�h�]�å�_w�y;�د���@����j�b�(f�c?E�$�9B��0�� ��[�����79O����%�Mϐ���§�q�d�Oj��l��
�9X>�-�nvD\?\A۴V�b��l��;�a���jI��q|���/9O}�R��Uo�����mf�v�<��̺�6lQ�?\��=zH�YH����]ȶ�qV�A�E�;�����W6p/�ːJt[6�Ϝyn�.v���*�Z���y`�3�J!g���%�L�
�_>�9��~J�|Ƒb���#��ש��AK��#�[2��C��F-��%z%)�%b�O9/����fKC�G	�/ԱS����`N��e��I���6AŬ̱k��LE,:7�>rS�;��ފӼy^�L*�;|���D�Mք�3�_�+á� � �/�4v�ٵRC�bJF�zY5P��/.gN���Q�O|��T5�7-9�P�\mAFԪ���N���Xg���|�8���Ƭ~�? �D*P}Z��z׷�	hڎ�r������&%}�P*�]0�A���]�ִI�ZZ�?�&U;��Wڬ�����ԗ����o�=m�N�L|��V����"��ى�a>U̯��/M�M���;J�NkT�X�]��VC�$�<-'���F�q�+��⵷)hz�yi���N��xX	��:�_ =A�V�h�%�.�7woø7/�d:�w$���Fw��T�|x^p$f%Hh�0���A��(>�_��#q����+��S�ƫ��òt��˂$Pƒa3�⽻�%�ϵ� )�+��}�y��M�r�,�m�[}V�@����1R^�p��엻������I���aa#��S�Z]�� ι�����w�E��G8�?r�e��WA>����Z,�y�������R*x½z�a�ԗ�-�y�5�l$^VvZ<($���R̅��B���!���G_�I���
���{��=�A��x��@�s����+�ٵ ��_sQ�^RM����]SX����NEȚ��ֱi>mC���e,�{d,�iM͉��F�7Y��p�r^v>^y�������Y�o. �>n��Nw��r}�����0��m�	'�߁ �Ap���2�M��ґ�������h����F�H�� ��f{\-��N�|���J,]t���jt��]YQ�?����~�V���"��d�3�kj(�w��?9��)�L����T����."U^���K9���OV������f��W�����H�Bh!�$��@���y�Q��$��S���'K��c��غ�
?U�A��OU��( ���{.�����z�����L<�Vѱ��ŕ�7u��p7Q�+�/[)<�!��"�n��%��j(B/8�mS�[�v
��;^���7�ΙK5R��[S�g��4�U`�_�
*���%j
�d�j]��}�;��
���J~Z�:/=�Z�Q:�#��?s���~a�My�x���f9�
�'.8�ulk���X	�u]Eڄ�m��*��k(5~��9F'�Z���w������������o�]Nw�](+f~���7�ʺ!�˙	~;����հ�/�����[ʗ��_<���Յ-h�KDu�Eӌ��uߘ����gp[�/8��f�fG�Y%��\���&�.�������W�R�3W�dC%��A{Í��"�r$�OG�_�۔��p�r���ޮ0��.��; M��]$v�7uaGL(l4%��5����P8���)�%�[�x
�T�N�{Cg?`���˖��2.�}J��Kyqlb<�A�/����j!6/��.��D�[s���[E�d�A=���$�g��l+C����VGD�O��f}�?
K��c���$őp�����p0��� ��Ӝ��4��9�$�u��N
oݠ�����Fᄦ�u��#�ʀF]^��B���oY?ҩvM�����x����`?�QjP\e#�4vP�b�q������׸� b7��������N)�$���U�T�P����������/���=U��≕~Ͽ����Uw�X��O#�V�A�C��<N%v_F���ʙV�hR��,��#[+n��Y�������>��u��Bڬ�u����p7�K�vu���>����z�\C���%T��W7���C1� X��>�l�� ~���H؜U��U�_�'�ń�q�:^v@�j�{Ir���Pg����1�C�1�z��U�!7�,�)WqVž?�Elk ���i�Id\�kF���
�V�I�z���\R�Bz� ��WE3?߄U��o�"�LƑ�Q|#�z�������ڵ�Q�b���zLkR�;|{�5§�9��L�i@��q۷�)f�����V�a�=�w�_�㲚$�
d�� 3���m���W��*�|�%֖�'!�t�ؖ���Д�(���Y�5
�.�U'd�l�8��n:�k�'B%�*1Z:/k�!γ����6	�Z9�6R�`g`1o|�o\Bq��"����@$�Y�2w�L�֤�I�T:褈�����&�d�J�!�����p�^,/ ���F9�"��E�ҳ��؉���w���Ho�]�4d��_�ܨ{���hBì@Vyu7��9p�&��J�bn��6]�M\rr2��@f�]��y���Xdq�U7��{�6C�B��Jx��s*R7�1F>\�E��=�ʲ��Ws5����Hr_{���?�!�I�w*/���9hS��
֊~i%P}����.688�wpiҺe:W~��u�PIL�� �	���3��-x��M��R[�F�X��Ñ6�#s\� ����
L	�cDhFEr2���;��h��C��1�u�:K����]��4=�9��{���@/zf����#۸<�\*�ǰ���5X:HT�E��w(f������3醪F<�۾l"W���� ��
�w�IJd��S'kn��/u��%�.�-�\�W �+�u(zҺ��� ���sZ���
෾��K.����W��a�uI�w��sq�9<&��/⋂�w�O�E�D����̯��l�(5wa�J}F��/����f�6�M5;�	8�7[�}�˗�l��4��QY^����9r=�#Q��.�b&��3$�y�(1�|}`;8Mӊ�&��YZ�;�$OɛfC��--7���X�qq�e�R���7�z#�p6��#A_{�L�s��ndV �j i�n�� Q�3��WV��*�Rr�pi�ۚ�1@lN����q?nq �rV�RB^���#ۼ:_DK�)��^\z�m�ր~����O)td�F�#��e*X��ug4�@y����H��q���>�j��R_d�]�l<*[�gX"�M�"pfʜG�.�ME��t��1����4�ܪq�J '�x�,���X
y��G��Vo�܈�l���>P��g�x���v+�\��^5�?�]pK�8U�_O�C�\�T���ߍ��O��-�'�9����H��-��@��T#Y��;�c1�Ф��5l)��#�$vzvne��ҠpA��tyP�ڶ��p^���4��&�,�YD��;*��p�d��ۇ���T�D��@�"���{F��5�n�5�h��W�%9��33{+��ci�h�O)/#͋e^��*IrT{O�V�ۿ�|Ml̕y`6�RR�¡�l�����RY#'��;��u�m��
6iq��f����ez!q�ϣO��/�K�����rټ��0��U��!���[-3	��*��l����#ٞM����>�|�j�l��[\�(�
6���G^�2q��SM'p#�)YPIO����x�E����<�}G���K#��-(�ϝ[�ҿ�	+�h������A"�L��;��Vw�zcf!�����P.M˯�-/��_�¬k��z��nG��������=�]���s�CB�+�F�7����<��܆�I����UQM:j�?�y�-C/
d3}2}�"���HWV��,=��SQ�� ���;B}JG�l�Ԏ���]��|�CH�x43���u�??�IM�	"R��"t3�Q,�}�IF)�܀�9�!��o1���I��<�礻�uT�_����V�=X�״���v{醴,��x"�9_��"�4�4�q��p��EJC"5Ӛsc��Z���5���{k��e��h�x��[�x�R,}�I_�31||�徝&�Q�����[)�z���ϊ�rg#�CT/��D�V����(�]��dI3!׵��S��qhʎ4�Z&��a�D���P�l��Cx��S�3M����q��%RH}��)V&tT��M�.�W���a�D��.Z�ͽ���o���C����(m4y���hi�s�,x��Y�N��fͯI�"F��T����<Bn�J.�!҃VB�Q:+jz9�A�p���)O��yn9I<��-
��yv�x�B����� ��x�₦��4[KM�i�x�w��<Q��$h�t �iP,uA����衯��~r�ĦU��I�|��֚�ڭ4�Q����Hۀy��'�v�; �����B��d�p���D'QE)�n҂i�r���탺�Aa~���<�^KL��b�F�9����!j�qNĴ��u��Rx��dܢ�[���'|ڸD��{�+�Y|G���O3�L��2��b[!�i��Q�!IE3�h=�T�X��ȯ�d���jlX�H/��^�%z��ѝa�����U�9�n�����c!�{�_�}�yڞ�%��!;tF�@�]�%�=����P��Y"��r�rV��C�o�?a�i�CS6x����b�rw�s!����-�"8����q��UW`v��9��݄y�l�Y:e�J����KV�t"�)��RPU�[+��G*�ǘ����?t��8F"����pgO^�B(����mG�9�p��n(G�+E�]�3HxKe��zޒ_�e�ph5b���IAj����������-X)�hŇݯ2���;��bɗJ���&.zRiXh��=�2�M�����N�I��&ҩҏ�j6I����B�澢��I>�>A�/�k�Xe;�Œ�v]>�p�J�Ʌ�:Q=��{��s�%e�.W�f������fy�r�) T�O9�|U{{�L*��'
\�W)+`�\�[o��W	��V�]gr�zw���x3�P���J��j��'總ß}s�`���ۅ�}}��+nנE�RƆvE�v�f|��~���[��7VT��s-���hğ{��G.�=5�X�唿��\I�W}$��2�1�"�+���������׷�Q�9�Owb�!�~//5AJTג����$�C�Y��:(�������up����y�E i
�s��:��,��s�Q��G�����z�Xd�Ɇ�:��MK\{����_�_��ZݽO/��JI�uw�����-��I���|ô���SΚP��:�ŋ�������c{^��mh�%wB��d*�`$�r�$�A��]V�i����o��BQ̯��B�Kc��˵W�#R��$�a,+���wJ́O�N��l�Ì);�F��^e�g�Q�J�h��t�Rk4��3���t�x`M2�fL�su��x�U�X�C�<9P&�q�+kt�$S~���dJ���PK����Р"�a)���`���Y���g-�ڦr��a������4����%���_���}#g����F��_���`��h-7�"����:��1"�։��%�,���L&Ť�Ԗ�6$+y�w���7h��i�3���z\}�����%�Ұ�IɅR#�֠�x)�����JP_@�T���4����z���n)/��MP/���?�]�J�m�x�r�c"�'�%���w���R6��Advex�/X���|[��s���T�g[�	�6r˷����HG�=�O���­�Y�X��oYE��[$��9X�RA���wԓ�ʶ�s�i���_�M@��	�����N%'��Sb �w�l4�P�لA�~�����K���i�9ʅN�\�sS�j`_��h�	�_���q��ͭ6��������7�&�xu!6�E{N�+�8Ժ�~t*���]<�����F�Ӳk�D�쮘�8`'Ryy҆E�h�cK���b �[VJ��H(լ����Ra�]�E�M��J@,���%>ӗy���k{��y�(fc-'��*&_F~�8�O�x�&Y�Mɕ�6���=j���q�1cw� 0PLUz� ���@�<��;6@�YG�Y����+���{�58�V_Y�0kD�|�����28k}�aQ順ş4�VIŽvw��Nޟ�Vs����.`�FO�G�x͘��W���Θ3��~�� <l�����!��og��P��Vˡ��>{61C��V��P�����K o���cE�Jr|@���y	g�f4��{��jgВ�c�Qǖ%׸?������/
���1�ݓ��W�����fF�H������އ��<�����6�28���?����W����s�����Z�l�?�n�P�S���<��w��-���>_�2�ـ}(�@�p̬��[aC�!̟D��>��|����b���vi������[�ݾD�U��\{��F�B{�LA'�¦�L���-�Cq�@��Г���0eM$�z�s(���IV��r=~=��G�5�	1�����!/&ym}�����~2����1�z#0��R��"��>��[=�����F�)6��Č�gZ��B�yB�π��Q<O7z?������WN���h-�{�]`���O�Zf6{�qJ��0�E�L���`>w([�dY����ǐa�9�M�,-�3��|�G�ꟙn����"�& �����v�L|C!]���T
�N����6ӛ-	��R��m�9��-��R��>^_���!� !�ȗ��?殐���3�-������Q����ʳH�1��U��o��k2aMhLNX<�Ζ�-��+Ɵp��c,:Y��:垷$Ҏ-��*MP���k�9��w#b|3���b���c�F-�w<E�a���d4�oMf�!b�r�{�rtM+A�Gљ$xL�����msP�b\8�O���Sp�m�R�E9���Oav01�am�zY�eg�K�6ށ��9��(S�h�-�D�`/�2�s������`�G�AUide|�5B�k����NU��=�_C����C�g�1Pz��Z� [��pU�����ST�?�o�C�!��.D�F�=]�7�-VX���맒?�R|W��z�a�����is[<�#M�)צv�-�%>�y�k�٠v��/��Z2�![����I��	1f���b8��|�Q�wՐ�/v1�7�9yq����eeW��xd�h��D\9��~�u*���~��%A����nO[y���i��t�-�:�U4R�\R�*�9v��Tv�Y:��f۴2���cq�$�Ul+����>���jE_v���Դ��[����Q�.���g_<̖�e��9�ν���}�V�X���쐩|!Q�r��B�F_9�Ծ箺ǣ���AΙf��g�Ƌ��Xa����DhK%%=2	e�v�ufq�������j,^h���N����~0^�3���]��3�䁳k�G���l�d9�{��=]l�����D�F�r*��F)�����5�����ܣ������Q����g�����8��s�@H�!:D(md�9���ny�l�����+ַ/ �2�ުt����<�W��Đt��Ƽ��	�������N*�q
����������ތu`��a�N����-��U*065&Lt�,�E�yR��/��GBVp] O.q��ڻ��?.�M�ܝ�jB}\!�Pj�݉���|�bKsLK�F�B�6�'�#2}�Y���{���M��?�}<��ߞ������lDr�������8��I.uJ�9b������)ʾ��ԄϮ�?��q�:)����ǟ��7*
ͮ��8�E�.��ݵ�_nR�^������T��ڌ�7Z,���7gNV���*F^�\���/���A?|�_�������eO�
Hڎƽ&S�,����>Y��	btv�i)���tÛ���g���Ew�b�k��}!��=����{�g�<��:=E��&���7�����(����/<�W�5�(K��!X|ę�p$���ɻ�'� \�QG�������VkA4Q������A��2��1�~_J��R�ݠ'�n�PsEi"B�:qn�->!|�O�^��a��ꤞ���N0�3�?��A�L'M��Z��i�h9U�:b���x��h"�����U�i}�zK��g�zK\3E�Q�f���O�9w���Rڌb�1���;
���4^�q���3^�v�Rn�^Y~z(�d���(��GYֹ;�e\}c��:?��$�EyhֺF�㾚�B�9�Q>�����bď�g+�$�<
9���uV�腤.�1ʙ�i�m�x����|���j S�B��*�Bʨ#0��ؽ4��{ BRo�8�6`�ú��;��iZ�Fc���'!.sr���R�XJl����8#��w��2�BMUSxG�É��>y�;�K'A��+�_��� `x0OI2��z~�6p�~<�ꋦ��y+����h�&���)*zAK i���f%���2����9�����h�]xbT�`H��w<�ׁ�^x	������g�/��߈*���5sHa��A�����a&��{&�vm���g&	i�#7ĔD�����6�s�ZU�:y�V�o�U� �,�-�ts��|#\�U�ۿ~���cs�x/#�a�8�d4�o7S�,a0�?jv/ah���~3=�7�l*�p�W���*jW妑T<1��>�%<��Re.��.eCE�g9��u�m�4v��Hf����ZꞭ���TT�:>� �g&$%��v>��m�J��d��_����ɓo��y���v��_������ �k�����%!/y��	�'�LBD��$D�K�jݙ�6�?[�s+����fG'^֝�|��-|R����K��I�ЃmxY��j���w�:`��u���:����!�]�V��>OAژ*���s���zib�P'�2M�X��7��G���5�F.s]�i�n�@���mc W9.Fd��p��vv�ۛ�vJ�V����=xo� *tR��3){V�ߦs0�EYR�}ڟ{�I��o8w��������0��9+�S�'//vE��*�ެߪ�Ѣ�AK|7�!?�kM��Z �KU�\����>�-�:�3]���\Jb,[��NR]>�I9���7$q_<PG|Iڶ��,,:vW��9ğ�A~]|;;�(&Ք=���D�m��4������d7�ш��l�+�mN2c年׍�=@�e�,�K��Y����_Wht=����j�PpRm ��U���dRR�U����Nxn��KUD�p���5��2�7�d~0\�$v���;k	r�A�p@�6`�?e���T�e&����ׇ䗕�c*`��G��A�}��̙.�Y���0�e��ι;M����|�V5��뢨9+��f��!y�ң����C�Ào�]��?7�5�`�gR��b�g�R{���ФE��r�`�- � ԡ�8{��U"�]��+�߿٣���x�"fi��Z�E0o�Fy�i�i�����͋���g*cO�9#/��>|�c�έvm�������T�Zy����we�E.Oyt�5��q�V+����]��׋y+��,���y��u(�0:��`=�V��s� 
�/o���vδb����karM�Ơl0���;Cy8@em�W��_�$�)2�`�����IW=6Y#;�V��udv@Ш��v�"�V]�aq߇�A�M�1$>����Ck���&=�E3�줍��9#�fG�\��]��ihQb�_��>`��f:Ն>-!���j��ߦ
�~LT�zk�Sc�����#���_n�7Ħ's¾W�Ѱu+�-fV6(�3�L(�GV�.�R/��S[��/���`��AǤߟڃ���j~)���<@��� ��쬉�N���k�=�Y"�-j����;���Ф�re�lWL"܁�(1�-6���^&�#g�/�%���4)ǧ����zJp�*�+"��)�ޥh����L��&k5�R�k����Y�q�Y?dS������褽E���a�����EJ��AY���>�3������g�=�Ǽ\)!�nv�ub��Wx|˫���,�tf�}���8�`#����@�B,8|�S�v�sku��9Ǌܫ�P���h����$m^��3���z��#i�?����ea]0� 1o�^�	o0%��D�G�(�#�(]^oТ�+Ƅ���7;�v�nt����`z�
��_��rL��ú5���;��ג�ܵ�>�;��k^�����Sљ�)�����aDi���`t��_˲�>e��z껚������,���K��b	�SZWrg<�c>�����<<����Ӣf.=���eN�����PK   �cW>R���5 �= /   images/e1c0e916-28de-44d8-b600-7ef9d9f2b881.png�{�_T���.RJH#|���ED�T:Eʥ���DI��F�n��Pb饻Xzaa���������yr��9�������JE�B  �^�z�  On/2��;���  E�����kee.-7g{k �'->�TKא	��lS�g�"o}��&�E����V�,(��GW 28��Q�H#h2��N��k���?�C��x؃�K�)�=���̹�瞺s �ir�����=o�00����	@c9�2�f
[���^�,�C%a=��Ň�k\[D(i�@�,��m:�zbv�;��j�k^^a�+U��&���{���ߟrφ�ދ"���}�-t��W.�3�ɽʧ�_�UIv�}zUAd���z�T��P��e��S<l�������U^A7�{�k�Q_u<b�|��w�T�."�5z{���ߟ�^��ѫ�r�آ�$�w}/��2*�C�_@�ܢE�܉�ݴ��6����$�1�u��t�֡�D��n{Z�kS@"��L�����1gKZ7-��Nn�K{*��E���+q�t�j�1�ޜN_L����V�����s1���W	�d�0�y�OmY��v	�k�s�1B���9��9���*�4�G��@ҏ�_�r9�kd�kQΡ?1��=�~F�l"���plar;�Ko�vf��I&V�1�D��:��Fؕ0�	�rʨK�{��ҹxb��瘓�Fd�#0� �1T����*�=W��!%�3v��ni���Y]���Y0��c)��d�[&9"�a�`���紡!��T��'\V}w���񭑆����� ��^��O��ߑ��d�g��ݢ'���Vڢ:a~��1�����j x��1�(�粐�H(����ʟ�)х\j�` ��D�~�:���g��P�����3������}�'Pm��V���8��=�Ȃ�d;�YZ�����a��p���CY�D�|���l�����w��E��꡷�'V�t/)2�9)` "��ߞ���"hJ����_�z6l�+f�E�m�!S�겛�J�^�rCu�qC���yyx}����� �-�6�$�R�ɫE�C$��_	d�6�R���:�����9�b?��LޖpIЊ��[���?���"�_��{�-��O�י}E)���e
���2y�����;���We�6�|�_�z�[���<NOཀ����_�-	=A�wC�"�
�ʾ_ԲR���qx��F������y�[�K����a���z�?��iE_�2�@�Z��;�
,6�V��k�k�5�52	Nj�����']'؊���\������j�>��DXv.=ef���<�ؑ�q������
�Ұ<}�"�����-� ~"�{6�L�^�0�lh78aTR��ʙ����a�b�}3�E6���-CM!/T��@�9զ��C�D��ƒ�#����S2
3^9G.�2���<TbQ�4������9�=U�zC�s���]*�ϯ?ߙ�}e�*,Y$�g��s�}����->|�kU5�7����� ��f��;s�@�PI�n��d�u�|쪀�a����֮]w�<���kvS�&o���U�l�V1�>B-!S,�?�Z�;����=\���6|PҘo�cZG��n/x�b�hoa�x�x�x-��vŮ']#��U�A/���#=�e��8���6ܙ[�����c��k�#r�ª��ԫ��P�&���;8-ܻ�k�|_o�~�t>�$�7��Y/3<�a>�s;y�qVw?�}\t��%|Pv�a�Z�;>U�� �S��Wp�����׆��� �� �+���8.�0� �8��	�EK���Q���2Wb��^��җ�K��~��>�͚N�UL��S�+��uS�W�~J�Oq�)��45WԈ���L�~1�ͨ��ù}����e�a�P����_���I��Ť���%ow#���F�9	>&���W}rm�ƛ���gm���`^�2�q�$��	��J�J����b����}�[��pZ��c����Y��O�G�J����k�O��|4>�q�w�J娍����w�i��/�zF�FY�0�3�u�<s�8m��������?�".D�0i�<MYe���������d**�8����d�J�]D�O�5>۠��D�p�y�LJԼ�śҝ?��O�c�}��M�bEJ���3q�51z�O�������僥p,w>��Hk�>�8��[Y=��9����wBgv�hTu�*�����ִB���vrY� �x��Xa��%�����?�ba�&�1�csid����P��˹����~�M;�@W�D�⽋��X�����������,E�E�Ŋhƽ��{��{�
�E���l/s0�W��2�⺚3T�a�E�ឧ��'i-�ӯp��iH�g���E=�}W�˗V�t./�ֺE��<8�f��<K������R�
��v
%4$��T�5�7ּ��C]�b�4��\>�LM�T�l���y�/6?;x�&��>++Jb���?F��;�ϑ�i���v���X|��^�y>�]/}(����S͜G��x1j@��x��r�ٜ���nn�m�����N��2�!s��4ǜ��r
"�9����E�����Vx+2�t��P=�4�Rfjg��lQ���|<؈�Ś���P3�~m��۔���q����k�(��y�u¿���\���;��Bl �ů��v����X&�K�����O׵����V�VVw3�$G(���x�6��8)��$�k(u���(�4�� ӧj3��p�A�����(��P2`^>L�em������8�^V�6�����j���R~9G]��j�w(����QpC  ^�Pz�c��#o(��I�����~}E������(4cNB�]<f�J�����$�)���r�o�b�K�E�(���+���$�&}�.�2�t>V�q����С�́�L\�F�^�U��U���N�'�����?�����?�.��5�*�e!���Ek����8��y�	�
�R���ҵ��B�ɦ#����N'�1��Yꖳ0�q�3+uފ�w�;!��V6n�q3�0�9v�~1�������7���+��k��/�z�ڈn�K'�� ��B��L_�<�#vj9�	)k�)Rv�_l(��������
p0X'��>_%ݫ�u��a�rS9|���s�z13���UOg���(f�I�T�X�a��鞓��.��RgSVm�O��4�4���HO�s-е����#P�mǉmW��ڮO���'�WV�R�_U�M�`��C>[��ĿhL#�]9�k�ykd����鲩��z��~3z���2��ۥ��y�]�P�,ϼZ�3�w2�&�A�=A�_	؇��Fv�������	�˝��/g,�k2���+������a�n�@�Q�K�(�+���ק:,8Ts�O��fQ��s+�P�@o����j�n�Q\�"��td�	�)gs�c��j�!�!���q��ki=��SB�o<U%��y0Qp�p��c8n�9�%���R�s�]�����6,R{_��qO>]�°���#7}7�1ɔ"K=8�"~dO=�R��6�zK���la/��|�^+ ���Ѽ��?�:ĥ9/��yM{&*&���J���3q�ހ4��v3�I�[���N�7�82�?Q�o_lf���t/��IL�5�^�����n���&�l
۽��%���<j�_����Q�eJ�/�M��^�,�/�&0� �~�Jc�J���J����\DO�+���_�_�AF�fF�s�Z�Fo|V��/ޥ�����p����� �ʇ ��T��+�d�ˋRE�`dhA���"ط�O��7Ea[f�(<�C�%����кkA��!��@?%��v��S[�_Vgedݖ�]�j71y�۲�+h��s��U8��i�::mޭҟ?ރhDo��_'\���\uu�gw��M�d�g�*2F�qj閐j<�<������,菑���iݵ�`
��pۅ�����t�tc�,B��/AT/��h,ˤ��v�L]�ʿ��"�_����o�.��c-?��2�66����
`͙�bOC�G�����U�_�����hx���=���K�J�"n;� mSn�]���,u���9�I��(�S*U�7��d�J����j�Yu��ӒCNr���۪�@�B�z:7V^��[$\t	�İ�mX��1{�O����3�g���m� GwV�|�>:��z0��q�Ǉ[��"��zA��4�űQx����O)�\�t�C1W'7W\ǆ@M�u��+�XΛ3:�>��0�� Pk;/b��S=�<G
�.�3�z��~\Y�����~�C�,�@��U]�HY�,u2�45�1gCTnPp������Um.�Y��4�Lo̼w ڱ~�l�gՙWlҊ�o���ˡ��)��CI������v�[�� xx��M�]ך���3ӻ�����fGR��M.]�-��.h�����Hcw�j�*+�/�n�H�y�m�D�!}<�eGs��w�?;mF�dbT�!����F�-�ydx�"����s��Ub���>V�[Ц�B����ݙ
��a`�&����o0�_�BD?F�L��b����|Uּ?8���\���8\�YT֫��c�у6>�-�j���f}��ƿ��n ������+sL�K=�+S��^n�4�qI�9������Y�'��*�h1��=z��L�X��� <��C}��Ju�E=_�����l�F󋬩
������h5t��h��D({���}~;�+��FwL�O�q4B��v��	��k���ϗ�b_"�Ag⯊!Ϯ������[��\]V].��i�!ŕH󫕧��{�D>�P�_�\�CK&}ɲ���3Ө�����L��[�ٔ 6���2���nA"�$�,Q!w 4qe�<��_�)�w#���F�/�(#�Q�����BI'�Q�c����gc�{��7.�s�_���E�<[�<� �M���o�1��T�ne�N�R`+֒�@<��ݛ���ዬ����� Ҁ�iD��s�
Cy��ܡ<K�j
�(�m�u桘e���r"Ed�V9��+5�c���
��A�bs�D��"�G�������l�d� iȾ
5�R�O
�~Y���,�~�.�X��L8���d+^Wx����B�g���؏�IL�i����D���g���`�e��AU��-���O-���@)}(���c��ب)��Yt�11�_�:�ρ��zX��(9���:�#��з�o:�dC�>�1 �����������B�W}]�NΩ�&���&���<tVY��
�;��u��"���1�孺��7gs�-�%��y�!60��[g_��Z1s��b�_�M��\��k,���Qk+F?��߰��A_�(ML�'>�ݤ4�E�)���E��8>,�ԮK���n��_6�]���*^g�k�K�!~ys�O_�?��r��}Vrģp�WӌVɹ<j��������9� �􇷶E��`�w~ɺF�K�1���s�(	p6�Մ���[Rަ��t�(��?�\��O��b:������lPèdwB5�
>�!����qm��<���^z���a�Dr2W5�R?z!sQE@���օ�U�v�.�=*~�)�}�Op&L�C����H�X�P��]	�}'s�N��|�w$��N뜙(B���/��p��{����;Q�b�M��X�y�����?����X�<����s�EPb5�My�7�N'�-�x���R�4r����3��<�p�����M���m,�r<�m�t�6R�0�2��hW�v��M='0�i��'UUz�w�W'���� �k'�R����;�>��z���8>qT��s`�W��yf_�]���9�dп(�8zFbTy&��(�S�ژ�kd��ۜ�d�R4��_�`+��_j� ���oMvF��w���$��	����)ݷZox��lY�	z���x��E2�w�����ݶ���҈dK�A�Q�o�>Ҁ��h�+��1C�c_aQ܃*t�xVd�L�v&��� P1r��hg�Dv;�Kϯ�OZ~Ϥ�̄j^��f��\q2�?�-���#�ob[d�����@_JUG}�$�Cpd����d�)4ؚ��]\�5���6%���eO�Ű/ٴ�os���(c�����ْ��/�ww;�>מ��V�G]du�d)8B*��|x�)3v��%�Y�ɛ>���Y@	1�]��S�sw���i�Ҫ�G�Jܓ���ӊ��D�8���g���% &~WL�%N�LT��z(X;|C=|_̭��[� �U ΰ���~o����V�^O��vhH��Y�(
Z�?���9���� ����2�fdW���I{,\�'۬�-��.������[�6K|V����k�mv�};%)'&����V���xL`��s٫���C%$�ұݥ� ��bD5e��\'|�e(���U?�����U+э�=�P�=re�Z}+�V3����<��^��\�-F����8�/�)E"��~.�]�F�\?w.3��w���Y: ���\�x�u�e���1�pE���Ć��+�4�'��i&�&�Qg���ڼXn{���&�g�\^��N��Z�o`<ݸ]�jFo�A��h���0��l�������̲а0�{ҩ�U��Q�a�IOZl����l�z%̔n���͔��u��rͶQK^q�2�"�n�)��#�bIA�� ���b�ԸO��j4�x�
� �������n܃����W-�
ʩI�����Mn��[i^���V���l�U�ўRmR�J������/]�u�Na@�A�j��;��˶���bl=�ت��ߩC	��S|�>�V�P� >m/����>��r��w:��яr���.Z������.�܌gy������;��`�qy����6�W�P�c�9`Un](EbG�[���O1a�&C�������#����b:e�*���U[��
�=�r�{�5s'0,����_���W����k*��n���֠b���?���î5Tb��L�e/"h8����p^�n9}���=��!X� ,�w�m�\�2�U6�x�-#J�H�E�g��x?u��o�.3CK�xm�/��1&�(^�ף9���r|����r�5fj��A#���+}���nM�ɨz���l���M3�&��ٞ���Nkϙ�h(L�rr����kou�ܧYB��c6��c{~���I�BE�C�4��$����@(;�K�3Z\��Ϯc[V"�|P������o����C����-X��u���ރ9B�Z�\	L�/�bݤ)�r��jt��Qo���z:C�Xw�]v�l��k����^d�u,�kׅ��f	����
�@.�m����>+_�3ik��IΝ��؟e�)�?��]M
�;2Z������J�l�o���g��e���83x��h��\w�;�A���=O�H�Ψ��~wv�U���EGŵ�(y�0��t���7
A������չŵ�L�o�p�C�������V��X9 :F���������=��l2��5��|��^| K��|_?S� r�@6 xD�~�t�	�w̷��z�~�\[K'.��#M������T͂1�$�p�<r�X��$�����4�
l�w���@��J�Y���ŭ�lnY�N�pе� ��
�yk��������"�9>';��F��j�;$��T�`�m4"�T�[!u	\�&���
ԋÌ�җ_�kX���2��X�ą"bZB���RW���G��$G���+J�L�}]�B���!]�U0)K����u��;���~��>���@�-��2��V��!e�`c�{�@/�˹6}���W�8�-F�(?��l 7*n�0Oh�Fd~� �i�N����m�[�7�J��;����)���A^V�di�)�n�}���ͬ)��	�?�-@u�3mY��bv��m'O�Ւ��JXC�:W�mv�H�ɷY����e�ԻM}	G��J
I���yj����w\��5�}i�5m���4��%Y5�F�K�������» �:q�T�ww+�7	�:���0�䴈�Rc���t�2	O���N�����1~�sRI���E.�_!	�=_�n�Q�ך�^�+�\F)r�XLJT����2��0�7����xcpTM�"'$tm�����[ͦ�_������𠗨��J��U�'Т�R���ť~����g:$k���a�����7�����'n�^�lQc8����7��L�63������p��m&����,��-&��&��$��Vאd�j¼+�/��-H�`؄&�^'Ng�ou-�}	c(�|���Q_������94�x���_��8��0���as�
!�Q47������r,�̣8ђ\�K���*_���80O4�ZQvbl���e�֏U8�
�T��1�&^�
Q���x	���l�	�~�����-��sL� 4t�u���2?j�tz��$�RAq��ΖA��@�d�so����.�_c���6���p�v�GN�~Nǭ��
�"�2���o~�Q)�{�Y>]����F;oU<75���*�_A�4��
b��ߤږ�*�n�	�e��rb��%[��n����SZ��X������\k_���^�q��)�5e�'V����	�R�w;�}�Ki+�� +�4�jt�\+yf��I�a�_m U7W�}�Ŷζ�}���2��<wv����$��!+��$��(:M�ݗ�������h�3��̦@i2������.�Cs��Dd�4~~JG<��h9�Iם7��IU�p�rLϚ��N`*!K�gf5�¾�ἱH��j�W ?Q��ސ��>;ڧ��j^�hX�	�-6�e��'��
�/����25�L�	��bJ�§b�eًS=�H=_�[�,��_$�yn�M=Q�uu��>��f�Z�͸,�@mK��d9G���6f9%��a���� �g!�>~de���8��*�:�x�Q!`!�r�ťF�����x$�4YA;�0k�>�PCh�h��̕x^<����'q����~�W�)p�z-r?$Ϋ���]�&S��|��'ٛ��:mU���N�[Ͼg�� l�t0jEڭ�E�䗡����N�];��"�J�������3E�.{6-�c����j� S�&�:�V��b5櫤�l�.���5���[�E�k�)	K4ȗ=>HAT�F�֮��(?�u^l2� S)�ə���r���J�uCIǏ�w�h��H���
m��<�)��C<1�>�]�h����VӲW���;>��֧؝6BDD�G:~��#2���5�H��a9�d^��N;��.���á�� F���Va�+��p���>��R*=�	��[&ؠ�%�ā���Y��WZ��#�R?���B[6�4��A��v���x�sL�q�'������ y!"Ӿ!��ٷ�4��χ��(:G�}[w2x�������uT���ē�A��P�/�q�@����[U�3���M)�u�ߘ�wh��f*��P��3�%�~ʬ��"e�>�	C��	/(��b���8b�B�����2�: M;�&�;���+ކkE�}>�i�қ��7N��j������Or�/ڒ9�����Y�x����7V�v��\��kAt�ꭞ��g�2�5Y��ʱ<?�.�b��Ɯ��V�hVUN���K-�vq	�\�a�o��^Z�X��=:�(�T&$u��:�{/�/���"?)�nO���0��l�ք� �T�OxՕ��POo��c=ߪ�x}��z�r;���܏?�/���=gܱs������V�l���'4A�����?8�t��_��sl�V�xk���Q>���#�F��I�1�W���ӣ��J��	>�I�&��["_���V���lSa��<��+�:y7os�iK��!�ѯ��F��sJ��`b~�b�K�p��I>نI�7q�o2������`d}�C�&���o��b*�L�b�"ewU\{-nJ�>̔G�����:V�buh���X��)��$'� g�`��V�$-�fV"��Q��b�W$;��}r��*.}�)�0gl��%v��/�蟊�i*&�����:z��~��4�9�u&��4�����~�>cp�@�6幄`z�b����&�7t4����J0�0�$U�)��#P&�E�4�P$=�g���������o&p��������I��Y�]�-Ʌ|����H�Cm�ȡ�OR�[����J,g.{A���9A�`��\~͋\El.gT�H]��th���'ƆdG�6����$+F�b�G�Q�� ����̙��ѡ��uD^u���㑪H���w~e5�*���P��L�#@4/��ku���Cus6!�=:&�)��\��vF~J�F0@�e���/l�f�;�k�W�u�Ue�*���rj-B�lHO�^]���H�K�H�]"���3^�� G��]]!3�^�¨�Үx�Һ��3G����ͪ|i7�����#�l�ݸ^i���X�C�j`ߝ-i_jއ~#G��M�]�¸��j&��U�0KGSۆ����*���7����q� y�+� [vp��&�?Od�1�O��.��6�*�!4�>yR/pۚt��&��h������]O|�a���$��Y���0�]�&��ֹ�XT�E�٣���q�+҃��Q@��d�s�y��������R��o�����ʸ̝Q��|����?|D��c@w���~�?;f������yl�����[�q*v��2�0�}�l��3���&!;���\�kN���z����>�I��wR�	'�WAn����P0���*���ےy�6��K��u��-����,] ��x{=ؿ�mes����D]�F���O���2�_�
��	�St
�M��l(��yE���XK�B{���.����ў�L,1��'�/O��k�0w�� ��/�/��t2pEw��E
'�H���
�׾��t�uR��2&��JV��7ͨ��?$ۂ��4���r��L��q]���� t�^���)���ɴ��P��(u��Uj�E*"�P�_��������>�7��&VO�Ш����c�R<�\`t��O����&و���?!t�;��O��^�e��s��!����M��9�bF��G���G�'��Gx�jָ�n�j#�`�^
s���T��3j�b�Çi����Z���l�W�x0�z���+1��Y�N<B����5J�9U�9�AףR%+�\4@�5V�����-<A��.s��]�c�Y�"�w b���7^��=D���`��RoOo%JS.��Q��z�k,h�'Mz2 �g�0�3�^;���b��^�pJlm�_)�J���𛎶2���+>��p���Za�Mi���c6'}�ǿ�M��[>�K����lRgŕ>��#��1ըr���Ł_�s�_�N�WRW��V7�6U	� �ԯ�h�»��5X�d!#������X��fs{q��\^�(n-�Һ |��"l��;�7o+���Q_](�ȟ�dxܐn[8/e�2V���Od��ΓmY�($:h�06B�z�bC���nd�Ŷ˯��)0h��;O߸+/K}���W<NFuϣ��F)Zȃ����D��G͆����W��K�b|�
\�O�P1��c��/�Q�;��AZV(�F^�n�EtE���3�wc�~=�x�����Ikv����G�J �Vm�m@	��li����-� q1�at�kd����*�5�Q�4�byKgr��(]��П,/UEo�e��:=%�c[���>��"9��&	KW��>�:�+v|�&a��v4~�@��\ƭ��7�oOӜ���зc]��صp5Bt�d��
�tD��^�8Q�
k�iiֻ��D?՛-�7ǎ&RG�����d�V�]IN��9��Դ��I�*�����$�t�w4(���x2XQU����Ha�T�����m��:ta'����~�4:�á?��x�F)�ֵ,:�����av��]���8@�m3)&���-�j��s�g�;�ٹ��p�׌}�xy�x����w+���6>���w ��lR�d�Y�%����;�*��jI ������@�It�y��\�X�{x�W"6,�K�Y�H�l�T����
ݠ�l�y� ��#�:���v�t���Q�J9���K��bi�A}L��gj��ƣ՗��uv=�~:�.��RB/��Q����BjJ�r��F�KN�����Rv��Z{�yU�������"$h�xY����1�AJ��`'r_���S��7�ę��z��� ��UM��N*?ߓ����)�w��!�Y��mHF�2ZQt�X�Br���s��oeM��TM&�&�%F������>H���6�#h�=��q[N�$Mɾr1�igB��d�|^�����0�X�4�f- �v�7{�-�p��j������i�����+#P�Ƿ!=����ꚧ�W.,�N;*��Oҏ��/v�o�c 4:�*�jg:����y��4U_�tEƅ��3�?@�L���������Ťպ��I��$GaS�=%�r��q&��k�B8Q���CV8ȴZ��1���u-x`�}�ո��?7�Ѣ���V	�Of���ѥ�=Rb���ӳ��!������8!	���2�5Y��lO�<K���_�i�jʴV��v*l*L׸��(��	���-J�">��X��:���T�1�G*J/V�$/'��)��!��-����!'>��ps� Y ��p����i�Ĝ�dn�Z9h|�W��m��00�A�R�Lgx��E�����N@���$OhE�U"Cd��@TBD�B1	��U��ہ(�8�;S�(�Pz��o!zP~cF�L��� G�+�H�px��G6;��p��,��wx}i�,�g�� ��ghi��̓&ь��:V��Xm��)�E/,�~�����"xU`����"�|��v �&G������d*W�W������B��V�Y�s���^�4���Pi\������m/)�R(�	mA=��p4s�/�ݡ�ƍ�F� ���oA�rfx�O>=Gʚ��G�T84Z�5v>�������Ho~UM�s.M���"�[)	ִ��� p��ڳ��Z9�Ƙ;~���{,3�JM�X���Ǌ����+q~�T�Ś����ⅵ�όl�~�^`º����W�4���;>m��8���o��X!W�p��ps�y��o��|��8�1����������ڄQ�q��sq�&�/R�'έɔ�tQ��/
��Ϸ�7��+4v�)�(o귯^��v��5�����;���o4X��z�C�3�c#axp��Jb1�8М%���"J���?3��J�}s�<�o+��֧^IR*��eS��)��3^��]8)������cv�X�sx� I�#p��{��{E�3��PK�u	��d�쪖���2��wB�oʚ�J��է��|װFݷ����X�R¦����}D� 9`�~�K���i�>;<�d��xc�X���	����k���w�ɼne��u~�;�5��>��6��]Fc7��x�֣_�������8��$�4mm^5���l��XTWI��S\+�r_�cf�edo���=�h��g�k��N��	��-o?�b�'�yT�X�n�;O�h�cT���T���Ü�ُ)������n<p��}�����˿�w����Tu���.�%��|')�xҍ����b�9������>3�w���� �Y_t�o�H�S∜�M�|vU�J�7F ��i��a��p�kF*�5k�XX��I���Hn��� �عL�߈�f��Y����1@��V���v��)���<���MB�Rg�/Ǡ��E�U%u�n�Ծ�a�����jA��[�iV�C���|�K9���2�e\E�/y_�#�BI ���t�F����J�����������;��z �ȍ����,L	�I]��/�h��%Som{��+c����X
9�˹�Zo�΄�զL+xC|���1�ϯ|�&@[ݳ�i!V��9$�EW3�+�Nr� �a���9+}�عn��׋�]��HO���Kcm.��U��n�����N�b"OkC�G����\?�r���P����!o��`<;�>��.Nv���e$n�'uը��b�+���!��h	R޻:��~Y���h�k����Mp���c!u-<}*6��<h�6� 
���l��2t���>�} %�f:2 �`�U8hU������k����C1��vh�A\�/���z֬��?}8����a6Yo���ST±���Nd]5S�̴7�O&ݽ�_ã���2]!�;���y��G�����R�Q<��a�姭M�}���7�D���%$��g)�]�Lٲ����A�S،��e�ZT;@�Ekے�8y=֓�R� �9P��ܝ��$�vgˇ�>���mX����q�	��M��~�w���-w������0,����ޥ��"F`��� ^�w��Q�|g5�8LŔ(��g�\}��S{�W379�1�%�����f�Ng�]7I��$/�)J��n$�C��N�0�)_�������sQ�h���$��Kj s�/3�*i�����<��y�LBV�~u�=7�D���:�	/�^���0���χx�����3A`Qϼq9���b���yi��5 �7:3%�.a�Ze>�����W/����u�,Y���=}��kj�
n '��Nu��7�Ğ=G�,�b�m�3��Geטs������v�_����X� �Ǌ��C}����-s;2����˕?֜��e]�/L����l�gK4��H�C*R���N��\k삽���#���)��t��[Q��ND	��i��sf9O������*�)��[@�q���y�ȫ��SB�z-ָ��m�����pD�y�^�ge����oТ<ľf� që/L}q&/f|=�5�Ƶ�\��lf@���������"�6����	ե�gE�<N:�p�3<F�C�]�[�*r��ϵo�O��z?X%s�@}vbҮ��ӤB����N���.��Zp��^��g��;;}���w�u=��oMb�>�v�������jT���߄_�{ºq��\��؏����i�։����A�א�ޅMq�&+�w����}��>9sNB������W��9�F��y�B4ފY�����ښ�SrǍ&P�Hs#VH��ԳW_����62�jʀ5���_�?9��H��Í�7&��B�c~g�2��l����
%_N�������l��犬�x�`�Xov�˗0�dV��l����P^���=$n�����Nƞ��I�a��Χ����F]gg>F���WWׁa5�*w�!4=3��:q��=O�e� �_��;)��/|t�{\��E/葎QD٠�c;���|��r������%�@;H%�}i����.�"z��h��yr�I�O�>��94��|�g�h@�d+f��n<�T
͒�he�;��׺��;��Ѻ�N��^���{t��I�Ʉ�hc��:
��h���a�_F�"t��D���ѽ��Ӧ�(��j�oJ��mje�k����܈�D]#gD���v����K��r����m=B���\��b�'9�!�%��Wb��4Ÿ�s|�TԆ7����C2�}�d�6�v���CהY%�0NF���^G��]&�O�LV�'���)��OB��e��`�uq�Z��/*�r�	��#Rʉ�2縠�%¾ʢ�t��G�f L�(���ύܤ7�!�m�?��G�VgI)^8ҁ	VuOZM��K�C9/%���t�C���n�ұ��;`������.W�`�НpI%P��]�"oJ��=�XXy�f��VZ���	=���=�E]I���J����G�C�ǉ����U9��PD<�r	��J-Sg���bHS����M�v�=�M��*h�31��~@��=���[�cҮ�.ͳ���G�|��Pzy�&]�y%����C_�ħ)�d���#p�)���hF��C�/4�u�������W���z��D��W
�gm�mR�-ᗎ�ʆ�`S��\yГ������KMy�DK��R�����zM|˾2�)/�^���@�w�c�;�B���� ]��Ja���uKE�r�s��Y�������=I7������*�*�.E�!}��E'#�y�ޛ�_�W-ۜ�艋.��Jg�%Dh�?�ws2��v��! "n/e#=��_#����ճ�B���)���?��4�l��J���D��Q��p�q$([<ap���Hj�����ݹ-^w%��Ӱ�ZD�+?L��o�������R3�}����$z�g���s]J5T�zp����O0�"���ԕ�u��7�el�d����Bxp��~[��Á�`J���j@�����*�z��C��ې����o�H������v��CP��}�@\����,[nj���� =7?:�}�B���]w�N�\�m� �A^%�-[>�I߱@[���
+�,�,@�����t��%E����V%z��845�nͺ���\_�Խ���<�����VJ<8��y�Z�\��f��,���L��(��h�͟���}a��߷lҞ������'=�I���/�x��vmk���ۏз�uI�W\qdX�O���"��pkU�Ao��5r�r���z����9" ��[�NwÖ��X�Y��,�,pj`�AF��V@��&�,��[��T���{2`a��nˑ�Y1`�p�gze��ꇃ��k���x%�q����>O�|t��s�Pe���(��6�[ M>�'%^�����`WA�;�|��� ��|l<��q�+��H.ų��w�k�Zֿ������������U�I��slj�p���m�?��O��m��/	k��X'?R��	��y��	��a��J�֚ /P�k�����\���@�]H:�fA]�5/�s�f@Tٶ��Qf�#�: PS$���u��dZx�����ڹچ˳d�@ے/	pO�<����n �eF�⴩)l5���a��Z����,)<��nO�s?[�)):��+��h�}Nxz�����D�^O�S��VWT[
��:;>v)�����s�1�|�_�����%�\������u@_eB�%){ĺ���g��W�[���'�E~X �p���\�vv-{�|�`X<��} �X#�[Pvp.	�\�w t��5k��%�����^��Z4�+)�,kÞ�������v4�����Ku�v���"⠜�Ǩ������,�&���^{/=�Ȗ�v�K��L��6<<Sj�	�oJ ��*�s�7n\ڴ�և�� ��������������(�Ύ��9m��&�t�����(χ1幤�S����#A����O���o~ի^uIHs�*��^܂耾 �r�K.�䠈P?4��ψ�`^`�� p�vv����u���'~	��@����rn] ��^ߘ�_c�>��tO�W#0.w#�yV�J�>��/"��c7w����d��p�`4O���E���|O9�� )�]k�>︶nL��:ЙKX��K|����Y���*�W)mt��}��R���/x�0�,���|�sy���sɗ�.��cy�҈�����ܮi�џ�=:������x�?&��^n���y睧���!���X�Z�rw� r��I�D�Ş�,���FPLصt5� ��0�R�<��� t�Õ���"��$�����NC��q:� =+M��e�Ƹe��]�u8�����Ǽr�{~yKn�z�{1�t,�`X;�yx�m���ր�6�slJ�y����Ui�F�9�e${A����>�R�g��<�~���Q��+�d��:麐Q�H�߈#d/�=캮����xX�vj�F�6��ʭ����я~�5���p�?)&���	 �`���{�`�
�N���XfI���2�gb#��,���΋�a��q+��6���s+�E�e��T/��y�ee�v��!y���G��W$ݢ��=�A:�%��Z�1�2+8��def�}���|���oxPh'�<e�: \��˙�2��q���i��Pw+���{p6��L|��?��?���z$�"�
y��>#J}�`�����믿����K��`�C����3��Ud�&P-7'֬��2�by뙃�[�����A��eavn��yBR��f��L`�ځ̖&yJ`Qx�f8xR��uh��!��똅��R��4���h��ܕ��������Y�.�'_./o�+�S��N�=8������]�z8��c����XǴ�AՕ�V�����A�算������,��;���x�y>��uZ`�g��R����K�n�w����.>�e/{�}�+^q�!�үf]�] o�	D�mg�K���rvv���>"ӟG&B���� ׿&��dي�U"�Jn>zȀ�F��] e�;	��ӍYD�5$Y�=(��V��L���u�;r���D������-���a����cb�܊��s��!�����z�'��{\J������
e����/<'��<x�<�F)��f�f/Ei��x��Ο��% ��ӡ�JO�K��2O}�P�2�k��7��氬#Y������[�=�EY����-�f�R�sJ[z�ա@�:����?���w�7�|n��<@���B�����݌=�x\xfa�׮%�KVx�����]˚�W��'�`��^-�`�e����Pj`5�n�SƘ ���v�����@>N�����RDf'˕n�\ϴ{�Ǝ6�_,�1@�<N�X�Z9i=cPr����?�E�#�'��f��d��#�)�7��,PO,`W8c矚��
2|ø�s!�@ꀞ*�� �/��+|(�^��W�:+C�ϓ�~���g^�o�+��8e�m?�#?�g�zֳnn��?_
t@Ot��]Ý���O��kCP�}rD��w�뮻��?S�]�e�:�� �f�g���as�3�EQ������< �v����U}ppv+��2��N	��o-@W=>�ކlQ*���v���#�s����a/~���<X�~E�V�j[�賏Ӳ2;�)+�F��*�+y�]i�>W��5��	����At�z�S��jmd��24�F�c{ ��+�[�k	�в�~���}�}[����:p�,y���
�=�qu����~���Q�}���`�h)�g�kK�w�a�^z�麶4�yf<:9��C���6�5#�����}�Cu�����<�E�CnS�/�+�G0�}O�J>�,�t��5�﨣f1 �jBS�=29[�% v��twd�����9��$�7�?38y�{	�iw˒�(��2�����j໙{~�V����<��Rp����xsm�c�-Ӹ"��P�?�a�7�m�0;�>�;[�>J��
P���UW2]���=ʗӻ�E_�r�0eΖ�k<s>v��Y�0O9!�����B���̿}�k_�������@y|J[{��(��G��[��8�w����	e}���`�t����q�-E��'>��"���A�N�<��%����b�1�k��۪We���..�Ze� j�{^R�2��a����J��yYG��'^����"?k�5��F7˥iB���XS����.������h�O	�Ɣ6VS��w>:�D���ۘi�����dE����b[*�>��~*=��2��=(/��K��k{����=���	����8�/��Nm_O7vJ@�[=,��b��������^�ǟ�{D���#&�E�k�in"�9o�`R:Hg�m�i�B�
 f.̩l�0��������N����'}����Z}���-�r��j_^+�X�-!J�t���[��=e,�#��2���T�� N�%C�]I��֘8h���R�jʬ[�X�9m��.��lG�+��Ł�^����1�wN婒b���Z���L�˘~�C�'�~5@�s��M����.��bv�����}�Qy�w��=�p,;<}�7�
��}�;��=���#b��8��p��2��ܰ�O	7���T�$Y�X晑`nw��4�weATzS��r�utֱ�^v%=��gA5Up�&p�.�m�i-k
aW��-���_�E�z���4�9��=�W����WIx&E0�������5�|���2���`/�s�5�`漥�9�<+Z�;����ea��m��������J�]�f��T�I��	}t@��Z���!��j��<�\Q�u���{E�Cǚ�&�H��� �{B�]w��jD�_t�'~{���۳���WuL�ѡmW>3���h��k�?�Ѓ=���3"��>�4.��*�o��n���) ��/��Ǐ	��9�/?-�� ���R_#�$Կ&��63� ������� �f���wM���
G�׬y՗= -��
�%f�BBi�2�!Д�6�Tcd;i��ꟗ��K	0J� �s;n.`�������k����(��v�R��q	�zB���*_�Ȱ�頞�|��g
�����#<��+��P������9� �y sx�1`>9���� �5�{�J�ȼ��v�@�o�%Ś�x���kVKҌ���¸Q�%��C�<I'���SJ/x`�to|���������8Yn�߱�Їv����u����?4��#& ���]���a>��x�@��]�-ׅ<�l\h��SN9��S~M#�wX@�ξ�R?,�X?5�e�>���d�(Z= }��%ptP�@mZ��M�<k;	 �����V���c�I��<I�#��c��e��� QP �<`N���H��J��ÏE9��ژ#�s�=h���^:��ӹ>��Y̮(��H��l䁗L���qA�P�*;/��2�ϣ���K
����Ӎ2|�J�Qn%��|+�g@�*yhP�KV��pI.�i+�/���W!�M%ޭ)�y�����R����god�WeͶ�mu�0u�T�o+�]C���.�K�����7~2@nݹߣO��f�8���b��K;N�~m>��Cv?��Ö��o��_��sν�j��Ywx�2�h	��(몰����s����O?�ʸ�|Z�o;��_��5G������tz��М���]�҄c;���I���[L|��@��xFZ\�S,tw��h0е�x^s}��M�г s�=������y�$l��܊�t%��u�y�`�i����T��r�[�����s�pЗ��X��г�8��-\���.�4�L��S =�J�WhK\Qm}�d��h������N]�hd�>�aVJr��%[� Aڗ��6��<�z.of���#�ے��J��qFYAaG��6\��0��n��կ~����]|ꩧ�	��#?f�ɮSut`�Y����c���v,�>�� ��^�e����Z��;x���#n����S���7ξ�$n��m�����Aq����?����Ͽ'���Ü�wx�u�)��
C"$J��}�z&W�+3i�^r�s}i�ة�	�kY.Z�=��,�ܖ������Xi?�f���KvA��G���#0��}=�<����M	Z�
$�6�xgX���Q� �;�-���ʀ��ƭD��㶕%�+{�@�Y�[)0ѷ�"���>�����]���1�hs�i��Ӳ֗\�>������x��f �}[-���������Ar԰�#���~B)��^#VH�uPM��?����y�{~!�����_\�_I��MA]}�܈�ze�X]�qR�;����ۥ�*��>����i��'��x���tvɁ�K��������}�s'��_}�'?��w�w�yW���O���Yض.+�~p�������~r0�118q��ǥ%�~j�t��D�� 09>ڰ�2gY �{v˂e*m�p�	���f��O;�Z�gҗ��P��%!_�0�˘�h��dK���7z{j�SJ�>g����,�y����P�"F!�K�֭���o8mJ ���ww	;?�+H�}� M�e�3��D9xz��g�x9�Ԁ���CVܨ��/;+w�O��y ��!���cs��()(� <;���bί���\�ih�ʠmY���w��!�?�7��������K���j�	O�a=?5���aQ?=��	!<蠃o��
r��\�&��]J��h�y(��a�������f���/(�vc����?����?G<���է�r�{��7��+_���M}o|n ���d0�^�.Y^;�p�8��C<΁�'r	�����p��T)x����o@/	��t!� �����1@/��5�s�NN��k�����@� � �Ł�pY ��}YH���ڽ^�򎒲�ߦ�㣬�9:��w�0e`�:r�10t0��� �c� O�K.�R�#@�ś�y|�]�)�ױ�?�>0W���_��ʆ�]��g�Z>�R$?=�5����\_i���3������O�ɯ��u��&'�E\̞��{���O���½~^�N@��,o�����/,й�O��̻!�Q2��Rz'+����c��_��R��/��eA�G��cq����O����7��=4�}t�������?�~ZhO'�K�p	k.�ʁA�.��Z�O�������4��1�*�����[`��ϳ��u���.��L���Ɵ������L-s�tb�[c�Ƣu����d��(�+�W������S�O���pa�=H�]�%��sԿ����1z�b�֯���q�"}�k
E�i���<�����E:SyS��eݢm*�Sb��P��;���;�����9�U�n5�𲢾]3N��g>�����@�?��c����6�������|�=��qY%W�iS ����x�GP�q���
�n�iG_t�E?[�>��p��8�`������Cb}�����-ό�xUo�p���)0���:���Y%�Tn�J�P�y�L�^���J_+Ɯ�ܩ��Tn	lk����Jړ&�r�S���ShWre��=��R{�6�e�e����m�Ƿ��Ã0ƊπOk|_�Y��C@M�mz���yi8Uq�JV^rr�h�F��z �lVZ�5��cޢ��cݗ��gxfj��,W4�6*�C�2K1[Y�aM�y�%:���%�s�4��0�BX*p,,���z�����߼?��o�;�o�w����x��w�w�
���X�~��ݴ�L����
��b��ϖ�������<-P׻[�r����8�|����:�O�	��u�!��%�u	��9�ӟ��!�]v�1������P?5�!N���AЭ�,J����*��Dl�~g��D\d�:��.u�h��:�j�9uׄŢnzYX�,�R�>Q�`�	Ė�Q{>Ex�P�M^/�����h^:�2�rj�~w�­tF������������7 �t��V�+ o��yu�^`�և�e˖�: ��yL�'���ۚS��%ЇǼ�YY ~ �${6�_.ʼ���6�-��k���e��2?��(E�+M�I��f�F�Um��D�z��,�7��u��˩����~I`��Vc;[`Ʀ��O�S�@����:7�y\����5.�e�\���u��)�z�)�����(��#��Ze�����)HN^�;�C�w�9��??�|�J��n =��)��������#@�u�ٜ;6�� ��񿫘��@���E8����� º 8#H.Y(le��#�����v�ee �����l��B++��+}>f�D�R�Z�Z�[�0�w������9�!����X9�j U��y@Y� M��߽-n��wF��7�cS@�v�v�\��Tpek[<VR�J�����g�b�\  �d����R|�k}f�?a�Ǒ���ʅ+U�6�4w�eF�}y��7��Ļ��(>o
p=5,���7��� �O�/|�K�?��_��ٱ��ĺ��#��ذ������n޼yp���]k�j7�5�rn��9��@\�8�i�^�))�K��0�o��bc"L�ã�/�u���i������a���}숟���� � u����������!4q�^�Q�1�" �@�ӿ�Ry"�V����,���$��f�3S,�<`.� h
#�#`���� X2�`������� �Mn��[�NE�����K���p�]�8��'oo��7֢�/C���mrp�~ڗ������ ����.[��1 ���e����8e>�����_�Bz�C��X��q^qe4�g�~ǽ_Z�rYZ�-%P��9hK��s��=�������;餓�U���)4�4��G��Y�^}|~A��)�>��d}�:��\����?���g��n�s�^�98D��r ;/d��V}�+�"@}��|fx'�۰����~� ��~���UA�� O��D? �����YHB$�CLG���p"2&3���Li}�e �	�yp#�Gظ�kNIȌ� zO[R�j WR�Q�����Uh%�7�e���=�7�|�=[�@�����ֶ�p̂-�o����1����rN<�Ň6Ք�V\挍�X����If-�����X�s�Zળ,�b��xlՀ6ϗ? ޮ��z�ҨK�d�����E;�r�<��~�9�y�5S�AX�]}��'��"��U��3C��'pr���fY���+��[�����ϑ����ޅ7R�-�����+�ᨣ�Z��}�,wxF��&|���^����b��@m��_���Ź�?zvmscXwK�4�惋^Ĕ����C��� hP�;�<hU�
�,�k���O�`S�;��0�	�����sYn�@�d!C�l��@ h�-Qo��Łĭ�)�u��d�y\k¾���+�3���5>�V����c����q�g��iT�����1p+0dUF��X�v�C;����xQwm�x�Ҙ�<�}Y9�{W���ݷx!�`�palJ~���\��t9����1v�9��L�8�h1�7�����mV��o��o]�����jE�`�%�{s�|:����"�+Bޟ��p�@S ��
x�ռ����l+��W)H:���Q�ћ����E��z;V��G�:���0��Q��^§hǾ���P���ȏ��_���}����Dd��.1�:�'1 �p�8X��X����j��;����e���;R�Y�w��}���K�RS����@��J���1�̖�w0p�fL!�g9]V0�%e��)O��s~/�FǬL�0���O	���,d�,��{�%˟�q))�5��U?�Qx�{9�-�96�(��9f�;�;��g*)�S�i4=>a����ۿ�T��d��ul����b��������c�,r�������2��)y,ݲ�P�(va
�/���[�����&J#eCGĪmі���cз�/��fzl?�#.�?�#�ȿ��+#�� �&LDĢ���Jw�Ӕ�rh��#�vP��DD��!`�PwP*���e������3^SpJ��ў)��F�ʘ�7��y~�}��=�.>��>����Ӗ��rZ
�{}J��lg�2n�D��]0�Gﾭ�VƘ���d|K��y�P ������xy�3��Q�?��V�+I�]U�H��<�4���)��y�>n�6Mᙩi/��w�_��_��8���׼�5ö� �M{u�?��7�r�+�}'��?x���_ҥ)��#�n�D7����9���c��Bgɖ��z�)yܪ& W��WweA��o����H}e�zX��E[����Ҫ�n� zD-��G�GO���?����\����N`��&��S��K���]իAպ��?j+�4%@]nwyy�S��na�30S e��EZ1$VL��s�߲���8D�
���|N��8yy^��%W��:Kml�O��x�oM��瞦�"m)!��N}�`���y��JJ�C	�J�B1s�uV�����@�̕����l�U�Ѣ��_	�[y���<��Z�N��9�V�+"�K��q������g/,�{GN�-^�k ��7q�K�Ȫ?�~�e���2���)�\4��7Y��2 �lk��<��r�Y�o��5��*'h�O|ߧ�c���cݦ8,��p��|t��$��hV�E�\{�7k�h�Lк�N�;[۴��:�OZ��&X���Zc!"Գ��*L� ��IRSZ�Rf�\v˲k�/1�[�<�����^�3V�[�(���[��<��+%�[��z���k�c�  +ї6d���O�R;J}o	��<1w����N���\oN�<��E������,+JG[��<�<W~_�GF�,!��IV���~Nu{<������^����+|V:�]�Q�].x�S |Jڪ�>g�}f�����������&h�]!�_w�,��}�2�$˹��i#:>��CC�a�7�����us���q����hx�Fc�zG�3�%{�9�FmU���^Q\,�������O�[e�����>��Ce���@�����4#Fr�<]&�[�.�q�@P}��]�M�j��!�ֆ���w�m9����%�/j�gY��nӬ��c`�h�j �`��<�$�)�<u��13�gI�X�-���E"{2��r�g�~�ʝ�R���ꞇ����D�#�k�iV�A����P���Cq�?u�w@~�K�{V��V hwē��+�s��o��)�*NU���ǹ�ǆ��Mۿ$�9{]�S���KSX��܈To�-)
p Wu�|���nv%� 1�X� 9�u\�-�!���ϖsv|�)�����7��M�,s~��PJ���:!���
��{Y �����	�	j�ȮI�m�q��]�	LP�C���z\`?��ښ���ܳm
��6E!��=2LT�(iK���I(�zyl�?�V�L�.�s;�E��c^� ��v��5zy=r�=[lS�pE
P/����9�(S�����R �ܕ({��ԼN��t�[	���%��>:��9��~��J�pK@���<����h����
�%����$����롇���&� ���G��%��v6D�G����[�j�`���1�����P��v�C����y� �_��!��?���ǚ��b��(T/�k8L gC����>�P���71�'pD�e`׀��r��EB��%�k�n��!:RGN}-j�O-�yVZƼ��bK��h�l��,�E�.�s�����c���Z��w��f�~C�m)����դc�,��N��@M^,a裏u%���E�EjB�<�;u�P�<��-�p�Opi�n���k�`���[ʥrZ�5�˿��S�Z:�<K�K��|�����,���)y�o��9��M�ͷ�q�pB< �,�LSs=c?��Q0fQ,�n�GwE�[6�/�Z3@����ݧŚ�kC�9��&D�DT��yI#bo^I���L&(��sH�@ 
�:{U�ڧ���V��~C)!�N3,�wy��2��t(Ok´�4��u��"�P�n�d�����E�˳}2LVlK�(	��f+���:�|�[�&����.�,��Y�<m�B����<�o���On�����=M���'���Ry@��{�F_��t9?k����)��2��Z�5=�a ���&o��l�ϮD�m%�����y;\�*����4�-�/��� �,�y�{ſr�W�^���2]V��WV;G��m�|�ͭ�U Ut�,wNv�"w�:u�/�N�G��>�߰���H�+���>�5 }�Y�qp�Q���� ?#@mP�W��Y�@[A]p��
�� '*�	z'*�A`W}bjB�в�=(��}	��B��E;^	ȵ����VY��5��ʷ�ϳ��"`�mB�|�����?w��Z�P	�ǀ4ϛ��kK	4k�����oM���0^��+��WZ���US⼽Y�r�-�́��Z�xu��<�������\f��?���Z�-���/�������8"|�3����_����ďʧ���V�s��܂ƻd8��{K��7�:M�x���w%@W�^
h��P(�t�+{�ךX����
��yA�CKu�m�������+4=X`�r�L�=g�~W:w��^�c]��b�h��
�л�]�x���ɠ�¾$즎U>+)kj��t���V���f�ڢ����f_,ǖ���5���^kSv-{[\9�"��,����~���Þέ���d��7x�F'o��k�_Y��훗�K��r�y��xg�1j�����3%��[�)���qroT�]zlY[��kK�{��U8%��Yy��f��hI�K~sM*İW�u^�gJt s���π�����Hs{�����)qjߪzs���ʯ�1re�/2g{ﶢS	�=���D���j0g���g(k�9k�j��$`Nm�L�&Q�C�����=ʂ��fQ�}� �2�V;���T �v[W�<��[��RC�� �5�c@�Ҿ��[�ާR�����%%e�~�b\�
��7m��|���)t�f�eOy��վ�%��xC�ʚ����y`��Fi�1pE� ��~��Kq��k^��������^��e�)��O�_��S�d��C������1���uv@/Y�� w��N#���+�+WE��#+���z�Bv�o��=9���R BXJD�K��ޔ�D�!�
ր����ia.iN��Y/g<��0�hM�c�p�Ha���hKڌ�Am`9�$\h?m�ּ[u��� _�
�=�BׅN)4�	�b�l��g:�4��eA��y�ga얏>��Wh[��B��]�]��2{9������E�;h������Zn���OC_��t�4s�S�l�O�V�<?��K"}��[y�t����K��Ng>g�ww-�:O���ׇ��#���%cj*�;_����t~���Y�O�U��-�U�Kq#�p*���$�	��1�e�d��1���%�����f�g(Np_�W} gܰ��?��vЁ�U�喖Lm=_U@���6_z��:V��� � �V�y�U-�fK����gۀ���z�ݹk���`|?�V�x1���#��c��1|\��b,�+BJG;j �ӻ��������Z�砕�u�|,K Qj[K��S�R�����s�B%���Вr���	��Di� E9(�U�s�Sf��ȣ��h�:Q�K��;@E�g���]Z�%?����<�}��|��ON��S�>ӿ���/�c�u����e�C�������{\�5X����4�v4߫^k���+�J�-��J���	�G���ٞ�����0?v�	�D�୔/W�?��O<;�� u��4u����ߢS�~����X�X�hK^��G:Y�h�D=�ݎ^���Z�˝㑲X-&����5�-iٹ.Բ�dlb�Yɫ�=��?o�b�q�:Je,Zo�n}P<�gc�Q�]5>hY�*�T/�?j��B�t�΀�i �d��f �N9]��rsһ��-Y��)c��}g���4c���ַ?G���u�A��yt���� ����ɛ2wZ�?���g��c�m�琽�y�Tt��R�=�ڍ$y��|Y���xP��Y>�Xc��Na����]�	�V���E����oW����SN9�)�o�Y5@��{��/�Ⳣs�Š�JD9`����`mu�I�>C�E�����F����vKdߠG�8��4pz��,u��ԥr9��:�d�ү�H��Ć!kJY��"�,�ߒ�H9c�[�ݖ��@k�j��+J& �e^�@���oXuz����@=el Ú ���:��<�>_K`��A�{ݴ�AZQ�
�s��#]�����YV���q�&(q@��-��f^e6��V��]<�<�ϒ��nmc��. �OXX�zǻ:�}y���5 ^�����^`\�*/<+0�߮%���/���N������j?��n8?�~�/�\���n�S�s� @q��bip���
�`8�Sm c��aPT�oq��u���3�F����B���Ba*}r��2I�]�py�g�_��oy��wW jBi�ǡD��+B�_����>�Ԓ�#r[��@_����n��h3�rYp�~ y�לoBYB�w��6��d��|D�����r�,){Y�3�~mq�*�D^�&��-v��	�{o�3��dC���W
��%�#��6��/wI{^=Gy,�wV"�K�˹��*WrZ�d��R�҅^8 �{H���At�늗Z��7���7����N<�p� c�~���@���h��e��g>�-*�s�U�8<�����A�} >��B|��%�|�Ji��� s���-���C��9��8cT��ط��9���TƘU�Z��*�4L�)Z��V]k�<X����Jy����y�Ef�vp��-�`
]� ko�t\����'���%>��^(���J
X�N�� IIiuo��Xb�2������n_��u��r���s|W�k���)O��nɊ�+cʂ����Ɔ�G��}��gIǊ+@N���{���Q�������q���r�z����!j���%a�uG<�R�{K�}���Ͽ��S�<_5@�mgEg�m1ؒV���i�JҖ�Aw���V��";Z��� �i]�7����L�ʺ馛�#dO<�ā��Px�,���U�YHf��zN}����8���<}n���e^����[J�B$�T��VwK�Ҏ)�5�,Y�c<��[`��/	���3�ػ@�t�Bw�`�W�he�/yC�[J	^���1�v�x�-h�s��[�%��5�3/�y���Wd_k��y��ܞl�g%!G.S����ͻ�.�䒥��;o��++h������r��1��,q<�S��Bg.�]�@a��(����͑���Ix��g�}Y�߽�Tʻ*�.������� �!��.��]�-�����i�6hp4�y�[�&�4�%d9�0��]C�N��oZ���k��-?p:}E�-u�y�e�� ��p��l	�Yn�oՁ�íQO��Sy��%��^��2�	0�E<���ď��nOW9�k���W��e_wP/�=ּʖ���yk�\i�y� ��̳�����2 �<\��/��6�N����`����N�#�튝�S�Z���˺�Xdy���i��3r\�4D���9]|��'��CWw���=��ޅn��>�������c�}�	'��駟~}�oYY�ת z����>!4�}�9������X�".�0�bJ���E�5A�~�0P���Hwi`~�=G�
�uL�O?�Nm�Y�
�v�5: xX6.��)	����s����4�[�uD.� ���?&�J>S���M]i�}oY"*���m��%��p� �qiYN>fl�hI�-�k�̣�m�m�񋏥���CC��~�7}�%�p�,pZ��9� oP������E����y�Jm/���<,��X���y$��ے�8˄�����iLDk����X�d����B�f��B'��
����X���:7�]w���4�P(o=묳��\�f�U� ��������S��5�ݬ`g6N��m��J@�	dI+8��F���+���IAX3Y�׍m*C��i_�4����o`B�3�[ɅY	x��҄i���`�Ƭ%p3h�ʫ=D]gZx[��ҳ1Ń��J��7��,�}
��[�[ed>���qo�7o�+r�&��ۓ-^=�o����(Q�&h]�e����ǜ:)En�g�����e<M_�k<�@���-Y�y���\RP��c�Z㐟��%���w�r�?�Y���%ùw�]�X�l�f9K�*�gX�O �Gc[l7�\�Oygx�@̓k����-�9�䓿�miGq�w�t]bG���m����Qް/+�5�kԧ��2(:@ W�:����v��2b�ɭN~�+k]�Ş�������>p�/)����`r&&li��YQ�1 ]�`�cBgkA���Sw�l9�,�����������$��,�,�3p2'K�=����^�r�J��y<](����v�����7�E\�j�WI�#	��=�^��c�߱�s;�z�J���,�)�5/���,x�&��U�[�^��΋_�򗗮�⊥pg/�y���7:ח��ݕ+��+L߳�$�?�q[�ȗ" ���x�L �M諲%m
�V���<):r ��p�4������|J��5t� ��r���{\�u�'Z�ρ���5{��r�����+���b���0Ҕ �R�kB�'��l�L��j)iS�q�8f=B5���������I����+%���ގ,xk�5[ S���g���-s��\9ʀC����Ͼ��p>s���VR.Z�*)
c`��1�G1`)�Doo�N�|o9G�:��[Ͻ��~+��L7���3���j��<�\����%Y+��KW0�vq:�˘��)z�.�\V8r��36.G�����!��2��ç�z�g�y����j�]1�Ǻ�~?��?��`��D@@�-k��0��%�x[�U�E�s�����)��� �%B屆�|~�mz&�@߉-ЉFrq����V:���}'`�bY�}~֢c���^��ہdQ%���Tގ�Ю�_���Ku@�ɨ^o[V�����V���oc^ o;����d�Rk�~'ԕ�\J}V�<]	hl�vS���!/���!�M@�o�E!a����6B��io9`  E@���K��y>yZ��c��Ծ��5R����5�a�/�(,5�4O�d|�Xhl�\���������?��E4�d�b�82��S�R��G�Ҡw�z}�����ۣ�K��/�@{�g�qC�ݵ�H+���k������=��̓7U[�uvLapͮ�`Lh�G9ꕫT�G��T9"���~p�%/��9�z��p��O �:T���3j��}�bH��<��)��E�(��X� 2�)�-�~K ��众���(����vd���C�[W<�4 ?��+��F���������Σ�b��-�î��w���@;h���`J���_��W�"��g����BV�E�E��<�'�^}V��"�u�g��k�=^^;����q�/�%o�sW��5��G�;�?����w�����wŀ�݃0F�w��5��e�ic�p{��'�P��ݱŁ�&��#*� H��g1�(�\�0��gٶ��j��mG�Gۥ�1m|�DJiq��)Dϒ�7&Hr���+��
@�'.h[�֘���%k��4+�_+������]��7�S.^B�O�����4v0�`�<
�c�;�Om�j̩1�4��y�<Q;�eҎ�&��o+z���WK�����+��Б�X� :���܌#zwy<�C�r���/Om��o��k�������|ғ�t铟��[�bl)sŀ�^���b���k�4���fF[�:ry`7.pY�X�D����sx,\��v<�Ŏ[_y�t�	��rË��l�,��?k��ZD�=9��75]�����Z���t��p��y�?e�(6�4.��Ѫ�2t����&��_���зdٖ���)�JP(�}}4�[� � �����/Z�<|�|Z��ۼ2���3���7xT���:�eW<�쾞β��{��L�"�}!�o�X�����K��নce�;�<�+�[n�e�����E,�;W;k����Ofڬ�:���S�,�=l\�c;��)7��(��_ʀ��ٷ�p0�@_ֹ�_�z���誫�Z
��/X��s����>Luӭ�[�r��c� �2�ϲ�ڱ����� 5�<[�-���[�J�t"�P��J��n��1�%k��.��|��v��.v����G�.�e�1t��t^�:}\�:�CXh�N_��$��u��M��yI�59��������|��R�Ҝ���,uor�4G��*{�<*��<7}��7���|@�j\���x%�;��Gek���R� �Y�zn�߿`��Z�x�z�����"ק�\�[1��������d枧!0�eb,k�Ғ����(Iy�S֟�i'�n4��I��s�;m=�6.�:V9�AA�
W��,�*J��RĦ�
Ե���9#����R �C,�*Y�.��,��ƀх^I�b���^;����������onM�f��������9����R�1�'���K}q;�uM� l�� �wܴ
�#��]6��K?���9+�A�O���T��qw�vL���_R��Ƚy�\�����ۼ�C;�E��)�c�~���2�ߖ�4�C^��\��i�D7G��G��=��τ������)t�^iV�A����CHa	<K�Um����4g�'�6�ղ�VJh�'W�bE8�ōv�����������	F�4H��U�< z�� �� <���uA7�h�aS+����3��&���1���5::?�T.��@�,!��y���-Z��E_R� >/�F=���mi�8����2��4��� ��#�+G��w�s���eBI x^�1�j͹�����_��<��G�{M���(��bVhy6e��h2U���إl��8]آ؜?r����������-ah]^ӿ����	 �),�m�m�Y��]����/�ҡA��T9w�/��kQL"��rw�_�����^�jL�KF�-���=��2r�#8�Y� �~�#�㉄�&8	
���^g���ۅ��g��k ¤Zm�_tl��s �3Bz�b���-#FS��|W�|��]��;߳`ʊ���92�v�{�J�\�W.UFM�f�/�1U0������%�����G�4i}���P�A!A��������*-7g��|Ք��|�<3�:����f�9PS���Z�a|�	�˛�y��P��b��6�l��­��0��2��?����ZkzT�j�dE���#&��x�����3t��G��@�9�ǃ -��InA�J.Zgښ �	�D�	X�ĺ&�,h�&��k\��g��+J�,n1>k�~��,s) ��.��^���9��P9$��?`���m.�ZJ+��c�}\��S�����\��.�ƀb*�8��@������+Rc \�T�'[V}���-�l���VR(\(�k
}}̦(�5�˜un�\J-t��}�[,X�/�뢡�Y|��-�c�~�������K1,�?5ު�e�st�U_/�,+_%���ֆ�1YTy�)WH�h&�c�!_`,@�����(Yʕ�3��}����B�~��N��x�)\��\m���Ѓ8{p���M"�oe���9�kѸ��2�˝"d�i˼i�؞�mkX��.�l-��
��=����r5q�W�Z�"�����~C4<W*���.���M�yi�¡$��5�,+ �قzᔹ��^����C�"�R�Zu��u�Y�{����b�)�>h��������dEv�w;�Ձ�����T O��g_6�c�<����?����Ted�:Z�k�c�Gi�:{ѹ�oi���h�%��"n���R���ݭ����+��wM��`�Й��rSr9�o���E�����E��ړ�v����Le�xٶ�z�
�9]����1���C;<RT���7љ�9���z�6nQ��=Z��(��r���P�.�j�^@�E�ve+De�ܚ.\K�\�ׁ�-�x��XV�����	�[��~
`de���F�o�@{$����
c�;-�a�^wg�v������� �-��XK[r����7����y��g�C~�}������-�x�y��0�|�1���o|�KW_}���~j�Y|�-�|1�������e�t��V�*�����m�&XK�k��g]s��-�$Z+`���@l	�9��(�]J�������@r��4�S��:1��8C^�a�KA�馛Ea �=�\:���-p*#b*0mo^Gx�@��)[�S���%�t\�[�skI�J}r![��ls(����AN��f{�wс!!sJ >��n��Y�)_�c�a�_�s�7+���W�y,�fpΊL�J���S�����ћ-O>�2���~K��/�m�9���>o�{�m�zN�"@��%��W�ڮX�+3�7�����5�x���KP�@��4�,�j��|2טA��W��t A:zF$<���u?���@Z�.�:AX�*��18�� ;)	r�k-_�z�i�q��=G�]����6ج�x1N%�ɚ}Mp����u>jYE���z�%�(	j�pM!��Y�i���U�1K��pP �@ҳl�K ����=X���ְ����k}��	��▬ٱ�%W|	�j�R4�{��K�7�"[h�<�<<�:k|��)`^���&y|��uf@#�_�_�Tr8N2�!,�����C>^�n_�]q��}��mۊ =&�n�/} ��`��}��hѼ�j�{��a�E��Ҥ,����-����EE�q�:1�M������G���D�è�}e}^��mmR�f��9���Y��ۯe�m�o�ƻXS������OY�OU�<�#�o�?�~x�J�IZ州g�� �`��@��=�[�Kї8�b�VC�ρ�0�m%`�����g�f�;�W�[cRz^�Gh��#/sy&ތ8E!���N���m��sy���� ��b���X#_W'�-2&cyV�"��Ƽgs�A�d��^��C�������1p�VQMmiմ��Kn}��-�Z��_��D�عO׻��}�v=G���Hx����`��)�Zf�Gɳ /�p��?k�R�cMy��P�����34��20���D���ϵ��-d�'+.<}|jnx�]�ǅ�怛�M�&�K} ���3.�9]�нݴ�]�S�P+��x��^o�OZu��ގ�/��X����V;V�yIq�<�"i
���N~mX�j�٢�[����k}�`v�?�ϒ��o��] �����ڕ[��Յ��W��/ ��]���lY�L"�]߹��-k�:6��n |��e����e/���i�}_O�Y����<m�W`��v�]Z"q^rk���8��Ƶ2�SI!qe$ӯ�K�[)*>+Ⱦ-�w��N��rw��4ǽ=�/�o*�RʁF�~���c5xsJ�]J�o��ZY���.dZ��l�+<U2:C��}�;�kE�@<���A�]64ךK�@8\�D���8
�쫽�[�S��9_��n1�w!���*G ��(9���z�A3JC�?������E/R���!����L.x�W��W����OM�B��X��5`l	BW�Z3�;�Uѕ��� tk9g��!+lz�k��q�~����������'.ė��/�����U)����+$+�*C�O�w����+�9`頙�>��wVB|>L��<N�1Ő�]++ϧ��V�c
��eO��ӽ��#c�[����~���s?�<�5���u��/�h	��|E����t/���i�4\	��nQ+H뷱1���J�;[A�W��X��������7qً{��c흠"y$	��Q�rǫ�汎Կ��+��z�˸�+���6�l)������2[s����Ҝ�v�X��J��*ଐ��5���V�ea^Z�@:�����߽M���c�#�� �D�V���h)���F�i�+;y\J��
������>F%���Z[ƪ���H�خM!7et��� �]Ǆ�<TX��<e�״LH,�����:(F��ڰd�kۛ Y���G8`i�^��6o�<���z���r��:Y�@�,�[�h%4�Y-�V[�tj��As�0�,�� ���<���α|%���RT�r�`����ց����-\-'��kW���aT~���>`�z�~���� e ��k�m�<���06�S��s7[�% �-ϵ��J��J�ҏ]v	~�3d�Jqn���f�W�Q��E@_�+���^mg�:�}�*���@XB���\�"7��k�j4��6�8^m�o\�t�G��,y�N��w��;Z�ɂ��~[>��� ��ܾ��,Y�XM%Y����������?��tdT2�dݭb}.��]9���v-i�h����xښr��E�9%_M9+�-)w%9c���J��� �����{��]�S^��ňLJ��9E��bdn����^q����<�TB�:�H:�҈`�Uͽ��ڠ�X�'ֻ�<�£t�u�ʔG@��Q�*C4���M�Dj��ǉ�	Y�j���S{X��`����5^���Q�\�S,z�1&�k�c���Kt��`=�%o�nբd:��<��.wh�L�._}g)�8�]w� Ӹ�� {����t��)�[M��-p�ӫ<��m� �[�W��N�E�u3�5�.(����!�m���BQx�).�:ફ��>��1yv�t�_��븫 ךH74e,�O�E-WY��b� '�Uٲ�9�N�C68jV
��&��1ٔFt�Ҡ��Ƽ��~v����ڤ�Y��\�E�Eˡ����W~�j���Zᬭ�:��pdLIp�������-�I ��bu���fF�j/�J�^�p�?��#[��+�N�E�1���_�XT���Zk���2�f15Exle�g�Jr��X�@�蹜Z���2A&(X{�X�n�^+r�l
Fڄ֝��Q� ����7����k*�z�dq!���8�^U@L���t��ṑΣ�]��7.��U.K=�@���	���@(M�E�k̲\�ؗ��c@;�a�dkD����Z�])�yl\Ij�#+�*��@%�V��/��-{w�CK��])c`���7
 �4Й�����r^i(7��+'S�)+�%E]�����������E�ϔ>��]�]��}<=t�cָ�XM&N�0��y��W�}���y�`�W�a�3hX�~OpK��@h�&��U���5��[�/��U	>1�����e�+nx��e��� Ľ��%��]��h���u��Ԅ�n�c�<�ҲJ�[��1P-	^�)�	�V��/����׼+%�Z$\/�-k���u����g�:�g)n��#�sf�S��S��բq��{i|�3��)L��2�c�V�ܶ�A��/�Ϳ�}�b�W��a�ﻭ������@�=�c�(	��՗�p��b���� �vd�)��jVSm)=�5:.r���ܦY�kN�S$</=S>N��w	'�C��"ޥ0	/�W=Z_�\y΢��l�jK�;[(%������h�ǳ�'5@F����mq ��d�a͔vm����3�)�(L�|_��9֬QWh�J1��I�*�H(s�����P^=��:y���>��r^���A���q�),y޷����7���cj�D����R�ϠG���w/'ӝ�e@w:���BP��%���˖�=�=d����A�O<�lb!%ي =��N�Y�ٸSy=�0�*S�IHk?��ٴ�\ .�!�(�mnX�<�`��M�t�^�	�O9唥��*0��.H�)��e{>��
Z���_�Ok`2u�](��͂����(M����1����o+cK� ��x�@]ef0�鳲_����|�������M�u�/�W��e�M����n=�����~3�skq=7|����cV���<u3���6O�m�v^��@P�Xs��Ю�ص9���~��Z�Rg߯���W��e}zr�M��nr����_��A}%�}��^r)�����󔲲%�>��J`[k��L^�-�\���N�. P5v���+���;��c��8[���������xh��}�#���%:d��	W�JuB�������pk|J�QH���e�TS���?�9mI�Ֆ(w̅?E~�hel
Yxh>�t�>F� Y珶�ڟ�8�Ε�'0W:����w6B�	����;�})
����U��	[ܲ����LX���40oy+IO[jVu	h[�e7ei�a����ց"�Y�E��6E���G����Q�9����d�]��1�ߢ���Ƶ�̫�,S�b&���E!��-����V��f@�5Х�5����jѵ�^�TOJ�WW�ó>����B_�n�M���Y�1�s�Kp�) �'��N	8jr��*��uY*������".s��+�MV��5��������}ݒW:�����+��ҁ4��������><s��ޮ�Z��Y�.�kֳ�`�Un�}cc��y��i��))��%�W{�'=�s��y�h�=v��wL����v~,2��;��;w����g�x�wi����)�6��7?��u���i�=�y^�R>��e� �A=ϋZًȶ���jX��n��K9��ɧ��fE�>����3�|�l :�YS�u�����Vp�˂�d�֖,w������b��=���e��xE٫�iߏ�u"����,@�fĴ����ZG���R�
���,�~ktp�G�$��U�g���J���������6J ���r�z/�J�$M�S��	�л�a���6LM3f���T�<�J��%���4oUFV<�<v-�՞��mc<���9���*w�>_)�?�8�BIPM�Wh5��)u��4n��M#��ZV�c��\���z����Hi?ІS�4�����{�|��P�&�RW]�9�Ɵ�,����<5E��	�+=oyZ;�Y�ǽ����Ԣ��JZ>+=��E ���\�s��N��g���G����9�un@@y�����)�!�S�+��K�<~�ϰ��m:O^�s���v�$^�V�"2���ʫ��YV��z<dߣ1/V��l�|{=_1�G�Wm�%������b�)e��d�i�Ip���N��ow���/P��2��V��]�*O���Yx�2�wmy��΁6�/�����%��k���%�/Y�c�� ��}m��G��P�-�*���r���}��kcQ����"��X��3`^�%z��gQoH	�Kc���Y�%�=���w�r�9��V�r�E�˞�e��Xg%�T��S�-�|J�W3��5d�c!����"�Hs�&Q�.԰LJ�\�c�[��(�|�zrk��m��!� c��1Y\��*Cnz�1�� Z��O�(�KZE��/�]���v=�M��}��?���ȳ������cc@>ʤ.o��<�[� >~k�#�Y����N=JC�~g���>��j?;G��V�����j�D��,3��e��g��>��x��1�������y�gw���<�<�;����2[�Zg��}��xp�k}���`Z���x�斏}	d�,r��6d�j��"�>���B�FȮq��^"6o;�U�Y�1y��ж5i?+:����VD�RO�1��)u�4cuK���T`+`N�.���ґ��q��	N�']�����ٓN:i�����# K�Sm���B(����mwz�Ɨ�zw��ߩ�I�&��7V1yݒw .�G���k�-d>���@�{ޅ�@�$������v7�"s �V[]�b�|����Ǿ�F�@�h�Znxh��5S�<�+ �vgŖ��9��Y*���1%�5_�o-�l�����"��'b�����7R+_M`� �y����ׂ�Ѷ5.r�s���lYjꀆ��~C`�i.s=W^��-��ӳ�o�y xy�F�����1� �2�[	��	x�|�� PH��@�����q�Ο��Y��8U7J}�`3bo��*������*��yY|xbHW��ܭ<��>�b5��o^����|
���/�M�}��e7+�-�Re��ީύ�lmg�h
�����<c
�?�R�zL�U����؍��ޕ�i5,t.�S�O��ث���	�@�A��m+���U.�9���>@]@/략sߋ�e����U�@Bn�;�c8:V���G�*�
LM���[z�x\��0�^��$x}�E}j�� 
���X����F@ �� -�J�[����K_;�sZ������<!�OV��?˖|�T��bM	(Yǀh)O��.�t�]^W��~eŭe��Z
�T�NM7���>5�FN�"@!. ��;�A8���b�y˛w0[��WJc��I�P��׌%��CB]{�e�˲��]�����XY�����2�P�B�g*K��`9���KG���{��}��wP$�
UF��E������U�z�o-��J�[�|�up�ҧ���Q�&�� ��L��+����.��� �ln����o9�@ <�Pxp"z۽g����B��������]eR���7�,_�2<����>�>�(��H{��!m*���z�\�+�- E��6P~�e�Z��卹�瑡�rV��)�b�$�v�׊ }������wB�f�j��V�����]�-��u@j2�<w==�v6�!׼,~���RX[W>���#[��y��m���Tږ����T�vn��P�	�8���y��$n��R&��Zw����^muݿ+��Ѯ�7�5�W����G�����eV��r^����K����ZSTKcL�&q�3�K��JE���%Z����e:���S繧>�e�SX���J]:AqE? g5�qm0����&+��^m%�M��`'
Z�0pX	V�~��nw�+/௲�ҧ<Y��ׁ4�ϭ�1:����1h��ϱ�Pl(�]�����am�Z�����+
@W�<ӻ~��Е���l�.��}�(%pr�g�r jѿ5�)��|�w@@}���jk����16� �@��+�'��)|�V3��t,w�7��A�BP��L����y�7�� M�)D޴�&��]�����)m�i���ܯ+�&���~���ﲸem�%PPp=��F>�������A?�[�-�^�Ρ4�z��)ty��~��$��R^4��Iv�*_VJ}q0'�_���]�^V8sk��g.s�Q&��:`s�.k��f��q"�)������.��5�Z��-�<>�|^�zYa�	."kV����R�m_M�X��픧��t�A�zL�!(�5L,��$q,M0_��Ҏ�y%e-��2Ч�!��%7�TaĤgTguK�+:�;�� 4nM��	�����h���D��Q~���6��7��Lx��8N���Gф�B�����0&�K.ٱq�Lo|N>,l��--�R}�Mt��X��  �R����x�X�pe�sT���ڭ2�	9��|F�(�)u9�e���\�{��8�ŉg�-�a\Xe��7c�V��y,+l>�N+��[��q���"�ۚ��:hiQ�r;J��n�R�k��#4�L5���%�ZF�X[f��.�����ј����z7�μ�l*ݶg���Q�;x��D�+hNV:�"�R���Z
 n�|R��ԋux�tҜ.|9���`��z�:p�%߲�ւ�%D;#��Ty\�u��f�2ns�A�� v��:tc|p�g���r�'��:xpJ�g`B��}謨��߳��qǽ��nO�Z�tg��D���YVvL�&<s9�� ��Mi�+���R��f����G���a���^��@ M�8W�i��ii�Q�j�Q�XV����x`.uY�l��)tJ+`�hXΐwP��i��2�'8-o����FU�^�W��Z�3V�����t���@ ����"�/:�7�:"���ٗPܪf,�둇��pq�:
E~��T�ϣxEk�#=ed�&���Q���;[�J�YΗ��~�P=�ŷ��M�Ϋ�c^ �Q��Q�vK^zUS>Zq�C�^�"X���}(ٽ1	]m�Hgz��S W9%���%l�V'�Mi��.@���������%�e�K��t9��e�q�K�v��~��|��@=��d)N��Z	�0�w��=̗�D�	�vc�cqa���c�+�[���}��Zw �4t����ɿM�oVr�|����,@���Omߔt�ގ��K�\Κ��
ee^t�D�x�@�EW��\�ɨ�����nE��Y�]7�p��h���z]�DXͶ�G��'���'w�:HMmCK��	Ą��0s��W?�_@AG��Y�H�q��L�;�өX���7�-w��IQ���QG���9,M���61�E�.c`����&_�;x��3 k��_�&>�1QZ��U�@���u���(�+ �X��ǚ �~ڡ��<v�� �Ƶ5M�J�l�����e���q�M�z�?�P�bq�n%�ɖ�@�Y4����=k�:pKJ J�2]f���;�5�bL�*��C:���"@����~����T�;�vT�EK�k���c�n��z���.�e����\ (���:M}�Rȩ�X��Ǟw�(P�o�p�,��jך�@��eD;8>gZf���K�O{����wr����������]���]�n�#�}=ܟ����v����-��N(4%Bɚ�ˀ9�����4�Y�2�����6�\�i��>VF	tK�Y}+�3�F�mY�e����d\����']�=�OI��Ӭ����f�!K����̱	�Q	�>KH�t�Ve�q���W����`�q�� ������&[��:<�Z��[�Dmq���E1)���y�ﭠLwS:��� :�.�Ņ�w? �ח��i[�2�p���v,v@�]��V/�����9&�Ck͵�F��D��?���r0W:�#}~��V�T@G���L��W*���u���<�Z붬��g����y���mŀ��7&�h��q��XY�,���>oǶU��Hh�p���J�U��2��^�Zk���y�#p+�-g��������?߷��/��|Z�(�,s�D��x��z�<*�hx��-�����9�c)(z��������w���R�E���$���e��sԺ��s� �t�0����߲"}��\hA�3y[|�x�/��S��g[����<��)�c����[)��,�\�����_��+����������Z�3S<u��ZW�.�_1���tO��tꕄy�f����,�z �h �鳬N�dq
�8 ąR�E����N?ԙ�g��$0$��#^�����rа�y= d��3�}��~�2VzE���O�� �G���ʡ-%P�)X��O�Χ�v>�G�~�k)r���l�7ӓ��%����|�бܗ��ٚnv������ےB|���V���;�3[��1>֦�O�����@��e��n�+)�<1>��5���9��
���;{�^����K�?����W��������y�]�S��/�V[׶�� �ڣ3��@��]+]��xJ�W�f0T6�t��Xsƍ��^ƶ�onw�)Qi�'���z�WN�s�%��e�R�U˘sG�Ja�3���뇭sv�~�BN�S~h�.� T��κ>�����`�A.�C�I����Wh@��ݿ�� ��>�J��oOw/7{D2��ܑ�-��,@o�7䛷]��׀��d�o�h:����=�5���7+٪/�Q��|���M���ǃ�m-ŭӶ�ݬ[���`�{B(>���ű�V���Ys��� CvaJpc����������d��4��U"5�L@��UY�D���]��w�������}m��D˫L)DM�Qߵ��JގR�[}ʴS�v���g)�0���]m#h��߱���蜯`�E���"�"[�ce �%@�k�q<�Vד� ݗ�jKm>n���o��Ό��;�g��ǧVϼVn�_v�{=k)K��:I�xȣ����-�)��#�6��p��cg	>�B��#��%�YKU��sj=�#�KB��]��?�ќ�N$�\�E,{�N9_�+��裏^���������h��䅇�� �J̪�]e�����]�*�Kl�y� ��r�
pfG�nk!���چ��⢑�J{3x���'�>��\9))p��ړ=��v����w	T3�O�y ە	oe,��,�o{ȝ9�|,x��wМؖ�Wl�~�Ꮕ0�?�+f�y��e�W��l���v���)��$X~+"�	���l
�9�=Ƭ�(����<޸O����$(�_���"��}��>c"`�Wi�Wz}��p�5�,y�C ��S�X�-=�� �:[��ܩS��Q�3_&��E����k����/�lۙ+$*���2u�N{�[VhJV�χ�B����v�w��������:c�u��A��6�K(��+ ���=�|�~�,���(�.�Q��"��(ژ]�c
�<�Z/i�ߏʃ���Dl��ЃB:C�� }��W������Wֈq�fC��|��Ss#
T�Hleq�/�p�;tp�J�k<'�X�0�	8��#-cp�Imy!��ǋ� �5��g��������7����������0��i�9ؒl%9���g�� �˪��Kk�6:j W�I5�6��*�����y]{��%��d�g����G@}*��y�o������S��n�6/���t�m9:^>��p���p��rv�2,��z�ͷ0��(#֥蔷h�V�kM# O�e��uYъ\��\8c�b�;�+(Neе�~�q��I1��)�����ܭ F��^���.�K��<π�<��K೅]��㓒:�Y<p�!���+��;W:�� <+S^Gɪ�Wn�xA�9��'���]�N���M�}ʖ8 [�̫�9���R�%9�s{���Z�|�H(�w�~����>���o�5��e� e^&�ضu���&�$B	��UZY����mE�
 �z�k\ !w9`.�;G�f���7�� /��ɥϕ��������;l���b:�W����p8�5���|�j�� ���r��E��&zi)+�Ա��؍����A^RT���ҟҗ1�Q h�-��t���ǘ�Q���<��[���恚B��$�,�v��.��BW����
!��QSL��~3�A]%�QׅCm�4�܎�V$(�.tMD�@�����D�+�@K )����{I�Oڭ�i)cy�>z(�/ط��p�g�+�_�L:���7��%�����U>qr���������΅P9��vO{�)~Dq����lŠl�eh�W��y�r����Ve�����<��_R�46��ܱ9��li�g n%{�]��������eGY��w���j��0�]�߳"��-�y��c ��\�(yvZ }s�c<�Ry�j���SX�\[�@[ey�K^r��^��kbm�~&�&v�,Z��|+m��̟��.0&�
0Ữ�q���E`.�]���^~6���x���D��9.L�����х#d/���{�w���]��΁0������>��Cp��KX�;!x�d��e�}���r�ӆ��-���}�J�QZ#w0oY�9�j �ϯ�� Hv[��<��nt�[�<wIS�1%G������l�9��۫���" nU ]��k����rb�p	ؙ����;�]���4W�����%�/���XMz���x�z�j�*$n���D�	�RZ��&`T9��*�Ϫ,�:�-�n����z���_���
����r�^��.�E*��[���+�{�PڲŘ�c��)Õ]�X������%�]w{B�%@�2'�X�ȟ��L���_�p�<\+W�� ��8��d�vk|�X����ZĒn�;f,M��=ݼ��վ�|m}Xw��e��[��L�;�ow��}H{�5iq��:[b��zM�'�ք@����9��AB�&pb��s���|s�A��{�%�V���H�ҩ�������~�ϸ��I�s��z8�n�}�N;����j������띣��.��FM���W�[��Ȧ��A0N{�����Ա�	��c	���x�����)s�E�)��e׬G�/�Q��f��=�X�YI��/ ��}��tM
<2f�-��8�� ��'�������;��N�㕅��G�Yv9�/��Bc��J����
�nq)A$�g�}?�#����,�z����5cEv�{�Z�Roi�Y����x���k^����9U���8{����w-C�%��_���:f]���|�+Kq����'�<4U����K@9��̟����E;��Y�م�� ��Λ���K;�W^�&V�z�<�3�w�c�'\��k�(P������]�x��'N?��{DJ��xe�^�P��Ɲ�5�{ɒ���;Q�j
ʼ20�g��;@��� �?��;Ŗ5�ת z��P�ۣ��5A4	�^m�hi��]�Z���0&����Z���G9��ֈu��NK��~�7��4������ ��Y�RV$��p�J �:Q�j��|)�,)
��nZV�T��b����u�3�u���X�� q��v׻T $�O��W���kk޴��(�j`�@��Z0\�K����P��|�i��V
YI��V��ɋE�ǩ���_�o�9���{4��=�㥻���N8�ᰊn��� �Ա�8
`�Ի��"xRl��D3_�h	��<����S:��{�KqR� �r�sLj��Y����~	V��]�z���~�t�	���e�*��(��w�9x7DgY�5J`(#�] /[|���ȃ@'Ϙ�^�>?���E���p_3�c�}9��w�;X��V���%��_W�Z��1%�{]��:�z���J|1��gS=`�~��[S`F���:���C[>#eG��jY��� �1�x��'w
�h�S�L�k��Q��"P�{���g�=�{��j�=��g?�ك�].eY륗�w�+l�h1�X!x��H���">�?��~;����3�=�( �k����� ����%%�ă�D������|�쳒��̲����������(��,0V��>��5��ud�§��V�8�j�ۢ���Ҽ��\�T�f%�Z�����jǂ�>�`�������!�Yg�����^�w�Ey�����0ц�������A*L����<m^��Lx,�,P�)W9 �~�
��Y�&E7��%֓z�K����?�m�կ~u�D9����!�U�1�Őӗ���sz� �@z��bxQ9x'8�FQ�J{�m�tTz��©��-y0p�^)?�c�9f��pi����o���0�[2ՙ-=�_��6ʗ#|�xsP���������|D	�s�B�(�/g�y��4^60���R�ښ.�xo��(Yͅ�J�J�{
xNI��86�[�u�i��l�o^�2��%Y@~��n�O%$�B(�qm���S$w[[��c�f+s�6���Sh�ǜr)��Gy%ln��5�SҾ��/�N����e���0����Z�ڮ'�����o�fE�
����4�㹋]�eՋ��M��vh�^uqȍ��Y�.�����Y�5��;�|���m,o=�t�C����:I��/�x`
�;@��AS �j�?�l�e/#+M�E�Q�x���
��K)M�ǧ�c������5��H��o�,�Q���g�q�E]t���� :��'�F����<Z3��&r��",l�zȡ�>k���`�R���O|b�ê�:S�nJ+�O)?�ܢB�e	]Y�,9t����6��`��gф�7)@���Ia��]ih�irJK��7</����ҁ[�S|�`Zk�D����1��m��{�Q�2`+�ڛ]���:���pow�-=�rD]����� �.�ﲬ��ו�	��z��� �4�����]{
����P�o���>/�#@���WF�{����o�x����53o��"=}���q8	푇��TɅ(�	��{����L��)T۶>���.]}��Ö8Y�����p��E?k�Ա���J�
H9eN�q|��HaQߤ�`��]`.I�Q�r� �1���~W:������>�W��=�ӕҕ����V��lY��d� ������u��/gh'�������ϡ�y�I[R���1@�J�j̝�(s5ڵ��x(��-!�������U	�Smq�}?�C?�����!XO��4u1/��%��L�m-L&Sm	]Pܥ��W�1_��F�* �w�2����#pS$�@�SN���^ָH�P�� ����缥��z���Y���`�4 -�I�>j��a=^e�C��[
 ���;��U�@]���o�}�.h��qywf5f�� �R�i#��g�sBt��(�.g>��1��+�����8_�x)o�*+.qW����Ͽd}Ӗ��\�MyPr�K�x�()��4g�o^1�˟7��������1���s'������usk��^=;&��2��"�����I�0_�!`��ʊv��������/|�C4����(�X] �6'ZYV��N��hm= Z��+k42�-hG���U��TVyX_W�B�r�z���p����@��b����'�)����nY<��O���XN�;�np��~�~��3 e�}��>e\ji��u����x;������ּwyty����"C2hfc�>0O\�8�g����{�1뻦�r��1�����a�v���j��Gm����C��/@cd	&�)zg�;B���5Fc�r�ղV�~� F��� ��wY�^z��N�<���,R�觻�%�e��9V@FD�,R�Yn����C��.�l�H�ވ�����r}�S4���ܶ&���h�ܰ3@��.R,��s�AY��.��w��%�V�2���q �S��ଲ�+ݭs�#^�i�re��������3F '��dk����BGA����{�\Yv��J���c������e�U��k�Eۚ<l���
�2Oǒ�4�U���{_��ǿ�lY$;�K}
�q׷�������/��]��b��ғ����8XnC ����u��K������V,�����R��l�ͻ���?�G���pRl u���=:�]tV^=�>u��2Kk��p��$��J��_��� �~�:@^򸔂����.�;E�(�#����ݭZ_#�w���z�)�])��[�js�b�2�=ͺ��"ۿˍ;�]胼XM��5�������rX8��(���:�k��\M&Y��RI��,����S�vܣ�9{h��.�p�[�X�V:����Z�}�{��s��ܥ�������%��"��|�.g\�R�w]k�\r��P�ͩ}=wM3f��y���[<9M�Km�2�KJ {�fy+�R��'ю�i�:����W�_ʎ��Ѻ����Hz�K_cf[ �.�� f}��o����OxǮ�]w�r ;�e:��f�<O�=���x��Ɋ�چR	P��v����`#�ͽ��'�Y�b��������Y~�2���yN�Y~���1�ԒWك�����zު?�S��*w5qe����!;u)�]1�w�=��*�N�25�*�1OA�G!&E ����E�yt=��@�×��R[��%b]��g"���F�3�}뭷.����_ҹ�~���ca冗�X�f���J[���L�W���W}O{�ӆ4:AMֺ�S�����ڻ��ح���Lmԥ��&�S��F�-��ė@��Q�.%Ai�W��WY%a�B���͸:(����P�/�ȩ������V�DMh	��z�~�N�y	��x�`Ϡ��k�v�\F�ʪY��r����;{[�,����vG��4qk�w�k_�r��sCx�5wg8�H�4A�R� O��!�	7���P�h�Y��Q`�����b�/���u�Gitx�������뻾k�w.�t�jgĳ�[�Z�Z��zb8���}�9J[@�2��m?&DZ@�����P�q�51E+�\�vKs�n��_
������������������R���=@-�e�cj[K�Jn�g�f͊&���m��}�Ƀ��Ò�^R�)/[�ny�W������=?+) ��y��Xݭ��Y�;�2?b�C�ʰл�}%��<�� ��c��.��ᥠ+,���̡ X�˩Bh%�^ͼ���Q�'�i���(	�t���J�M�9۴D/_�������^����W��T�%�A���Ξn����=���:�\n|���,]�����W@��\`.tU@ₙ����2��q�J#Z�� ꀫ�E4�.uэcQ��M,s@ �w\����Ѣ���V]nu����� ���T����[���AT4�B�6����x*����zݺ�>:�j��JƠ�]�l���퐓��uӊ��i^���.���������ᮼ.&�.�.ց��6"MM�U=fݯ�b�Y�����l�?}�wY�U��pҜA.����#O%�8-M`�|dy���^����<ѕKMRr��Zճ{�g l��J+e��O� �ZW�Isꓞ�@���j�ż��Pر��7��좷�J��L��r"�ֻh��u0�\�l}CѪYd�'��cA ���w�Z���urw+-�P������A������VR̨ہMe�g�5(��(�G�o�#@��w�5�)�/i<����>���|� _R=-��%#�sa%�g�ꕴe[�u�:��3����u��ݲ~��V�E��ҿ��+��|V������5�:�j1��S�G�)`Իra��MD�A��]y�Kq�-P��,𕋝KD��CiXC�����!^Anumq(���@���p��g��VR�_J�����) w��%�~��;U@�Y� ����U��C`#H��r�Ž�� ��]���&T�tt,sbs�;@���e:8S�pڹ�OY���Ǭ��\��0G���b]�A�rJ����%+�r����t����5^��l�g��ʿ�5_z9[S@<�����7���kg��Z��>����_��7i!�p벎��z ��Z`,�/�#K}Hj���Nw{�y�[���[�@aIy�:dͳ��>�я��i����{���X��,��VV�p�W�N{�ƗU��zy�P^\[�`��=Fꃃ�����7���R���&�\��h �\ʙ^�Ƨ�g� }�g+�� -��T��������P��Ю(�+ 䩍��η�9���c^J�8���`�5��Yi��Q28���
�j��))��l���������������tX��~�ѯ?�IO�G�S�ߚ �s����'��7�r��!,��J��1"�0'J��#�! +j�<iꋄ���	|�. �� H���r� ��s�Y
������ew1��Z'W0��^.e�N����z�ڻ����\�"�R��b�MvZP?>���/]~�僷�5�ڲȘ�2ӵ�t�:����'�D/yDC V�`��!���|z���|�}��Y��e͒�`������u�R�� �T���ӭN\�X�YIX���K`�A1[ܔ[������՜���c@]��=OIa���k���-@1��ܷc~~%<���l�Y@�l�[.���/��tv���r���D���j�`!�ӳ�v!��X���\�Z.5����*\�"k��pǂr����6Q����b&�p#\p+�\�*[i����]u���c��g�Xnuڨ���=nw\�j7@���Z��g>3(�ұ_]}p�b�9M�
����ٽ\s�S7���R~��R�'Dtt%R��>�����R��(��!z�z���S��pk7[�5>CQ(��x�{�Iid�P��L��Z��k���@�u����S��ҩ��d�������%e���:Z��)��r�c9�ܚ�њ��������z^���\Gi猎Y<��Q���~��#h�ڲ6ȇ�� �oD@�c_�Qǖ�/�֞q	��jk�ֵ,W�E��
�p�'�a�`1�&=�^n���>{ ]��U���E�H!�#+Zk߲����H�����*+�;��>�8h�M�W��H�mT���š/Rd�
lX���-E�0+��S��N��E;�Q;~�.L�D_�L�w���G��b+A��9`1ƃ2 ��7 �]� ��{��5:f t�b(�&��[��](����t�Wjx������`Ͽ6peC0��=!c�
h�֖��f����=������$ ]W�.G��,/ ���)k��}��@HPHX�O�@W �A4����� Dֺ�XQ�c8XF@��r��6pi�����O����,�/k��/}�������\u�j��u�Q��}�{������ �	�� |�S�ڧ�)?�-
2�=��j��堮�J�k�R���+E@�ߔOi�D?@p|YV�rev׭���lQfZ�|Qg��{��\ـ9V8���>�V]s��w�g��,��׎��t�卹�͐C�>��sw:w�Fr� ]�?�ϸ3�S]��[�gzI�	�4q%dY��`��$�!I%P�_����\�)`��^s��5qY˲ص�.K\u	td5�������Y�Ǚ����Q��S�����&�G��,"�Y;F��w�#�7@핲!���+��%�����.�J��Ew�s^���oDг��+?g/���ROXC�ip�5�y:����X�kY�>}��}]=��z���_�y�f�{�SdΔ4󴫧]��%N��H��U�,��ء�}1��s�%��c�>�W\y�+T��$|RmLIXy(�w]KX� �֚�j��U^m���?��p�W��%�Z��60�*�[���Z���\Q�ZW?�3Жk��\�Ջ�9�������{�7
�ʰ|ܩ�X����l�������M{C۸Δ�K�fSz��Wk�0p�--�{��] �vr�*Z��_>Y���s;p�s��˳��^�8�u�]w��8�L�^�m��5�7��ZC/Se���k�n�� Q jk�އ�(�h�ӽ��'�5����-p_�5��k=o�
]I��Ւ�2�N����;��űe�������"���y��B������n����'��۳�@��<gA�#07�!����q: ,7�h���*����W����^��e�k�]�t���˥���0H�Py���.��������:7`���.� ��qU+�T*������������9��q�����>ky%E4x��!:��r�A9�o,Ud�3�9�8��5��e1��-��\�0�X�9- X[���Ͻ�K�LM����e���4*ѳ%�Z4�ϧQ`�K�
3gŸ����l��;�kM]� �;�v0�If�(�/i�~�%�L \I�ki�-�oʘ��X(�LmhjZ��p����X��*������|�3�b�hX[ז7Y�J#:����8p	�s��{խ�(�^yd}J���pY�9)8�V&�D����5�,o��S�Q�x�h���KQ��UM ���C'�]
�*���q��Z��E��5�e�o���i�e��jc�Aq�K�^Z{�t�����@Yp������x���Z�y������3r�t�ݕu~Q��/�f��a�ybt�j0�+^�oX�} ��Apm)x���z8p�uf��_�5ث��mY����S�,:jT�H�8��`�	T�.e�Z���d>���H	P�����"Wy\K��p�
�$�T��������pڜ\�R2�p����Ku��R�*GmҶ6�ծ��|Jڶ�m�.ZJ<Bj,lx+��w��9�c��y�W�;�O�1�0�� ���-�նE˛�/+��z�ކ���MN���#\����_�Aq��v��kn��dqؕo~��� ��}�ҥ4P	HMH�MH��������Բ
�,��u��l��)@��2)�xʅ���	t�6��,p�hY���'0����O�u��^v��/����E�ѳ���:>V�t��]m`{����(�>��E��H\s�5�����g�L�,�[J���	��@�Kc�E(~M��pd�<��h�:�@\i�� D�A�ndC���rh��޳u��^[&y�s�$8_ӆ.��^j�~���Q����<���܆����dť4���o�BQ��T��HS�^$]����� ���9���{)A����-d�_��W}&�^��;J�m�
����� ��@9@�_� ��L̚�����K5���[��, �a��9��zW�	p#hP@#%@��X`�@7ݕ���Z�M�]�0i,T�&����ZW9?��?8���W^��
U���o��ל94��/�r�Z�\�׀=��}E�Q���Qv��/;��p���&<���S��T�YM���*+���2,X��7�d�RG^�&mIy�@����Z�%Eb��r9�$�r>�He�7\~0o�e�ٮ��_�E�%������.c��M =� ���o�>��/�?2����HY��Fi�k�8�C�F��:U��" �r����#a9_]�hr�����.�vJ/0� �馰g=�Y�)rJ/��d>�Y�l��<\e��-o��q�C�J��i�X�gg�~׸�>Y��yi��Z�,1��}�����C�
��:BF@.K^ �~���.��u.���++!�o�ʬ�qW��e����[�(�K��iKc������,���,ˋLߚYj_��Z����~�n�;�ݛ��{̵��yW촹2�Ͽs�NJ�m�m������ ����9Wsv�aMI(
ؗ�2$`�^BPoM��s�֖���v����ek�����߱��Ա�Fi�r��r�kۛ>�U�>�by�ڱT�ȍ/�@e��rT>Ǫ�v+�`d��Ƙ��L�y�1%}i��ꀦx�(wաtn��e	��x��!zN}�f�	��|��VUFv��@�����P�3�� }��]����c6�0������1Z���Ϸj�4���Q���ƐCo�c������%�g'}'Bm�?���pʻ���_��^�~@i��[#�p��0'a�V�<M���=B�RS�9(���qы&bz�ջ~�Lv}��nZW��n�] ��i���%P�?��s'U� ���`8�N� ��a��^���׾������K�޺%FK++p��-Ū�q�y���W�P�a�k�h��.�^��κ;�R�d�+XP��M�w܄��s���y�d�c�*�\w����}���h܌6�}@�F���cV��$��Ql�w�)Y�yގ)�%%�&�ZAK,������[�o����վZ���::����c��+�2�����C��~뷮h�sgy�����ᶽ9���	oς=:�s�BmށAP�w�qA2o�k��6�=̀��\{̹L������볬f���ƵO\y�W�� Lּh,�[�Zl��s���M���x�;���a]��/����Vt+����R,1h�{]���p��g���*"�E�Z���HɑR���$|3�e~�ZfIŭiS�<�&�.R��(]�9���K�c�{�3�}���G�>���-��׵0FPx}}ܕ�Mg�E���߄��������b5���]���}q��G����O�1(��4D�{K���l�s�K@!%G ���c�'%A .��@7�JidE��}�"ѵg�S� �������U�.��a�^��ǘ�� ��Z�J��
�b�;�y=�}鞆��J�u�(=�����[Р��h� �۝?뻃9�v_��r�.Y��J��ǬG���u�<�{۟H�1�n��Y��<�3�؇��_��^������t���UmX�7Ś��{J��}-�604}2�J�'¸&[�^>cB�U�"�U��@�#����y�Y���, "��؉Hw7��~:�E�\���k��qH��-.h���ݕ^w��L���?�7���3n� �'И�iDW�fBdH.�c�O��+ڊ�\�#��.{�[?���e�-�x��ju�.�1}r�,���G�:��f��a��\���_��
���w�*�����Ӷ�����g0:�w?��^��2>�c�=��H���s�����Gm��6]C�1?�S?uZ�n��$|i��/��ࡴ=ӀK��ҕ��ob���~���E�A�ځ7Y��ga�v#0*��&� � .h�8�L��o��s��aߺ�p�E�r�f�g�[��Z�N7�}��}�pʜ,S��������k4�j�2&S��s�.(4���˃���2(��	�� Nm��t��H��AA�#[13p�f��yo�C����Aރќ���"��{����{V�Jʆ���w�1夤T���\�s{Q�5%�j��g�������&j.�;�%��;q��C�1b=�2�wc���G����ÎT�6��E�p��p�%��E��S�O��	4���E �}����Z�s,S�6����W��$�q����9V��Y_gۙ�Q0���v�9�+h�+C�~�s啢 k]�st�{��ޥ8�w�u�{���P��y�8���r��2�x栜�x��XxR|�x���E��*��g��ב��>�X�1@�Q�c�����:�Tk:�y�Q
��1��*�Hm�nk�[-��Q����u��<|��!oW����D���o�����W��W��ԇǌ��v��ՠ��O�����{e�AGHbMj��~�*�A�3���>E L�0�н^��}��a�80h��wF��['�I��׈*���0��.�A���hz�i�ݘP�W�N�СK�x��d��Yn���K��e瀀Z�H1��� +]����p��i�~�y��,r��d�oe�F��>���������yWI�Bw%��k]��
&�ǔ���}�ߡטB����\�H�ԏy��T�75]�_T~���v��3b�X������xgȨKB��a���_��_�~j�v�t������z�_��_yYXx����!hv�rd���V�D�ДU�a(b	(Y�b }F`�\A��F��(?��"�Fh�\�5%�͘t(ݺ&k]tU ��s@_�䷭	�U��.t���%�Z���e`�:�9_�Q@9�$�oR\��s�=��@Y�*C�9Vt�tͭ��,b��*��{ ���u��m�Y�م���m�sЩ?���٘2�2H���Ӕ:v�4��Ғ_��-z�zp���;k�(l����� �{��n�9�����!���s?�s�l��?�d{������>��!�~0o3�[@ Ћ9q�㖑�(�b�%���a[b{�oLc�"mDWY�rє�X�zWzh+����������o�y�J�U���ٿ.׽��U~?/`5,��x� ��Y ��D�s���t�F������턜�(I
��#�Zz��-�>Ղt�V����W}����l���٭g�)���v��xn�=��z��ͩҳ��-��h�t�ȍ�|�����B^��v��/��s��]��/���?�+�?�������k��=m^>ٮ�~�E���w���c����$0p�{�����kz@�jN��,k��YIz&��H�� ���Mm�1��J���#�u	�em���t����sa�.ra����3���`�K9P�ܼ
ּ&�oY�д�C��.�a���?=ӿ�)z":�`�����~߹^u����Z�̟�k�k.��ik[�ܚ�6e�AVB� s	н�1Z����6e��S�Z��z�txS�X�X媛�v,�x�F�֕1��<����f�{���O����+�����˿|X\����8,�ce�9������WV��Aغ�hM��9�͓�q	��0�:��	�I�w���g]��e�j]]@�9�J/KT@&�K��@_�kޟ>� m�_������nj�tX���#@0s.��J�WCt��q�E�Ѓ[v�dk�f���[b��׎�̀��� �G�)��˫�7�_�z�i�d[:���\-��X欝#�gy�|qsȉ�l��؎����ٟ�sZ�z�L���j��~��>#"��c�sp��עm%H9Ɍ-TZb����-�X�2�*{[=��!��N�Y���OjR_� Ȣ�Y7��:UNAsڢ&���¦4R��ܾ�Ǳ�O`��v��������.U�̉%�o)E�3V��'���~_�ց/:v�A3�_c�]�ꥌ��<�%��x.�zj�bl�m@/�s��՜�V�lK@�v�_n�������[C�\��=�|�3?�Y�GKw��
�c] �����?������?M֟,qY�~[�����g�V�@,t_K�)+��Λ^����������%mM�u��dQ�K}�Ҕ���]���t����tY�{�js��<�E�y�ע�[.wO܆���)E�g�Y��@M�.o��QV:���?ƛ�G[Ji	B#����2 �5v��^r�gZ��hƻ�l;_,:Z�Un�y��Z�[�k���ߪ�U~�9��\����7[d��!j]<2桘?���X�{g���:��n�k��m��?oS`��C�������o������c}��a��a��.T>�� B0�$���'��b�6�v�y��nqY[�5	�s����}.:*�,s�����ZUY�u��5����v�}ǅ(��?���;At<��U��@���P��[�57[��x>���w /Yץ�Sd�?�/��>?7��q���x}����HwGȇ�b��M�)����]��?��}�|�~] ����׾��pO�-N;3�`��{}���T8	 YI�Թ�����w���� .��(Ѝ��$	�݊�pU-�\�
��˥�-nq��h[�~��d�����4Ղ�Rv)��u��=p��d�wv_�w.b���&%Iֻ��6�v������T0��aQ��9��,tsQ�5�^9>����k��{"��O���Ǳ���m����X.w���{�;����$��ق�w��s��_P�2�˽d}8)p�qk �Z�ZVf�p����X�r�x�R�<��T�$@b/�� q���?���X\{͵K7�t� �5A0���͟ӷ\�����ᣜ���]4�2�8A������͐��4:dF^h�5S��;���^tW�r����Ҽ���2~�Bo)6����ߢS��V�V���[ϩ��RZ3�=��0��p{��]�ở�\�����7��ԟ/N�u��F���q���r�پ8��Z��FL#�b�>K�I��]����;��&�T��V9S�[�tޚ�q��g��,u2-L^�-R���J�u�uu���Z���Ҡ����O���e�?qb���~~y>$Ը�υn�#��i�rK���Y�:_;��F��^
~`W�9�u�BR�ݕΟ�����ֿ�y%e����<a~���eH��x8�㎐_�9�g�}�s?{�o�����~��JkB�u�a�����D���/,�������ѡ<�X����$���J�9Z�j�g7���.	��KB^��p�	е�\/H)=nxY��z�kk��������%�Z��Gup��~w��]�e���|H��>y����v>��[�f��7���d)��ہb�o%�{N_�)�^t�^��(M��зP�����7���2��7�"vļ+�v��_���S�Vʨ�;@W������U��c��Iޗ,8��8O[�`1��@�Y��Y;;��~�����Ж%*O�h�����gX���\ͥ�T[�ŷ��`n��.\���	ys ]t]f.��5s���C�#�n��gf@v`���v���s��B0�cAo5��^��R~jYح�[�[����O�гg�����o��9��7q*��|�K^�ո��;9ۻ�;I��&(���~�����E��H��gG�����]�R�&�! ����cJ�F� `��-��"�<�����uu�N��?���%@_o����y�[B\t�8x�s ē���]
@���2��4�����7ڣ8��v�Lm�[�K�&��� �[��>��{�?���V���|;0Ѻ��E�}�C��?7.�?��� _#����)W�T`��/�[�y��%`�-�����xw.�Ғ�ȭ��ixbDg,B�^4�" �s����%4Z�)kQ�b^��<6��������y�XK�.t���� ���lS\��υ���V.��x��]9��m�9�����o^~���ŗ�M5�����܌KH:涘럏�طǁS���n�u��uz}ߡ��t5��o~�����}!,��g��J����gW��.&ص&,�A������t�n�F ��������J���!�s�U���s�z�<>���2�	�9O|%RiTʥ�-ăJ������6�}Y�6�n���k��k�Cm�h�uG�+"��G��7����<���~E<��8���F~cl;�gG��؟u�"���ƣ���/�L|����N	���̥|�"F0�+���:f	�v&@�@��ȸ�MB@�%��� ]
��
]�}��m~�l�v7	J��緯��,T���-mUS9%�����ޑ]='^e<ߎ��r�����:��Ǖ�~�|����~�F�����E�W�����6�_�� ��`����&� uܾܵ���2g��[�-��eu�����`���`�u��hX��Y/�1��V��X贷�z�k�q;�G�E�}U/{�������C�D'�N[��`m)�%@��s��?f����S]�-Zn��k��Ȓ�Z�9��ܶ(����nT���
���⒦k��ۧ���l[
l@��޶�;���}�k_��������Kk��lk���ɉs��J� /�a�{�6lSB�V�-V* @�]�傗%�w-uh}�oƛJ��ҧ��>/�r95��w�������Z{�8y6ă���CYA�����
`���e�C�$%>�����ƭ��q[��+��nϼ��{� �C���{��o�9��X'�y����k�q�6��ێ�2�=w�G�G�kV?��N0������8E��s^	V	Y	Q�sԩ�-UeJ��6mM�@j=oEU�X�%0[�[k�9?H�.`��%{�9������E�V�%��:e�z��[W~ڕ=@�o�Xrr�֬�Kt�[}/=oY�+��"mڑ󬔞S�I�����ٱ���<yI(�������/�9��{��:g�a�C��/�����G�V�O8�,�  �Cf�g�H�:GŪ\	H����PomjM���N�y�g@��3?���Q�z��C�)Y5 ����y��Wh�R{rz���)/���FR|�>�q�,t�Ξ��a�O�����
i�Bo)+��V��-?[�[i�V������μD5��x��-��W��?�c�?��׿��z��J���o
l(@Ibk�)W^y�υ@�ް�҄ K���"�I��eUr��ޕ_���U�Ήs��hM���y�61���j����d{  ���X,J�y���w���;�ap@W{��]|Ŷ?�\/�v�����3mk�n�:���ޢ��y���h��(�S��)�����#r��C�^�c?�cw�����6���]���Moz�3b?��������r#�<�!��I��:�S�q\,J�(�G9��c@Z����b���o��Z�k�_�������rϿg��~�"����w�����7�)�����C�h��?�.l��|oA�������S�t�kؽS���V9��mͿ��Z+@n���\�,��@T"�k�I�x��4�]71�|����a�ֿ�o���o-¯��b�i���?x�w~�w�{������ψ��1��A	�>3��54�%p�v���*� �0��Rj	�u:�YkHx�l�_~�.z�S)��$W�0yS[��5�V/z�R�#�Q"[�Ԓ��V��B�%v�|6X� �������<�*�?_��p:���_�����ַ�,�_����'���|�=����\��r�O������r�7��-����:+��*�X�v.����x-j��BR��;n���8bW�J���D��ƣe!O][o���v���������F����Ms�[�s�}$��r�s�{o����~&�i�9�yp�Ƥ���(��,tH� ���_����_���1�:�O�g�$H���'ui�iv��u���%ЖE�<XG*��m"����}�-����)�˝z<8��w7�.��Km�>b���6��- o�TW{�M���e%iZ���w%u���R�B�!��q�]wE�����w����#?�#�D�[��t=�*�a�Z�����t��_���?�����r��JPK{mi�NK,(_g�s_;�g,t���D"���l	����<}+ճ�����5௴���%K�AP�ux��8E�비��J����;�i�>g"�h�� 7�k5�[-�\�rj}nr��Z�׺���[�W�K�0QZ�i��(���ߌ�7F���t�Iu]'���ЦL��f���n��>����dlz}0�)X�X����	$�F���	��IJXZz�@��x�?�Ӛ؋�M�?�r[�[�n�o	�V�Z�[��4�5O�Љ�k�Gt��Q
"����^At�=�ik۔%"L��}��h�o�~k��ȭ��w�Z�/ʿ5@�쒁1;���[#�'�2���~�/G���-�������$��?�����s����!8,�� �E&��&+`b���͞v"���H�&��e����5�p��|$�b���
~�5���T�����oS{,#&����UwD�����g�}4<�7�IoO-��ۘ�!,tH��W���K/��_���� ��H��%�x��E�uO��'N��@\��0G��TK�&��*"S��س����SAj��Ӫ�U���5���\ �.w�D�4BY��'���t=�HV���c)�����j}o�g{?�Vz�Ϸ���Z�l�=ﷅl����~w[��'~�'��=��n�q��o
�P�����������O��g~2��ׅ0=ѭ$Mڼ�ݚ�<�KǙƃ��
7<��@Ԋ`�Y�ر���L�E�T�V�+�Ev���Ω��E��eN>����v�(?��*�7����.���Z���J����������Z����X���Y�/����j^���o�����K8���Ǵ^�3?�3w��}=�Ƣ����/}鱗\r�?!��:"6�}W��i8P!�� ���!�2�(����U��^������E���t��~-���=[�зF<5�l�,:��p�P��-�n|�V}��O����-�.
�-����[��9�rg�>�9sSȤ���W��_������Z���;&v�5�<4�7sC�|�?������O��=�����#TZ�o=Wd��\�N��3� �Q�K�ɧ�[x�d���W�@)�?[.w.���"Z��A��Bn�2Eü�E/z�g�o~�_����k'��i�3�o|����W�d�g1�O}=kM�/8���V1��b���q�b�s&<AQ��-����mY�k��-�d*�-j����=���|�_���?�
H�����Hw	(H+��H5%$�Ew������9�a��ۨ}����>����;���y�u���ڎ��T8=�/�������hܑY.C!���m�u���R�2Q4kl}��nڱ�����+,������b�8}�sx����e�R��]�DJ+/Q�Nq;�}iJ~����/��*�C$��,	Zr��,LgىR�U>	��>�n���f����������.�{tu��
�������7��KO�Ɏ��r~�L_N��;D��z�P�̇�C����F���&�>%�F�W��7�-�;�a���VBĎ�ӆ��8�R�����6��{o��~�����W}���O���ׂp>�H�6ۛ�e4� ���y>[H���qI�q�Y���V���M��*�*l��3ޜ|�$��������杝�*�5vY���Q�� ��&°��d�W҄؟�	�B-������ ��":+�5."�X}�v��=��|�9�q4��6�n�O��$�nT�W}���XOi;�������+�:��
��Zc��˫��ULҪ�^�/̪ZV��9�f%�W�v��X�c�w�c>b�=z*	��V)�`���w�`�ek��&���5đ�+̗mBO��cG?Ă1$)4&m��=2�I$gy���I�~Vo� -S0i`q)i�/Ie�\��.p(�$�����y^� �\�����;��V�����\���ަ ��R���O>�/уP�w3&2�a ���s�lTP��@�;� ��Tf�/�֥*c�j���oXu�Z�-9�\:\�2��.h
����$�FR������'�h���g�|��؀����rly�q�Uȿ|�+����|���}@l5NU�h0.���qM��h���kR��W#A��-mh	f�sK+@\@��D�^��q6��-p&rjU���������Zj�+|��p�F�����'uJr����CS����w��I}�w���&�õ^��!��gz7E����ڻ����O��;��Ұ[+�	F��S��©�t��������¼��y��u���6��e�}�� �(�e� ��H����,?S� ��!���,UY��%]��QLM�)�iۣW˞����7�s��Ts('Ѯ�1������E3�a{ٝ֞��W@WD6yW���|�k-�-�s�a'�<�סi~Z�n��>[���v[t<��7�_����'ҋ�g�i|�1�*������Չ2�n4_އ�:��Ev�GŹ�V	4�I�K�F�F�wVܬh�r����ט`y���dbS�ן�0˃�{����,��WQ�*��'1���64���v���:����!͟���lN�\=\Sl,��[�g�_�q)��fX_�f��7U_�B΀�Ҥ�n*p�o��*���7���g�P��!�VK#H�>�"l�$K�ɧ�7���f�8��(rź�����})?ڒ`�0,���8�
�g�#��T���~��g�E��=l���O	g(q6�o�<�"٪`AZ�����P�v"W�TЫQ�y�#í酾�e4�#�W,Ro�����]9�ޫ龅���FN�d��n�q�M�͑�Sg�X����(E�S��HՃ	n����m*b�(P��A]��"�}|%� =��<�3���/�������0k��	����KE�}���쫎��wՐPO�V�+��_���K���C6Zw���]�k����[�Ȓ���k�~W���O�TQ��F��N>-`�n?�\��,��#{�zU�C�����@r;WA|	d�&�ȔsG&�1JE)��o�� �:I����?�1��ѫ�qLA*�`	Z�-����"�C.
Öq��ע��'73�T�H搨��3�n�Q<v<� Ǚ��z�И���{�E�X�.�D�}����4S�M��!7G����6<�e��N�������a"�������B���^vHږ�!�xl��K�R�����/Y7�J{�㗛*lY�:>�e&w���>�\��Or��~�u&�wEn�����R�8�:)ٔS���"��@��뀪0[`�۲��)ڰ"|��W�X�Ar��jI(7�����Io�$R$%�8����?깝�?
��$���ie�M�M�}��j\�gWޔ�7�G-�;�5إ�[8���c��N�����V���+����8�%g�I���aD����P���[� �/M�O3C����$�6V_�N�i۴�f!h��$�_\�T�!��.��5j���M�����G�=vJL0�OB�
�`���3w���_����1e�~c�1���>�a5�d��.H�T4V� e�:��ٹ������T-̏0������v�ViG��6��仦���x�#�9-���tpk3~����V{�(6e��~uʇ�}�;���:�6{�B����G�w�w��c��% b9�GW�79]�y����p�*���W����n�;Y
)�a�����U�=����1<�k��&o]R]f>/���ʧeJ��%^��nt97H�,���9pe�����T��l��A���G1;+ �FCO$ ��VC%���~���$��}6���
���Mu�D˭�y�Wp�7��cƏ[�J\����;'.�yp��R�hZ�9�L�u����z��\]���݂v���#��������P��d�'��9�FQ]@]y�M�JoUpP���c|�M����}��jf $pdp&�Ԑ��%�x2�?m>K��ؿN:�NY�!l\|c�	����!���@���#gT��t��JqDk؄(�=�]�!��V�0>-�Ɂ���y���o����k���t/,�z�n����3��,�F�HsE�WW�j� mdy}婉Gle�"n���|��Qsc�m�5x7�1�
N�V����_�eq�~��9���~�t�n�?̤l���L��2f�c>�,��=掅����p�W/;�4$�b24��>�ֶz�"�ϫ�[Y�{�Ib�O܋�`����DK��4+V�s6�fH�Ɣ���(Z�M�r���7s��j8��~�Z^����3�k}���xp�}��I��$�!��XR��C���gKk�g1aumό�8A�#J�(�aM�/���DH�<�,�s��`�����г ��Y��Ï��|�7���'�>��[�F�NMU޶�����(�`�"���d�O,~�6g��|�	u�I���<��.:�9eec�<��`E���pѸ�
�A#5oc��7��S� 8��&%��+k�#��'-&-A*��JM�Ϯ�G8�<�M��%i߾�����.2��ٱ|���H�"����7"|��9�V�1�D�P��[4�bY�z~�4��'�}�)C�٬?LB�A��Hfh]�d�$IZ�kI����ח����,R�bKR�Ϳ����ש-��(��̨��Z�l����S}�(F+�z��(_X�~Xo9�cM2�Yd�T-fn{�+�!$�P���H6\4����}�`%�WX!�b�aN����E���x]���kG�׻b����/�������=���I��4�J�5�Ԋ����~����y�ص���o�{?����}���yn2�'��0U�/�/L��� �u����ֿ�������Zb��{��t*��*�`���H9�bݯ�ڴ�:�\����R� 	�{���������N�w$�#e(��Ԕ��N�5O���$�Y^�K�F�ִ�Sy��5Q���v_�[�2�ۓDc����%b�x�V?�f��&�#̡)��}!��M�q�|�^��1 �VS��t^��E��dQ�N#aj��}!lV;Z���t���_�m<�,/{��$����4��᱂�	�X|���L���|��}�)�4��,���u���k�8gh%�����A�{��O����
Q>n_�]�ۛSr_j�����2�,'�z]w�ŗH��;��n�%�'�>զ��,����Po����+&���V$Y�EC���q���̈́�ŭ�0+g�Ǎ+��(+��[�oaS����W�!'e��{�`�_�*.����X���A���9�f�ԊU���or�vz'}���_
o��~�yt�|Q<&�;�w���LA�u�4�l���k�z��q�� ��uT����΍�����BD���p*5���6P�հV���k؛u�t�a��!U����d��Py��ک�;�S�ER��a�^b����TH�G�wX��(!���-O�y1�_ |k��J��KƤi�/��7��9��/7se��X�O��X]��������Xc���<�tӁ9�"Q�b�	�Vl�{��0z;夾�#��m�Qs��ԙ!��_���|���Z�x*>@s���;��/`MO,�?1�t;@`S��I��*��ݽ�
�W�^'�F�`~���''pl�
�� ���!���f��&�M��ŢwP�e�t������d�Y��2��&`0�>�zG��<�_*Os��Yd�5p.o �8�1/csZD2�I�M��ۀL�we@6~���X+]�!����
ꮼ�?�|օ%U��!��+��u,ݩ�,��y4�n���]�0�I��؎�3���ߣ�w����
����U��v�W
kʟ��C�܋�6��EY�k1����A�|�5�3n׊��N�z􅍛SÙ�@��Rs��1'�dOzg췦���5�"�Ti�rW��g1e�����S�&W�qDA�����-��#�K?�F�ct%�H뚓3��b��0����u��ҩ7W�^��(�;UN�X�4Rxvw`e��R�EO�CI�0�Ǜ��vh�����|t4�����ۜ��ڡv��cO4� ��$h�9*���
!g6|��WZX"��]qf���_�6�q�1�l��7c�ci�?�����њ<4�����S�1Щ����5�3���O�3��n�c�����u"��JXg��101�<�@�C�@H��1I~��3^�o��O`:ktg�-E��m5m��GܭQ�i�΃���9���_�B�������	��Aꈚ�h,�RJ������Ƒ@@U����ק/޽�ߏJ��u�f�+��^��o�oxq_��"�ya-�w�E\(�3gD[��p��B��25�����D�m�#nk]���B�eWm���f���o���j[��U�u>�z�ˣ���̈2x�&�?eH�V��n��vu�~-�@5���!<���2w�r�%��{߸�m��ێ��Q3�N�NH�[a������ِb��-`C�9�UY8�J�a��^U�xQ]�FW��a{�WU�Q�s�Yǈ0,��{����ֆ���$�.�[�Ti�%�+�L8��g�v�in��b.�*��P)��G�;ʻ�����ܺ��R�獊�((�KMq��fOc����XS�$oD��/ehu��^#��n#=�Yi��Jr�~Z�������i��δ!*�%�#�E�����nU!�!�������V�uE(�'�>GR�ěR�na�"U�}:� ���h����ԜAԬ��&O����|�'+-�G�#93_];1"�����Y�_t.�*�K���W�S�[}��ފ�wA���g���7S�6����j�vm�o��_�iC4�f�{ϣ�]�V=VF��bBM
	����F�����oL>��Q�a����r5��W�;�6ַnF�Ԩ�!���}��:���6�o��P7!�DO���f�^gm�˷��5�lv�~+`�b1�/�r����.Ŗ0?e�SS+�V}��K�|hw�L9�(>����~4K�W�A�rY+H��C����Wݿ3KWo/Z:M*�|ė���b4&�>gAQ���bJ�u`�����P�W��j�S���(�yi��J��ǿO�
D��y�
ޅŞ��E�$X"�ʛ�ͩAp���8i=% �ش6r�5���X�U�%q����Q��!�r�1�:��ܕne��\F��&�zn��?�.]^��˒�ʨ����4?�`�����A	��/�OE�3R�T~�\�sݬ��� d��WpT5�!��P�Iu�,�ƏGoBR"���ݹ�|��n��/\�ғ���l�ڕ������y�ֵP��Mb�#� L�A�%�#�"'�����&�������)�Z���I�U���>e
�KWP?G��������,?e[��6�&XO�g���]�����Tu�z�r_� �ڪo��\2�|��@�1�3�C�#�qB~�ب3:�J�I��a��N�������Fg�B��/ޞ�w��Xdw�VIz��^T�3KEG�zXp=�r\A��6��J��c�?c!ng4���=,�r�Q�~�P!ԸV/�nu+A�]QCzӰ5p��;�)�|�N�6E�_q�aw}
���9[�0�z����;�XW��5܎a<Gr�1.��u?%�0�n�'��@�/�1p"W�}C�6��h�)+a6cG�qR�JC��ZV���������B��48U�,��?�)(�R�/�7M-�E��E�4X�%����U-���D�Q�*�!��*K��1�e�M �/_�9����M���K &���5X04�$��Q�w*����V�$�/�?�N�۸"=^!������D�n��gq�Gu��Fɓi��ȨԔ`�u��b���Ս�)�I��8���h��C��e�\EL����.�FBf��jN��7b�$We_f#ɭ,Y�A^W�\�G�5�R�K�M.].��ERN��:_."��K�9 >>��/̠�:��@���ｮB���FUr{��g%�U3�Ȕ�M�ѲV2@S���X����t�h��߷%,����c�h��C}V��g���̦�!e�6����Gp�������DJ�41ug�&={�D��bIk��9����?Ɯ��i�+H�uT�����%W���S�!�яU����Ԣ�["&}\9z*A�mN�G�{y8 4�sA�(�-�B1��O�q6���
�w\�᫛�w�9����?�P��&w�^tk�V���I��~�� ��}$
,�M�����5Ք=T�ߐ2�e���!+J�]�2�}I���O�b�j�$US��7��n
ߺ�}���~��wu���ދ�&W�DA�X�|]�h|N��T��w�-h��X0�|{��v\�4)M��T�[xI��$���	��9B.E�m�z��e�����A��H�{ΜI��&�.�𗣜���F[�=F
����l��ޅ]"�������� ,���s��Y��e��gE������ŲT�l��M�$?*�I7<E�E�سT-��d�CFec�Ō��fMʳ�;�2���\=�?����4{���Qf��5b�6�j?��Ѷh	k1���2G�Ru3���*<�^���ր�=Lǒ�c�����0W

��] ��q����-n��>Rn�ZLzv�Ď��-M��PaR�Fh��D;��>�	�=���D"�)��n��P�w]��Iqo�S��TX0����DgX�6�5���ڭ���T�~�WQ��<���Aby!{=b/�E��Ζu�`�{{�*�-zy2_�Fo�2��s��&Wt���'�����.�	
d�z�OLj�}����r�PZ�׋zO�&�V�F�ԗE�}yoV�,ND7+ǽ8Sf��k�ͳ:��ԆM)�/@��ZW\�����󣥖D���t���WS�B��H!�4aJ1�"A�[�����,�U�T^W�ag� }�d�R�O�u�`��������
F�� $��g?o��Ae� #�B��,��d�l��|�_CA��c�ض��à�l�At3�����ec�>�����ˊ��� j�-�YGف/�$�.O�G�U��G��I,��2:�,��f�^c�l�(�b�� Q^�� #�M欼<{��x��8�8�@�bŊZ�ڴ��x�o�^%m,Sڛ�~��evuS!��z�B�c�_gJ�+�WӍ9�5ƪ ���Gl��H�"(V���H��e��D	_Nc��T�9[r�w�����;�Q��p���xlQ���`�H�q�Q0��QB0���bjy�kTs��,�Q����g�l���a���iE��9�u:���ݞc�8�G��y �ښK�m6��:`f�{��D����>'�ޙ��hU|�>n�~�X�ϑ�r�h���1%7M���j����J�x���Y4�:Xݺ-ja�,�;�0Iy�٪统���;*V��y&Y���a��D�Y)������񩰫�0V�ۋ�?��&����l���^H���Ǣ���r
�����NłA-K�������ܭf���vc_�u3��	�P�$Uۂ��=4�tvZ����ˡ�����;�#6X�wO����>��c�w��(�T��݇��p,;�q�}x��v����B��
�1�Rd�	{��n��?�;����x֯"f�kQ�T�7�z�\%fjK���6Ln��cjZ6]̳Rf,�.i
�#���0>s9���'�s˳vDk䍈R��8Y�YB4�0A�b�=���7D?yMi.�j�	�/?>��2��q2hMLvcZ���Gex�)zb�a{�k���w8ߝY�il �����-��f��֡���,�E�Zq] U��t�.�p�ZS|�\x٢�d�b2��"���4�D�V��.�9�#�a��n\��C��a5L&���62o/B�vQ�]ph7��*7�2-�},��#�;�k6z�iQro�It��sH��%ӈ�0��T{�H��["B���0b~���m�ɾZ� R��;���)tf��=K����(S>���5Q����O�H��U ܇�)��Җ0�P�uѽ���Y̝�[.�Ԃ�� ���*�3:�,�ȓ��/��D��H@�j�6����R˺ ��k.M�8�\ܨ���9���դ�B ���z��Y��(��ϓ]ϳ�\��(��J�6��`��iF�k/�`�w��u�->��k��Z7��us�T�V�"-��&�Λ]���Œ��S:��Li��������]�{���e3�+��4�9�C��koG���x��h������Vfv��Q{��x��i!�����ح�ol/#al��X]㤽�������_����l�&Ze�0��	�9ل�����Xf<���N�;�̢XT!��*�Hl���7�a����W]��I�.b�:ỔA�S���sʿ��5�~�_�����Lgf�؈bP���BF�����w���!wU��>%���T�������@����K�D]�k=Q4 ����e��/{@6���@�w��'��G�	��W �m�ɴ�
C� R�����h�lۚd���躌lw*�螅I�oI��xPq[�i,d��@�6Y\/R]]l�a�1�����Ǳ�~O�U�${qQ� Q�z�Bm�Vk��ql06��k>�o��Z�lx��w.^�{���X���U�;1֏�0w�ې��$��%�J��!�k�B|b�ޅ��MȪ�ȏsQ����5�����{G4��TM#�F����:4׍X����O���0׆�'�C�h:8U�����1.Ϣ2�E�j�
i��)�+W����p����Ѝ���zJj��/�w�	_D>?�f:ˠ�;�:��E�����ɋi騼9^:�8�rQ���s�*�D܉�&��=��}=M.�F������4K(�$�����Os�F��s_]O���E�aZ��pn��۝�e���dD�ZV�r:/�J|��K0;b+eכ�k�����Pbh��>������k;A��&
���
�}cɑF�O�3��Ɩ�Vsv��˶��%�E�`��-D�� �Y|�?��L�q����8���+0�ap���q����YZ]�9������,���/1�]O4H<�M���yw��������|2B0U�
�C_���'�4|�9u:
�X�cY�S����	�R�?��N4U�G1
0k�O�Tݣ>�C,�ߦ�%v�)����P��;e}�>C�{��&<��A�>����C�>�
�RׯZI��xp�ZU��)�;^,J�Cp���mRy������7l��x��1���j��������=/hl}�r:�f�B�;S��@|t���I����>X� �V7qA�:E�X����a�ƿ�M�U%�QV��]D*�����Grm��&Fb�݃ڕ�^��%��Z/函�(�|���� Y���_J�g��
�w��L2W]_������K����2�wc�v�6#�I�#X�V������2؎�nS����d�E�F"�+[֯�v���0�x/yaP�?����c��qC��2�K��l%V�ŧf�*�xv�8��U3��֯2B��W}��@"�Im�f�J��zݎ�Nb�N�K��Zhk����f��!�"��+���X�0���	G�ɦ���# 䳽ۅ�6(W%������Q�����GWM*[�E��{�ɉ���@�,R�
�e�I	�`�	r���Tzu���R�
j���㊷����R�~��� �9O�j�#Q7����=:�̘�vb�GD��p����Ϻ=$O�z��A����7W~����mpo}�ܛ��%�� t�V1�{�	��2d�|@X�E5��7����vh��ː�>RƩ��h��J�e)�ޏ�y�����i��`N}Ɖ�_��6m7�4�����<�A!��+a(k'�##�*ҽȼ��۶��0mcu0ޝ�4E�*���SlH{F����#|��\F@y��>x���r�K�}��ar���젙���/�g;]���̪��VBꟸ�����H[T���m����țt�*!��PE�&�W}__Zn �Y�4�xB��:��MS�<iN�_����-�����Vt�+��m/�kF�I��r{��ċ�e��u�;��U����{|����1�5$!M�đ�G<�9q�o�I��H!U�YN>[$��	fnc��������(q��xG��sge!��d����Bo��\��#�:�`�1x���(�����cd�FhV��ܫ-j����� dV[4��^�����#7ML�9���;�?�*kj��r;zj��%X�[��Y`��UL��5�S|��� ��8MU��}��Q����Ĕ�N�wC_I�`D*���Ͽ�h�4�Ч<¤��yy'���upB
��ʑG@�@�"�����\���3�;i��u�Ʊ�&vg��y�y������G%k�"�֣Y���M�s�$+�Qx�=������{q�͘`=:��<��ϪZ�X�;��1b'��w|_����~�|�������)/rR��|��w��@x~�f叻�h����<2q�m3��Y)�N>��)�-u�P[�YXW��kO2�|r̃.���lS<C2���MQ׿K[#�
��C�/�ԯGs�S\��ԷJ����)�9&�4��I�옪!�D�	��A�{��ͭ�GG�D��#�-e�էms��yـ}�	G�Wk]&J�q��7�Z�:�p&>u�ѭ.���0i!Z2{G�ؗg1�ȑ$4�������\���Ƨ��l�ѵ	������;;xA�+�t��i{HjϕPf^�w7�ɋZa��'�ҤϬ���*O\��!�&�P��+]l>"���m 1���d�3�>�g��h���ӌE�[�d�si]�+�����ك�����h���B�m�-�xJ/ŗg��Ӌxz�&����=�� ��[MBK��wda�#���<�W���l��*_N�z�JO�K�ӿ����"w���6�	�It�����+���Z�Q[�;�-��r��]����<] �j��y��q�2�p��ʥz-w�֟��9]wW���� 1Z����m�hc��8�:P5J�,	^<b�r�G1ՠ9��䉄�Y<3���V�eG�>T(�/-�ͯZ.IJ2���]��lV<]�t3���8�&w����%(�b��)o�nє���5f0�(��*������d��ڋþ���z$�m_DP㐤G�#.��ݼh��-�n�����3�t���[��o˾�f��oh��q��+Fv}݄��г�·
�q��@�}���q�$��D����/�-�����ª�ѝ�f��H�;�*�w��`���_\:ا�Uy����������@��P�^U��|0�*��+�8N������aB�+�e:��|��zn�����ĶrJ�~�sScP�ɧ���h��P�(Y���̥�*R���<�O�O`x=���������4� ~s9��1���+��g�Fv Տ2G.h�~?fi��o$��lu�C ���2+P�vȡ&ئ��T��*+��}�Ukz�yz�[�N�o�7�cd&K��&Thd�vj��#�ES�0�ݟ��R�و��'��V��2�;�ne���������7�9�§�|sf^;,��0����v�������j���-a�G�b8�8/S����ۚ�U������X�*�iH�&�/���:"�lmf1<��_��'�n��������a|����b����A<G�=9x�3�.�����1]p8�ꕤy�w���o��C@2%o�ׂC���/1?�6�-�k���8��������F�a�9
q.�t7���C��Ȱ�a�ȫN搿�k`���֏�Ԇ�dp,�yI%z�K6�g�v a�X��B�����J��ꪘs�ԄT���M��x˵Ҹ������;��3x������o�V�u��8 ����S�+�$iAY��g~���{%:}5�����$��s�Ǵ"���<���	QC,)첾��ԇ���5{g����݈�E�V�n�ٳ0�|�T^uN�Q�>��D?7�����)� }�D�e�8�*@�.tA���(��Տ3�,��wG"4jl:m�٫��D�7��<�ќ�Vc�w����W!ݏ�e���e������G���t�,���=n��Qߒ��R@��ó�F�h�O�#��Ϭ�����z���Gd���=јV��xM�P�;��V�$��cҫ
����.�k�;���$f-՞�~K���7(�j?��,��X(ϗ�|%�{����3B���������zL�#�Pt�\H�%�^i轨V��?PK   �cW�!ߔ�� @� /   images/f1137482-0179-4042-abd2-21e421d54476.png�Z�WT_����K���k(		Q�Q��g ����n�Pj�f��k��������p?�u�>�~����N��  �Uy�  ^�w�`�{2:� �*���*(0k��X�9~ |3�`k�PAN�	�p�Tp�޺ �L�q�`�=�%Q�	ɵT��\�����l�����lV�c�'���<���:��<o}��P�9�>�������� 
.M��e�O��@��b�/�3�B{�	�L�᱈�)��o�B���*��Qȧ��h��ql ���v�8T�N���4=@���c�/��V�\�U��??��&��c��A�6����He� ^��	z��Q���o�Q��Ű��ƪ��IDI���@��b�1i��6ٸ}���Co�}V��SCA7��߿�f� ٢�3���M���(�n��ۻ=�r$y&~l�e�Gp4��|p�J��N拋]��[��%���T��c���o�D�M�{}����N���I!�l����̢$�:���XT愈�w�@�ڑ�]6��-f�z�l���|`�Hy� 	k�Jѐ��e��?�ڕlo�u��g�)n�VqW���A	u2-��8��؟B=?� ɿ0�t�pR�b]��xi����d�I%7�X ��>��!��Y�D.4�^8��V^�.�~�U9o�qc�kr����
�� &�߿�;)t�O��$l�L�q� �j�'z|�eH0��^D���
!/.���	�e_.�4��jބ������te4F[��p���p�$6�8c��'��IB8����7Y}�~"�v��}�M�R�'b^�H���q�A�Y�I�=�Y̵�<�=�+��O�D��쵄c�K����|��Ĉy�,�z�J��
����QK�����b�{���I��8X�]�����r��a��M�Z-��$�1�yi�܍�$�;��S��?����=%"�Tұȯy��ԢT�1o�^QX�4���Ƥv�����M�4�Ys���f��h& Z	?���*���6�N�����zܪ���j���,�[�2���yn������2&6-�!QyN9Y}�E�Ee[�U�+r�(�7:���SU�5*�EH�ȘH��U^���}�f��cb|"���9��?῎��y�Z�qʑ�
��)��d�pQ�b���~��&�'_�F�^�/n��ˏ/�_���/R�ѵ���0�ë*T��T�M���������?A"_^�N��-�w�������Q�9�MZ^5�s �hk��ɻF�ƠƘ�`�dg��i����_W��������dM\M3��X��믧i訕i�b��^y�u�a�kbZA�N�/�l�q�>� ���OB3B�v"�yy��9��&����I�-�#�`��o.���m���"�$�����r~��n�D"���G���59���l��A��0{F�D�y�`�u�5��gD���2�:a>-!#��׷_�V"�b��xD�E�����iJ�]O����dV��K[me__.AaW�h�F_�Vŋ�g~ζ�y,�t����R���/�f�f
��ƣ���}	��i��g+\��tK�5ǧ����0��F+�+A����C����a�F���G�bZ���b�ލ�'�Gn���ކ��;WsK���R{�[���m3�L�YUY�x�"Z�ݥ�Ɨx��KW�NtO�N��r����2�\ts"B��V	�?����VtN�N/�����xΪ��3t�"k�
A� �U1n��@�n`7[wVpy�v��`�G��O�O�hɘ��X��x��sm^��)������#�G�K�S>�N�_:;�]ʰ�I��R�*��� "$�{���v^\-o����D���d�T���e�'o{~a�d�����P�?���*��ZO�W�q���f�ߚ�k����[���h��n&��ʆ_�j�0���e[�Sq��W ���L�O��������8��u�Ej
��/�o�~~�!�]���ط(�� J,_u�p�w�`��.��afh�j�N����c����[@����1ި�B���r��+��yk�%�z#�=+Ok�����4��nnW��>$G����5���f�a���ѻ���C>��N̀�쟓#?�*��U@��Ԧ�J8]�`6c~�<����}9�w��|=�R�b7��t�P~��D�5,��������{�2}1�wxwX��t�3�iu�c���V���]�ku�^��=�a�b!��6��}�i6}����ʾ�^�Sf����y����O���rZ�SNعE��n�	���ܫ\�B���d����l��8����f���8�h�֭hn�9>�9C?�����n"v.�8�|����x���W����>���A>�O&Bвw�W�F��9�-�jznq�Ư��ɭ��?�8V׌4��:���wY0ׯ��gc�K���/v�Np�:�ޜ��K{�H�a�u�AM�y/�2�h��u�_p�_
�:h,dU�܍﷐gMdi�;7�zv--W����<��=#v���}:��N�{8NI��zr�Q�a��ėL�?��A������K8����LWw�B��T���i����?G;�'��t8�~|��Ǉ0S5�'z�Tv��g]��~Z��X�@.L/X��w�v��6;���~�8�%sޗޟ�r̗�Cr����}Aew�Ȧk��e+++��$�)��D ��Z�$�2Od�p`�?b�2�����f�� n�љ_3A�\ �"r�4�ɜ�t�DD�s��7C���	�?r;�Ř��N/�%X��}2�= ���n��[  x�F�Qf�Ǐ����2RR�G�G��GnG����'Θ���(P=>������D�W���� ̡橪����c��?ދ�������/�$ �}�,�9&����]AN0��|��:���E}�oОu�ݝoҝ�-5�ͤ�gI4�<e��B\)�<^�Y�$D�f�n+��gE�n�o���\�h��,۸'�)*�V8}��N[����q�N�����bX ����R�Y�&�MW�,�����v.�˳���Iǩ�T��%�j57ϰ}z<��|��L0��*5©�\F�����0WCo��jf������((��܎�a�k��2Hb�%}�l�� ��$��a=��V&�O�Yk;�4?ՙtx�wxKt����-;~r��;������;���H�u<x�r��M�~�<c�l�"�ů�H��E�@wQ�E�	p��8e"�ƲtS.,Lk�t]I�vT/�1Ca����9��ڨ��#d�Lڦf'���f�(#����m���Ň�.�l���O��6���v�ח������k m���M��g��ƿk�Q�c��)��K�n�>���nR#�����_)�	4�0���T��{��ʹ��2!���'�m�I�����9��]�����y5���
Btb�&�������4Nj�%�������(�Tʗ���>Hev���[7��#�q���-ENci��d�r�3�1�%Dl's�P������\�g	����t��b�䧤2���	�ۇ=򓢹F�k�r�6�T���b�����#?x~/��9N�����'����v�������i�@Z~��v~h��/�����S���6"�1��0�$�c;n���{��E}�c�\�<�=v]��w�S��{d�eO�`���a"���](I|�U]t�Ng�R��rA�\y"�h'9�]=q�����e��F����x���fW�%��K���]<sy�����(��X#�����]�">��з	s��F��������?+����R�U<�3��C�4q�[�F@��)��.���viփ�Q��N��>yȊ*W�sX�q񬂈A���Z�(o�Q�ae������M����7��BQ��|}�Uzk	��¬{y@�����
CsOPZEr��z����	���l�[Y!��{X^@��t|�|z�r�xa}���T����ҟ�3>[!4J8���m ��ڝ��Gw
\�W�i�2v�H6�N{�&��z��Z3p�����X|U�]<�x�WSʄ~>��aĔ[bI*W�1꼀�ˀ�U��ɸ�ݗ�O���Ѹֱ�6�C>OaW���*/�V�!�#�0���ї	�y��
P�DXx�Hͧښ�y\��$	��y+�'5��b
'@	>�Cg��6���f�$��9[T^�ʋ\��z;N�W0�woa5�a&p'�����I����ጐ�AC<�Gtϧ�OUs�G�]j��7y8La-�O�����C������� ���>����%'�Q��#��hK-�h8�n����_�����^��2�8�6�;�����eZ�;.G��ܿ�M��3�?�"
�Y! ıi����~'#� ��''Ԏ��HN��J /�=�+�ݫlX�����m�ポK�Ž^�w�[��68q�2�J{�h�^���V#?i���\�	��׭��6k��k��`t5�-ړfQ�`QN�l*�R/�G񭴸�F����-�WT#�G�kM0#ĳ�9��)T ��
)�&�8:��nV��`�S�yBM�x_�Dz-�k4/�$4�(��4s�V�b.��Ĳ���6zK����=�-��ln���?�>��4��'Q̲�$�urx��춁�$���D��J/�2� �q�~C�k��7���4��-�z��Q�aBP��ݏǭ^Z��������F�yˍ��h:���v@�������1��E#iE_�x1_���°�=���0�[�@?����;�\>���'�@�))�Y��G&��*����-M�9�R`vk�>4+�N����z9p����x~�����pM~���$��\�		f�Iﰿ����o�h�n��G��hP��kP��<���8i�x8����`
n�����Jҳ>�d$�G�vX�&O�����'b��kˣ{�hx:	G��㣓�����6�,0���֑e>�>�t����{�h��]��䉍n��D�J�i�F0���t�]��Mq���(����"Z�*����6;gr�����sj�JJ;�QPX������8g���U31�џ��i[�����v�lz�,�<yb��)q��#PEVZ�,P�4[-�7����^o©?Q����+��KA���w�3^���x?l�E��@�|�a�3(���O-��(I7����*j�X7�8H��x%<F�o�A�V���y�]�����3F���6�(К�׽�u9����@����~�8��V�����W�dak���V���-���]$[O҈� ����W���R^Mg��v-|�h|�s�
ߓ�J��\d�S�y��)����f�*����m��g�ʨ�6o�������g7�yn�v;�g���1ȏX ���Ź\]�G���+d� ��)"��+�4åN&Fԩ;D��9i��Z��pz-�*���e��'���P�1����A��묌@%Z�n2x�@|�p��#F�ިu� �|J���Q}nͽ�S*�#�����G���j��c�'���]c���.iC�<W9�]�9M��b���z��·�ԩ�]��ٽ������^C�w՚�vM�8:�d��ae���|�OA͒H��S�ң$�~.٣���C_r��̵{� e=�?P<����d"VD�{�`h��W�
��d��O��/�<��DB��?p�Q��
+�hM(�q7���Ґ�Z}ǔ{�����A7	KC��N��oB����@z^@���6@����:��T~dIu������G��ħ�8�r!3���}k�1��Eڶ|n�I!���"�����X��lHy8N��`'&�%W$+ ��{���jCy�?��#���y���Q@pF,ܯ���o\�zΞ�0S�nj���5�}���"M=p��Da�y��0R�=�g�p�|��:�fm�zp#V��!��P���8��릜��6�� �"е�	��`���W)h�y�|���m�<�^�+v'�~Po�_�%M�&�DU�$�-��ޒ9�����ŷ�$��V��ƚb���1Swh[�2l���Eģ�T�>SՊ�~��~�ꁮH`�Qج�?u�p���}���*��QYH�T�&�I�\����� �i-�/7d�r��c�	��^׹s�c���H�g����B�NE���н`sۆ5�1�&(�ms�g�4F~�����q�ٳ�n�E|�	�v�4*�ש��_�y|��ҩ.� �
��l%5�_���*�m��~��H�����o���~|�Ϋi����A�Q5t����^cٓ�L��!�4��9�y�����x�e6z��;��u�e,��U^E���ߎ֘I�Z��< {K1p�� 	w��<�Qu���b-�h��zN�.�[��ŸV���s��i�_��~K+W���.�A҄�M��y%D����E�%�~-a�y�C�R��M��U���	��/���b �Pz�����5�	����vˆϐ���
�x�����a��������{�n�[=bj�� ��@���<���E�̞� ���z���f}|�z&�mTt]����j�������z��v2��[�TnZᨶ�Bz��;{���Rx��'���'k�?,�aQ>Ob���H��Y�Q�5�=���Q�U���d��t��Ƙ��rꄀ�%�I�����L�[b�JA�g^>W.�o�_<R�G
>ۗaq�����z�_BezD����Wt�dy����M�3 ��y-�&rGOu��>�����f/���"�z�A�Rg�������/�3���׽��2��މ&*�p#���k�4&!M�!�8{�����C	?����)������~)�/{�X��Z���K�Zx�I�$���ǪX`Z�����G�9|e,���1�����j��ޜ�Ј/�?c/��O�O�h1�v����J��淮W�1O�����sN$m�㡑2�2�6������7t��E�ޤ����9�}-M�&	%� .;{�{T)��x�W]�����	^PrVj�}o�(Y�PI����7G�B�թ@Ƙ2���D��|h�\������,?v�F���"n�qk�7?oZ��5�[U:�����&���ä�N����öǗU�2�k �d�z������N-k�Lq�ة7_GX[D��&:YS��;pb���'��V�6�±H�j����Ն�!:��5���P�Qݰ��Iۮ�j�����T=|�(��X��wl�� Eu�64�����<$��qֿ�*�����s��|�]����u,�u�ezQ��	B�`N|��l�(E	k�ޯ�U��~m��zƓH(��B�uس?z&�sp;��{�ũz&TM{`��~#�κi��g�W^�V�\,��z/}���3�2��u��92�Ro���{���pFS�wg.+2����x��-�{���/I�g��u�W���[	����� ��a�%��|�M�_���-��5%��<�o�O�a�K@͢<�āpR���[b�W|�?�r��x��=E�ʂ�Fe��L�(��T���ѝ�_;�;�;�������O���e��:x�K*��jrl����đ���	@��vV�)�u��Rͣ�!��s����-X-��	�>`�]I'�!i�5&X�8�Us�P�-��YJ�NX��i���U�H=u���Ԧ,�YTC��^�)��I�kZ*������J������f�e�qv����;C�}�&��H'���� ����>����<h�>��,�6�y�����1WTփ^���@�x�{�h�{�]�b����d�xHj+��>��2(��Z���f�[x�M��#,T'�#1?���Ww.HK��I6�UG�Ӈ4և�ݜ�;���ܥT��M3�	7��h���]|�ki��Dk�q�wj
���d�0�܉vjB#&jW �i෇�I<�$q��*kh�%��*�d��]����~q�m�:������&.%}؎Tz��#[��4a� 9�Y�	)��Ն���E��$����{���=M��l845��T��~_�5>���sk�[�S������L�=��$��j�������x���0f-/�����R�:8��<�h�Pt��(�f����}���|�볖��>(��=�Q�%mΜ2h1N�=~�^�$Eݍ�ώ�3\��q�)H�C]��u[}d;0)í>F�M;������N;Ñ��tTJ�T���ʈ��69�v�|/��ӟţ���j�)�Eg���G�0�{�7O�/�H �����Yy%�t���S��Ċ7��MZB:�V���B�1�ɻ&�P�
���?1=gA
�q���:W�b{H*O__��Q�?�5���;�!z-/?#-�i��J;@s�bh;�h�[�vH
�0�� n-�S�ڶ�����[y���S�.q��Ij9���X�7��!���a�~ct|�6���Q�C8��L�[��tVp�L�ܤ]lQ����V�
b�Y�*�p}���"�K���x���fjaۙ	@N�����[�H���~Y��U]{t
�U>�h(�&���뼅�z����hw1B	��+Ơ �O��/��o�&��^��2S��
�#p��򌼭���>vi���w�$� S�tD{��>;�1�l�T�Q����SI��
��N6;�
�������FX�Z3އφ��'\.XsƬ(ܯ��w�"���k�����J�t{	�1�D Q��%�a�,�E/�/�Ze� �5#����_�n���2�?�D�m�5jl��"fA��.W.� �}�^�q�,�� `�7���e���������8�C|1��Fee����`A�7b�ڐڌ�L�����nf�MAOή�t�2����e-會��ZJ� JٗZL��x,��OI/�!2G&��V!���^�3�˳+�__�:w�t��J)��㴙��q�@kb�׫Z`巳:�<Jߒ��Z�%h]��N!;�ڇؽ�6�W4��x�bP���.d^��l�f@������`�^%:��j�q	�Ǻ��nGzF����!�}0\G݈Vz~s�^�v85���$�<�ӳ%�\>2�Q��<�u��n����g�Ng�K��d�1��2��L�����c�Sl �_�,|�zp�"�C��'�*���АUe� 
ۿ�Xg�&C�.Ҟ��Ve��Bf�L�o��(�����t��P�xl	�B���?]#F2���	)���Z�;�s���zMO6xr�6�VP���ǌ�R<F�����r >b�:���敓oU��\3�5A�[y��D�R�~�&:LѰ�F�<��x8�a��5	W��\?_�+(L]�"9 ��p��m_������C� w���M� �2��ЯXtp�`Q�g�3�����^9n�Cë��8�Ko
<��v����S�bm|uμvح�ICI੼Z胑/�:PϷ
تuu�K�h�͈я{�@��_�,�۱f��s���)�=O�t�{�h(�}�.� ôV��(_�3�	�l��o�= G���{3�^h	����έ�����/@�Fd�~�`0�ٕd��B�HI\W����l_���e����V�	�I/8~��J�����F�%@�5Ԛ�dζ��Y���`��e���Ԁ�F�@ÁƤԄ����"$���4�t����r�h�rBx�S�L�}ݝ�sJ�m2T ���&�|߯�7ϟ۟aY:�!�����<��ޖ^�:��9tI�~�q�����(����"�y<�2�-۸��ߠ'#����o47e�@0�y3��K�6�a��6wH��vR�rz�1>L2y5Mi��6g�p������*Zx76o����q�O`�Fo[�6���H��,f�,t�}3�;Í�$�}�Բ�i�Ľ2��p�G>9�6(��n>9
DҖ	;��Lr)>̾g=�=��"]�����R�������1Tlr�o<s�>v�n�t�H�1`�	�ˣt��`���O�N{�/�}�L�pC|�3v-ߕ���� {1��]����UQxc����R]�\�='���~%Q;:c�2���2)�?9��@G�%�9��}�8o2ݳ�j���`�S�Uڛ��x�%t����Ώ]���k��2}$��<y>wd:܌8�@�]��'�I�]�s4�@�J��ݓƵ��]Hz�9�vP�}#��V-��o�X�%�� ���.�c6�p��p�טwK����@W8N�;������V}UN�d�9 .�s���D×���
nQ�E.�/�cN?c
ʂ>��/���s�X���4��Y9�4�ʭ
�T���O_���ۉ��o�_���r�M}2M�)E*�w!���#z�����j
T�< ��\��	cFc��ь�R���H9s4���@/:�VL_�d�bl<�G����l]-E%��aQf��Ʌ���T�ٖ�L���Y3�O/�10A�M��/^[��ƈ�˸a����;0'���z)�	)U�u��g�W����k
����d���[�Q�8:�(�vx���"W6L8��M|�$��e����v�NS��R~ ��`�X�@���JT=�>�&�f�Пun�~�5`���ƅg����j�e�R���:�~C�mG��P������K�Pp�9����9�r\���f�m��/'O��`��ª��w�|�u�6�8�;Y7���S�מCL�Kw���,�4�K����m2�3#���&I�J�D0�o]4��[ƽ���Ǭ-k�v_��A�V���J'���mB�N���oY�3T�ݜ���J���|���~g�Su�/l�aW0�o����H���dmn��rٿ����9�儫�ը`�����ԭ��,;��آ�����:�9�����!0&}6��FtN:2pq��<�����^�� ��v��s�F|�V#��Hq_�v��c����i��]��L�Ըi��a�X �\�c�,#"��Ʋ��ɏ�Bo�5��v>,�ᛤ�`���~M���P�Μ?�t��\��R!����v��a:��b�F������iH���fw�Ğ�ez�Hz�*#cAp\mj���l��!��;ۡ���ad������xgU��S�9�2�
��ޗ[��K	ým�@�H�|�Z��O#��z�E�����w!1˭��aW6F�x�]XFt�L��g�l��o0��U2y/�0,��
���,!풎C�u�x������u*~�$���PjY�&��:���mt�����Ű	��q���L'�
�1J�N�&�Լw� �L,�7�m�hA�N��B[�Y�ɳ�t7[�ۮT)���^�j��r���9w��bt5q�FH<��=�*&����ȣ0�1.S[��dBsy����r)���|�nq�j>lvJ�!�[H)��O?�H��ė�N���\��Me�O�b�%Ϻ�5Tï��7����U^1KF���'����0�;p'W.p� ���3Ά��߬��b�Q�x��;)_����(���8�X�oj ��+���h��dd��i�^�l��*0[�8�FTɄ/ĊkԋhM
g���>��,�e�3���Z��3�x�?|����?���"^a��!r{���B����0w?���CQe�Ǌ�B�6����!>��t�1�����+^L�\r�&)��bp�򏲴����;�}�L�*wP۲}œE���Cҁ��}y�l�~jw�{�A�W�d����ԀSE�
$���l<�"��i� �f��K%�HҐ]��x��o9�]�pTl7�G��^-X�#��
! *!��(����K��''(1�{�/5��x��M4�WH����|Ьz�ϰ}�;.��M0��o�Ϝ7m�Pع��ΰ��=;3��}��=�3JZ�͚0��%�����
za[H[��[օk2�#�Ov�x^��*�\�{�`��N�@㹄���C��כK�Þ��4>�E��o��8��{o�Ժ�ņ�ɪ��G��6�{9.����|��DB��x�� �|N=��	���[`�Cҷ6c�h�F��1f��q�����]�����9\k�l�ꚝ�&��4N�?c����P@�\��,�>ш�d�h�u��6K(��°N�P<��}�q�a":���n<�L��-mw"
�+ys�����Cڨ�Rs���}Ήs����h�,�*�ݽ��z�����r���A��?��xbݑ=w��Gq�Ü�;>Ŷ�����o�8x��Rn�G[y���,V-L�A���.�mM.F��@Y�����sio� ����[1�j-���m�
���:��sCx3�a ���E�Y��~�ߒ�Ǩ������y��Mb�̚�)�h�FA���sr��r��uqXf��"ߩ{�� ��ߤ #�W�&��(�,�����jѤi9�������OP�Zr:o��<�Xe�b�'�
^.��mkb�2&,� j�~S�`F�a3\EDz�@y'^�A�V,�ؓ�S헾�8R:X��y[�.ǖ:)y�2����o�q����$˷O���OAӽ�n�VY�#���Կ^��(��t�z4쯮3�t���}'�&3��2�m����a�\�K��Nkl�9�(��ӌ>�ǝ�qz�Z*Ӳ�f��([ž03`�pZ��>�S[�"I�2!+�����U�g˜ȈV=�RK�/pv�3�9����	?���H�BO0��_'g�|�A�E)��k��ě��UfǪ��ŉ�6đ����lF�����?�N5����q��H�F&lߙ��Oj,�q��|:�iv��&®�� t�}6?><��8*�:d�s-�:�ў�r���|ٱ����C���Ru��I�NpB{Ȁ�qW�~����Ϗ��M�>��_�U���aݟ��3ؖh�SX���g��_������I�#4ϐTa}`5��%�V�������y�S�W� ���}�b���(�)bX�I�!�׃��ٚ|-��0�Ȼ����%~{E�J�r����c��''������ vV�rd��}&��^���c��ga�����B��s�X���9tm�����7��O�UG�[i����}�M"vud�3������v���Oz��v+$��&
���ȿ [ǂy1-����Xb,��_�[i�p��o���T,����1�����ua��)�g�V�i����K\�>��^AB�S��>*��A�ƃW�y�N,U�
�1�����ug%�`U|}������� WI�[VR~I}e�E-I{�c���
�Zc!�!��HӟJ���e�a��{�I�σ�~�p ��KCo$���wޙl&����N���`p�N�ǲ�?%�����zD����rg��.�� ޜM
|��dנN�<��l�1����x���'�H{� ��9L�m��5��~���x�V���p�rQ��gc�;y�c:���H
'
�s���1E!�����%Vc�m|+c�;v�����T\G�h�?A33�\�V ��+;���w�	�n���˙y|8y�"A�|���*	[=.�&Yn���G�pM��20u1�:�V�B���T�{��xn��h,'3Տ���Rw�Ĵ���!ْ������%����2*��p9,0�k���N�y����f�5hޯP�^9�D&oXZc�t��o�O����G{u�����Ю ��0t�Ě{N�/A��f"�Igeg��"X��p��x���=�Ñ[�[��<� ���>k�qid�ڑ����g����}�������4�5g�c}�������
��Ǌ�S�4�$�؃�r[HyfEB�B8Oi5����s�M:0��EƠsy9{&��!{4����kS������G��s�Xїz�D�=o	�,�n�l|���Q�o N��͔֘]� B��e���N�~\4;��C���b!�z�,�����|�~�&��?��҉���=��yh�zb������{@��
-��2�����	8�)�*��(	,ӢK0���zJ�v�F:�Z ��p�([��i�{���	U�V��.�p�-3:�w���J^�e�#^��B�̡n��~�6~�.^ˡX(��9�K��~m����mT`v�C��%R0�?{P�E�op{�s;��$���=1|0C[1G������e�Ʒ�1��<�;�`�v�=��7O6ˍ� .�瀈l�Adq򔲆�έ7�+�̒�T�Ѐ�>}�
�][` ���5&i���������,��Ǽ���=I��n��cniv�O��� �:$��(��VAL��c�r���r(�F��ʤ��r�?��2Uf)s�������&(�3�T�Tד�����,��U�X�f�V�@��K���(��k E�,���_p���n&s]1$�(��C���͓��k�������6]aM/X�V�����JN=Z�� &Ạ!����;c�C� ��І8F�M�tl!)ZȪ+��淛�u^W��D��(��)����N�+/ �93�I[ea~?������(]��!J=}%䝣!5\C�����t�˯��f89�o�,#�ӣ���ƙ�d�CZ���,-�'Xo)K����/(�L%@�aݗ#��:[S5u^�sN�K�q�[K8�fߣ�Ѷ�-5���X�4�#j₀}��!��]L��k��'�t���
&�4�p�f��e��?aLhb�bp�����;W��і\�B�u����@��1P�P��ř@
Z<��4K:�p���v��Y�rj�!����:��_�[����6m��������[�+6�&�w_}r�ک<4�S��$������r�t"�"=�*����%���!��M&m>&c1b]�X��|��O��j�9��ME=���M�b���NY卛�ٝ!�?N������%E�"��U&��K��\>Л=E
/_^�^�G|L�w�IaY�iC�N��{��ō�*q�)*�;��V�l�@�2/q�b/]�������P��K_���H�>�ׇ
�3b���f��4�,�j6p|��k����h>�)�����5.��/G��D�_��n�	B�AN@�8/1��/�ܣ1�w�v?QJ��!I����]8/���=�|V���v��l��#��Fe�:p�d�f����KWj�o
��zOX�v@�1�<��VX�JG��P��T(����m�J����e%���g��x���jzE�x����@1΅�^�&Y��a�u6+�-�_�U;A�O��ͼ�<���anlcF^���j��'~& ��L�F�Jp��u��ʻ�%|�Y�P�R֞�5�c�ܶ�#�7]��Q:�w��o���KC�q@�q����B�TYF��q��K�)x����s U�Ǝ|��X��*f�F0`��kb,����05
P����K/�� 4)�ڹ��G���*;��\s�a7?�`�m[��I%�4������g��J7f�\]�yS?j^~�����}Y�tJyv���z�%z5�ނ���Qw� �'�TP�Y_MN�f���^KN���{���U�w�h`��"N1!�����߽��
=���N�T/�l:L��4o���=x����o4y��į#(�`'�R��0���ζ�Q)��if�C`�+,�AL�mD �<��K������+���}}y%cD-�H�V��-s����X[L֘���<�9r�T�Y]4�?k������HQ�Rk4�ڵl�S��?X)o\�_&x�ɹY=�#_!w���j;��]��܁L|�� ���B�כ����*��A<���$��cv|v�#��Sr�:���2v�aѽЪq�5jb�ʦ+��y���i�7�9_�[�/��#I%�ԋ=h��B[d�����F2
V�g���n!�q�<=����Q3�%��'��wR}JF̶�����Ytr�r^�y�țܟ�	'�!-���Qd����}fq�H��6��~�)"`!>��d�B�'	��vwK��f|��#��u��� �iͩ���غ���/ݖ�A���r�1<P�KS>�A[v���O����)���W��j
��������V�o-��[��uF����,���@rc�Wz�BW��CAl"�-/@�w�����{�D�X��r<�����CD%��Y̰3{���a!��Ow��{�3K���S�4��Wnh�2y.4�Sƭrh�U���U���
�K�w� #�[��	&�M�o���P�=1�b2���8��$Grt	=��n��'���+,��k�HcM��6B��k; ���7;яף	��
-���Þ���xXAVz������@B���>�Qa�������2x��2la��JpY���Y�u��mر���	%�8����G�d.��a��d��~�?���H�D51u�}m�'N�����By�'O�T�6��@{���j�#�������n�o�xg5��\�KzE+D,�������o�$����~׳�b޿M��=̅gH�����s�f�}(��:�	�K�;=�Q�^^~���֣�Vz�7ٚ�B��:=��!4v���@����� ����.�K���(UQ�wac�Tʒ��b&2����.���C��C�(&��12������V.����#w�3稙�!c^�V�'b��F������f�d�Z�)�q�O��~D-Ӛ�+�q�W�󪂆tO4�96E�����;�������0 zt��u��ہz6[���j��y�8�n���F��������>%��6�/��
��Bﯡ�g^�1^�xO�j1zM��M�tԛ����d�L� O]�J���[�d�-���{��5Ж���蘿s�-�Y rP���QH2���VJ���*ש����" ��7��ù]����}����~�k랿qN��`K���Zj	����^6��<�y����@]��v۝��\��sK�t}�P z�б�Z�_� ����ua(�8~���n6��w�/���[��>�Ќ�r������6��|r�ړ �VT��(@�i[�!hS�ڶv-F��ZC��c�o�@@��Vs�j��Kߞ���@	�wI�#���G�I��\ðl,���\f�Yk��(��6��wjFn�G�Zm�i�x�\��������s�8��q�� ��q*�鼧1NS�ݯ�H������y/D��q]8f���k�OsȮ��f5������n��-����kc����4�'�ם5_�}��D��lW���:���;�>o˼���S�%[走b-ނ��1wťh.ȧ�5�,pҖ3�oS��s�[�Qg��~���K��ߘTy�.���E��>�rM@���B@�P�kI�yZ���]������1W��k����͇b6bh��@��f�+��?j�{�'l��#���=2hР�0�j�َl�^��nX�F+Z�X���Otsq�����:a!�Z���N�{N��;�����O��1vo�m��#�1�A��.\E�s.�а�^��7��|c�S��p�K${�꣹�y"a�A�1�Ѧ��Lؚ����w�}r����y��²�6>�7��S����3��?Q�n"ib��ls�1+r��O�|�J���9�9���Z�&�u���U��e��*Ƌ��Y�?I�翷�v�ˉ�Oeb���V��W�k�N�yջ뮻� G�h��VӐ�Hv�Y�v-fi����~3#��f��d%���:x��_P e�A�Y#���l"u��η��ڋ�(�����/���7~?��O1���v�Щ5[��d3�e���(��>72|]�&��u����Vn��`��[����J+�A�#�z|���4��D/O �'b>-j��ħ�Ak �v4��9����' \��j����5����ޚw������8bZ�k �:� ��n���v�D��Ӽ����>-y���$��՟�����P�:��%�ϼ�[m��ʄH�U�v�i���{;�ꚳ��Q���;��=_�"�K *4��Ze����������~��� ��uQ�,u`�H�>�L�g�y�5>�-1k��mk�@������������ʥ5ټ�b2Q��Lڌ������ۼ���G�c��5�A��A_���D*m|%0���!V�z@�+qK¨7�'>���-1t'�^t�[��>��&�yunԺ-��R�}����6&y��2��|��ǈ�/z�
�I=��-��6 ]g�K 4��ehى9�z6��^�%��e�}��Oc`뎀�m2+��6T]�MaM>V 4H������@��,����3C��.`�h/�K�30�x4��,_����U����+vew]�k�ge�zy֭�?�b�Aݮ�Pg�Q�"{����9�fg��s��	Ћwl*�g�u!e�hI[����	�e\�����&��Y1^Ք��V Ny�Lk�u����[���䨅Fӡ5	11�XC�YÏXLJ��޺�%h闪�=��q��/P�ulE	pח9�01� B��y�6ֈr_uY0�c�D �0M���um���ҿB���1y���{�t-j��}��<�l�6�x���
��(s��M���e�
\�6��ct?�\�jԚ֠ES�g,1@��6�+p�B��ڎ�\u�������h���h�H{��&�(T��s������D�_�uԃ5Y& H0�`�v���w4��`>��~���.��
�SZ�i�s���@9���1�bM{��n�W�|Hm���ݫ��:֛���ˬ�Z�b>6�ۯ�P�[@��[9
��f*bf:�ҍA^f�1H�Z�����\l��P���`D]��+U�>?3��
+��6iF*J\L�m1{.�{L��f�6=1��&p�$��}�Qô��l��-
?q���������f�Gc�p�+��Uq�O}@��Pg�J�[�����3���Z�M�Y4���4����噼M{�����u��г��L��զS���w��=����kv	X�t?���j�z��ѽ����~� ����� KPF������|��

��½6�.Ԇ����^o�*��Z`G��&G����AU̕�f�Q z�Ѻ��t�M7-���d k( �đ��d�.��a���^3?o�*s�L����5xu�M��l�62gk֮c�]k ��dm\}��g��ߟ ��䭿Uѝ� �z�E�-�o|�`�3��޵}/��c
b���}���;"�Q�g����?� ��Uu�_���Z�8�5m^��ILAK��E鄀���a��yӑqk(ЉZ��fs���B��P��ݠ����0�_sL��2)�Vt8�G-\e���������V���9��LC�m��g�xJ(�i˚L�?�Ή�W��2���ZS?u�k�km����v����U�A�l�ZP��
�NW�X�������\H�'���u����e)��/���0�:����bb� l.�oR�+�H�k�+ILJ��`bԶΌ��f3fԮ�i�b06�:h)���~:G��Q�*Z��q�t���T��Ж�h��l�����+��gli�)
�O��T�!�h����� �8�ׯ9���Z�Ӏ�ۘ����P��zTB�6v�;��7�o���[7Ʃ�5ר�:N ���g��5G����D��������E�ڋ�w��y$��-����Y�砺�>�`F��c�w%6�GZHӖ��eZ��V�L���cZ�r8�im��ł�碭J��[ ��"P7��j!��?���)���Q:g%L���\R �\��.G��Ni�!���Җ��ʿ&P��QA�C�a�9���4�$Ř���TG��Auژ5T3+kK6��	;'\��Aq���:�#c��ԁ>���O?A�-�= }��0e6@�yx	|��U.��M��v?�o�=�#�ͼ�_�Sо3���~�(S�� /��0��"�KB��|}�օ���7 ��5߾����"��yDm|f���i�'�&5���EU�S��i���*�M�\9�ۚ~��>q��2���A�ڨ˸�Ǉ܄qj�x�
��!
�k���BbpZs@F`5Mb<��@] -ߺ�d?�h)�Y
�^z���g�}t_�Y��~s�-bѯ�1�`i��)M]���(9�Ԃ����H�<e�w����α/6^8?�'�<4�h�����m�{cJ^P�E`%u�Ya�[LC�� ^�&q���s{53kW�X�8�y��9�� M�6:���*go�|�4y#%+?�g	�D����&���0ꅢ6�~YP1s5�����b!�ϣ�x�g�C��s~
3�30a"��3G�ժ{J��xG@�/�34֥���ZǨ���ǣALc(�د�s��ŀ���x���G�H�f���>��� �w�����x~���r~��y���m�y�	ܧ����� ����Y��Uɯ�,<cK��������/ 8p_��Л���NǴ����T��m��n�-Wi즏�K�B����/�Z�z�yjM�B��(pڪa����Z��!P��|�v#9�E��jr�#ޢZ�>{��S�=���	�瞆E��h���B=�a�=��%��_h��~3s28h�L�29�x�b�O�`7C2����GV�ޭM��fzk �5�o��&�6 �V*r}��Os��F�E�o|q��-�,���{s��7M�67�N�@�������_;��}�ﯣ�=x?I����T8���'~��cdJ�?|��@�E/ƻ��%�ڶ5k�y}4�T, �l ���ڸ�G4�-��{,s`4sasG��}F����3��d��dΛ0M�*���0SO���RL�	B��X�&���Mߞ7���ܱ cAGG=���:���k����p�e�}�ɂ�-l�g�R�Ċyq�Z>�+��=���mv��Z�2�K�1�=��j��ޫ�y��?{H�>{�*ʳ1�w&5��hZ�Ø;��Q1 ��^Z�q1[3����۟&��jo�q�p4'�lM�fb"����561��TlڇA˴�:}��m����u�l���n�&� �+�n�T�R S1�I/a�����g�}Լ�%�z}�9~���7 ��1�>��U�J��HA��� ����!zQL���q\=��S����\�-3��񏮖�p�}��T�z�ø�d�|�\| y	��
����4	at2@���_�m�.����W%�`+��`�L�zY൰jP�|��N~�"����Ն ]�<��eZ��6���Wľt}w|��̾|�+4w]3B�:k$�P{j'�@��IA���jv;<���mU�8�_yH�^y��������v8A5[#ݷ��
���m��5sk�:*mF�C���Wg����ΉG�Wn�\��^���to���g�unA���<@��䐿5�ҥ��Orq4���<�G�Z ����C[����(�3Ӵ��ZK�5ꙿ�� �<mw��S�d��R�`��Uw�9�Լn<w��<jwQ/q�)Z/�ϻ<�[B�j<��-sr�4��-4��ݏ�����Q���~�d���P�=@��T�g�d!��� i!�z^j�X��]� Ĭ@�֒^nC�M�B��-����c�5r��%d#g� �\���XŎ8���/�Ɩn:GH�>Gd+����{P��x@mS���NYqZ�����s��Ĵef�)���fF?�����1��\&�`_�}�6e�=�Z.D|���ή�G>b��6�il��R�z�^X���m1�1uV۹�1J�-�fm�An6�����I]��ss���}��u|�w0`@�~��+:�V4�>� ���*�_�0s�+s��d�M�f�Q���&��m�@�T��	`L��5s�s���ǡ�;h�8���W�rfFo�N�1�ĭ�.sR����w���9>Z@��oi}@3�_Z�L[�Lw�� ]����\e��-L�]�u�1��V��z��j��ؑαk�kk����y��s/�W�H�^����cb�E ܉���0�jH@.��s̵���������Mn;1$k�Q��F��fDk�fr31��2�j��o:m��o#��u)��G6�t��3#&º���4�@��@�6jS}P����Y+r���f�z3��!�%�zs����!�}$�cK"��4D��ixY7l�d-c�8��43 ��,�k=^���],��s��W��*q� �	�����ʜ2��о+��=ǋ�/DXj�/ɼܗ��"멻��1>�sΖ���[G��IW��Z��v[�� 6�4X�T;2ۻ`Na��赪5l������T:����y����=nf���^{�o*�|��*�@�*"lU6�/���_,�X̍Ĝ�⥣�j��=�ix�t�赐]��LÚ���E-���̿0z=��2 �P�jԖ�Q�hs��ɸ�f��o�u�]?����KU_�|U�-	�l�>:������>虬��q"y���-��0��G��GX
�U��Uf�����<��l'��J�¤�E����(��Ϙ�e�]���vA�2I&t����PL��Ac(�2 /	KFe�����r�� ��
Jy��-_1F#�ي��Q4;�Z��Z��VV���ssR6nޅNcc��py6�k��$@�\��^u��\'��Ɠvw�{�q��͸V�ܨ�6�����w�yg����4�ua�P��\0FRR��L�b$6A[�7C1�G߶��P���V[�:l³�`_�@Q�Y�� j�$~�>�O_���h�`�V��?��j��K��*0�-�E�g�N��]Gk�1H�AJ6=�2�s}-���3~B�^@+�����5f���u
!�-���|3r�W���֖Ѳ0�@�i߷���8Q�n��q�����F2����@˓�)��q��<Sz��3y2�c<6UʟA݂��\�s��M 	O+��r-�G-�8��۴v5v�ʥ��]�S�4/�T���@O���=�Z��F'_:���vծ�S�'L�o�^w�s�=_�'k~��%4�w�q���4�z o]-N�����5��+Pv�y��cq>�� �� �ĕ����l�]�o�� aA��1�o��)=
p^���J*ڏ�`j�ooa��	����țX� Kx1S�afia����\�C[��(����|���%aR�ؓ�+c�@��Z��L�0e�F�9J_����haΚ�i�l�!��ti����3�� ��h�c����~�%��*��Y� �a�cl��:VW�е
��q&^C:j�G��=�W�R�⹚�^�
����5 ���ܖ��2�/^kJkS���Y��MSv/��HIpv���T��G2�Wꬩ���W.=��5�j�1��J��0���`[[uZ����u�[u����^9�g�OP�Lq(�E�>>/p��Ao�`X@S��-��U���0�����S뮻n�)^0�fh	����6����@�hh���h]3�����< >�F/��n�|�<�m_�J���fy��:������jk[L�6�Z;�1�om��V#�5��W�0Zk׷����$��a
����K0˂>U6�K�a��"��e����wT�E�b��l��cbw�Uc"_:u2��gTT�p��k\�Vk�n�Ql^W;��S����D�����J1D?�c���Ćc��n��[n�e!��� h�e��B�Bs����i�اn0�]ڷ�����),�Q0�v�i�����;B�L�̖�#sq;�CS��o ����w�a�O�#3EM���ȇ\[p�Eaxu�T,�X�6��"�h�r����\���|��O�U^�&�F)~�&]p;,
���4`�#�8�͂��![[-b`��_��Ӕ|�F��w񇿀~`�L��u������.b~�@��-0�異=u	�G�[Vg-<�E�qu�F�a�,��<U���S�v�ѹ偺�룫Js@�.M_��t]��;�V<���l��Λo��;5N�ԁr)� ��'��7߼0p�x� �u����_�Y�og����Q�?��F�A8�y?9bĈuH�9��ڈYX;�Z�M����S����0�z]B��7��'�ͣy��^!e=�څ6�(h�e�r�Qts4�5M_���ȳ���A<ñ:|@���|�˺G]��]� Ȫ?���V̑�6n�K�}�&����W�8֋�Goa�� ����X.J�\m)�'c� P_��h�iKS�v9�$���O,��\go�Ubk��+�]½4z��k�]�Κz4���X7@�w�ՔW��Q��S�p]LۑX�u��¸��}L�^ģ{�7��g~&�amYm-@-X�9XF� ]��)\��
p�I�*`�Y�� v/A.��{�Y�;&�-Y��~��}���`��>k�N}��:د��]��^��|]����	l�3m@@�B���C����bV�t?�,��_G�s�X��&�&n_j��F��a��Z�G��l�|���kTzF�ƣ�#�Tc��ͦQ�-�L��뫸An��o�8朢��pb���!.�D�5��Չ[����ZW.:�ul���kF���ʏ�
pZ�2�GM���.>��ũM݋�l�	ԝ��]�Bs��,];����W!�R�sH��sH���3�"��s��0��b� ��5si�s�tU_s��;H�ﯿ��÷�z�0.~��W���
�`]��k�9ߚ���A����r�[n�&���L�������Ql��aC�����}�sk2q��&�k���}~���� �Ƕ�f�/�zl*�} �%f��tۍ8�����B_�Vf!�fM���a͜M�\8R��H���;��݅&�V߾}G#�}e�ʢs1�C@�@,/�̸��FN'��K+�5�S�q�읱�8��h��b�6�c� ]��k��K�&g+��?��:� 9����Y�W�T7�_��O���0�B�ـ�;H􋠙��润$x����\8����>n-j�����0��Xb�k�ʯEʞt�u��I��� ����ڼ��ǝ�f�ӝ��s�����@����C��W�S����쨨�ma6�Gf��o��`��8K��i�r��p���_�Y�M�����M:R�m4ٍr�K9Z�Z�M�v��;����~V�'��m�?����>��rM�=�����Ӗ�5��{�^X��I���z3�]��E�<��B���	]¹�:CZxs0�ֺ�t�]'�]��bV�~������Q:��zUJ�3[�_ra�J3��׿���$g�u9H�^d����h�g !�a���o�����n3���������t�%��y��g�z��^{�/�����c���;��_�h���N�>n�	��\a��=�C�-$#5�B`X��/h�K�M���Yt?�u� � .�AL�`�?�L�p����&��JS���8��h�+滢�Ĳ�Q��|��q�'n��T�TvP���A���>��6ANw�i=AP�(�ɜ^Dk�B@ݨ	,��V��\��Z�][��[`����<��t�S�4��7�NoR\���1o_�J�ӥ���L��=,�;��sn$�m?���E4��+������lS ��h�gܲ�d����\\�MM��Z���x��rMz�wȵ�����6��ˣ�>z��O?�P e���#���� puЎ�l�`��R]�V�0����d+�x��Ba�]	B?[�h_��;J]Ϫ��~z��ϫ�M�o"�<د_��t��]�J�84�D`��XEv��/	�[�?.Z�������q�������|ocb}!�N�|�Вɭ��ER� �_��ɿ�n�ij�YsBk!��W�k}�*��.['Z�zY�vڛ�Z���:�CҲ��k��B�Վ�u��=�u?xG��H[u>� +�[��w����S�Oz�'>�AT�;�|-R->I�.���PZ�޺1��Θ��r-��l���C@���N;�i��ۢ�����,�1�]ѱN�������\���-}������I��͓O>9�E�#f���>��'�\u�_����MB��Ƚ�D���0��p��Ɖ�������o�F����]�E����f�6����A��7��ډ��g���I�f��Wpw��E��+��I�˿ �ͱ`5P�ֶ�D���u�u�=�uTe�hzw�vݗu4�����h�i]�5��Q:�7��y~E��o�D��y�)�?���6�B��_��i�Պ�x���4������[o]R��,�U �.6��[�����L��ݺ��;�B��g�qƊ�{�?��]��#� 0�´�`��&;�À��εO��o�W~�[l1��bo����?3����,( ��߾7��f|�C�����k�J={	�ߝ�}o'��K��$ʲ�.h`��A��F���!�5�&e��Q,	j�,jL���s�]�-�	��*�H�"XfEՅe�]��c���Y8K�V+k܎j�w	�
Z�&.
\�~����  ̼��&���Fa�Z�S�n3��l嵳AQt+�b~� L��K#��������qg�����:XEc��K:�bqmvoĐWs��}j`������gQ��E@��.��r�%�\�;��#�%]��w�#a��Ş��X��n����򗿼@��2`E������|{�����K{�@�Z�"s̽��X����u�F��� ��'5f����{���'s@@��v�s�5r3a��eFnm�}����:�J7#�<��W�_H�� %t?&��H�Hs@wUk屲�~sp�A�l�̽&��ְcM��+sl��#
�������e��ڴp��]�I��B������aZ�dn1���X�v$��E�<%��Q�O�?�~�ݻ�{ڹ��+ka��k�tn3��RG�� $�,�-�6
>�4t��1��{q�G!�o�ha�@܅b��m@�����:r�ھ_���a�Ϩ���H��J������/ͬI:G�@.FS�)�g�˺�D^CАi�Z���K��	�脦2 �� y��Eo�a;`1�(��V �h��6B��z=uFPG{�[���4N��
���&|�xָ�^,��Z��ڷ�@\kdw�U��6�{+L�]T�	��Ӵq�m'�����	���,\ۂf�]�W �d�R�sfsS�B�D�EK����晹 C���(� ��9��;>�S�{1v��P �ť߽C��]��<����	�m��{1�_�����M�����D��t���{��|hy�YֆK�F�����h�C������w���F�h�F����ɛ^i���wf���Qڮ/�{;����{0�����D(��@��1��u��|%�|OJ|�˂�bQ99���y�������g`�W��B��6�������$��,��C=���n�π���Yj�"�UL�A�ZW����V��߲�˭Z��գ9���N��,X˷f.^��}���s�lF]��M��.���$X5���w	Ыy �7�4�>�c��\�1�ٵ@���k�.Zӓ����c������|ǂ�w��g����Yd�c���i	��)m��/�U�yp��,��H���C}����oF!�8��s7%�j{��a/&�����]F&Bׯ�v��g:�|�~�O���x�O`j%�#MPR{��x�UW�D{�����U��g�oҁn6�k|������BeX�y���䘊�T����ۑZ�|�6��>��eWDt�����?�)	��ԝ���u�ȼlϩ��F�8\�y������N�;�Ekٚz��[��]��]���2����y��Q,�gM��~����=��	Ыq6 5���9�0��������p��h�H���|�l!cb�ێ;�8|��~w���n��Gu��h�[#4�5Z���`ca	3
������^4�+��%j:K�\���\�(�=Y���~�X���t?3o�� /Gg�9�ҧ�1�_�F�1���-Ƭ9��!����$pi�jG�m]m&��$h-�ڸ蕏�8�}�������T�@5.�y�V�}�})�{	������g����s��Q�^Π`�u#�?����|��
�@��'�#����h�w;<% ��J��%M>��:.��--}+��	��-�4�j�	Ы��HƍI��V��E6Go*I��j��M�����?����QL�&
:<��aYU��O>y�s�9GQ�+��p���k��R���95����w�%_~�I'���+2�p\���m ��a���t:�,m3V��� �B�����g�.�������@�J�cWȒ ��5 ��zިe��*�cU��1 �&�����W�v�p�`
t���*�F�{AQ�S4�X�Kh��=#�u ���0k}I�v�k�oo���� �/�_���}*V�L(�KsRmi};7�fwӪ��Z v�:_�����h��״��'%=%���U<��Յ�"룵�
�/��ƥikqzkB�2iQz�C��6濰`����ɝ���;��J36Dk> �|/��ǈ�u-N-zk�:WB�L�,�w�ǵ�_A�,z����׺��+wE���uc�(������V.X�}��'	�m�e��J��3&�~T���)BS����,[U���x���E(�) ��4�g(���ǫx�R�G �!�@6��]�bM\J{d�X�w[�.(8S�=�Y�1S�w*��{�m=�k�d�hy��x����h��^� ��h/�zw�}՞�%@��ٖ �
�O�R�����j�iM�l��4-D��b�)L��Yhc9�^R��p_@+���������;)#�rMS��� �٩)���Do)?�c���0�	78���[��nD�jS��qS��7���
�R�
f����<Ep�0��7�tӱUH�Jo�;� �;�}���8�Ȗ	�5c��*k�y��d4�`F �\�%�q�%E�J'pj�\
 ��� ܭ��h��R�Vs.
��_�D�젶<�7n!���6+B�V��	�����5����蚋�a�Y�[Z���T�F���m��U�^n��R6F���U@x���ca�M��*J���E�{i�	m��v�P�yQ��Y�7����^�S &�)���b/3�;%�Au��l��_���^h�3��^�>��w��k��sߦ�\s�.,��H�Zw�[z�bw�G������&օ�%�z��+��i�{�����냰l���o�n�:m��W����6yM�J��E#O���`��KM2O�"���Ű��p���ֲs��S�>�@�9�|�������6�`�ט�W�Oi�;,k����W��JpWQ��U�F�(g�V��ؓ���ЄL�^Ʉ��P�iu{"L�V��*K�
�:�䭅�E����d]Mp���2 `6$�eW�>_��Z����,@���:��[��sx�{?@^�e�m�ʅ�U�����C���:��*n�}�����>gqߋO�<���X����\��a��M
�`����+1^��|1����f���Kֺ ��� �W1uހFsY���"58�P ��s���;)���+�Yw�X���<�+	mYϭ	BPۏX�C�� ��,�M¹ֽxJ�<Yp��N�ev��^�޵+� ]�p�	�ے��:�+%�:�L)������<����/���C���j�u�IJڹR>� |I���"��oh��p����62�����~�q����������7-0�x��iv���y����B��QI�+H?���n�E-�6h[��/{�� ��ݿbЛ���t7���~kÖ�1%� �J*:��m�д5�.�m�p�+�ٗ�w��Q�����eL�J=�gذa�Д^��C �;,f!h��潀7dX�B3*5s�ʑz�>[cV���'�K�����`_�y\Gm;������mef~���NFM�K��.-]�9�A]��BG��bv�7�[9H�^9t�EN���c��+�Ui3inh|�K���ڮҦ��MP��2o���_m0' n���_� h���z�����9��i먗���Ч,�g)@s�~������$�
������ѿV����T�b(�$���ܬ<��^��\K��-0��
��%ґݤֹ�����1-�&�x3�|��2����د)�f�:V����~#��)j���|�����GX�hN��q�]�Q{�ˌ�כ�O�ܢh���w���w�������������8���H�r�)H�N3>�({�Ă�Y������M�>�D��Ԉ��u)�p��2,���j��� �ڴ��偹���0�x��$o4�����_z�c�h����o���\���^��Y�7����1��Tބ�ݶ#%mLgK�V���0��u?:b��@��>�x��.�J݇sI�j������8@+?��[��ʾI��v6=FC������^�r׭h�7C� �j}�t�y�l�����~#.�u�)ݵmz��u�o��ҦY�p��?�YG�~+�D�/��u䋗���ծ}�.r�5���^ɇ.�;���=s~�!b��G0����O�j�@�� 5EW:)
	uG@b!���4�\M��$Z�py��XN���C~�y�L�_�*���.; !a{�����F&{��.]��|����,�iWR��JL�3����)���+�2�;�w^����٧o����5�y?Nu������h�䓋^���`I���XO�YPq�t~1mM���Y����X��x�L����w��\L�ti�@�@�V��w)8�]Z����`T+ �\�Z��.�m�<�\@W5'� ���C���ģ�;�:d�!�+�����<��|�R`X��}I�����a�^
$@�Cz�{�Q;�H�a=4�6�F�UQB2����p�#ڝ?*�bЋ4?�ۤ2]��{���~ �b����.7���|���<���֞�����7��5b�M69����cD��&5m'���ėp�-^���T�:�{-\�j�?��;X���WR�()~��VG+��R0��.��r԰+$�;_�x�{	��79���9��*]�(�;
�ͺ��9+_zc�U�u�]�U<�w��Y:Yn&o�
��}��(J:ƚ� ��1$�:e���?�rj��S�w)1�;]�h���z�ߕ�W�dN�>4W5
��̤]������Vk�Y������p�U��Z y�P4�9����S�]�k�@���k/G_�\:���&���]w��L�����H��_���� .���@/��t�ܼ��<�	�\"�_���o�H��(���������tr�-zN��]�ϦG��	�(��0��"��A�iMz%
T% �'0��"�-��@�9���'�;��e�7�����Hw���nݺ��Z�u�Ն�_��z��6�FQ��/]�z.4�ݸ�˛�~W��Im��	�gcF�cل|�bq�D�$S��嘙� 8-�� 3������u-�ќ8����RY]�\0Ҍ����������4����h��p���_$�m'Lu��̫M��o�l��k��_�De8e)�S?�����
�[d���PЛL�����ń�Z������	_"��"4�)�1a6�M:5Q`�(�y�+��g���q�tĻ�zc=��d�7ͱ*����)�vسX��dE����\�B�����:�p��,���jԺB0@�{g.O�>W�?{'@� ���s�֘����UG6>���&	U���H\�A�p��@]`.@U>'>��^x�E�z��,���}�u�����`�R?�%�.�r�-oA��K��AX6��ʣ��jgnӁu����پ�x'������oQ�uFIU�)��|�B�#���
z�����QG.�ꌄ�V3��X`n!�h8c�"wk|t�`�C��� �5ަ��G��7����毺�}z���#6����ha��B����XV��:q�4��B���KO��W��w���'N�^�����l�����b �̿�X�Ԓ��0z�����Z-�5����k�q�啪+E������ru�7i״�%���O����eR������1����`�J���{�@.�;��jJ�^L
�"d+@�;�����5����S�O�wz��x�y]B����t�=����#�.���
��M���^c�O7�2
`!z�0�5�P��E��%��=�sK��{�nk�6^��LU�h�#����w���ɸ،݆zH�3A��.� f�L���4T�hx�u����*��o8�,M��"_9Mom����D�7�*,�R�C�.��HtK�.���O�Qڼ� ��	L���uܳ�9��뷼��t�Zo҇'Io;�E�ÿ���#�6Ud|wk�i��]�ɾbK�y��w��u�ꫯ�*EbJF+'�>9�+ �M�h&����g��u���?�i<i~�⺸��i�|B5��t�D��R �S��w�h'��P��wU��сm�]�M��t��8�q_�e��]�q���mr�;�^�q���t��2�k��Bh靸w�j��	����_Y�(Гa
HfE]$��_������l�r�@��I�;�����d��i̛��]���=��U�����m�J?���#��7[�����a4�R�̩rj�>x����.�W�{�k.���W>�裏��)8�����.h e@��[ \�u$�S��^�e��[B�^z��Ua�hp#��T�u�&�PI@���>���J�+:�m&% ���� }��/��}L
�l� 8G����׊y�s]�F}��"�&_���u����VR3��@�r��א෵x�&=��'0�)��,ECѝ�&�$��ݚ��'���\�EڼL�.8c����x}� ��+ r	R�{�E�>U߮@3� �e�~2m��x����q1%����k���L�#�Xc�R��b�
�B`�2�EØ�o�H�Z�+��"߀�+�����y��H\#Q��(���gU#t����/>�/\��X����r.���)���JF�ҥq�W� 9W�sA�.�8����n��R;K�^E��E�� ��R�B�3�V#F�8 -��w �|sI��e����8��e����[����djwU2����.�kc-v	�_I������ޱ�>���.l#�m�b�f-K�W���=oͪ��HQ���7 �����͎nߜp�	�75~q��=R�sa/k�v-�&����]D�[��쓡�vB;_���%�`��l�@y`]O��4��v���26�ۊ�BT�i�J��:�NF���׹ؒ-�I��n��� !B�t�˗���d�h����0��"?���]�I��6K�p��&.��j�^2��̴$p�y</Z�E���l���Pj����*�(@wh���(�<��s��WY$7�O}��w�]k��wߟV�漅PZt�6�^,�jM߁ua����/&�z
ДL�F��1����>��2_��7�qV���%[��gw��h�#̜Gf�gհ��-��mK<9�}׮����.@Oi��S@��i���苷ƭ5$�_q����En\��io��	��|�ܻ'kv�����~�/L��ӊH���8?�{c&a33i|ލHd�7W%&�~dS�4�' ����u��.�~�5J-�&z��dfM0z�{� t�!����￿#in=���[��zZ3����{wt�5~	�#���9w���C9�]�^�)Ssg��=��wD+�z�w�_ܯ��-F�1p�]�)�01>I0�y0���C(�"95G�t皤� ���NS_���6 �(������lӡ��X?ST��U}�۲�KB�~� ���m���.K���	��"�&
�c|/w^M����;:�#�iA�����g=@���5d�
�i��sYWi�rK�������:O~s�x��I��w�w��k��:�� ?�"z��C���G� pꩧF���nO&v������B)���o���~���.c�f�T�<o���m@���XO����y�P�T<���͙y��h�W�㻜�|�8�(P
�I��G����X�n-�|���@
ʟ=#�CmOuy�XH� �,���f�B<Fµx�x�x�x�Rؤ����w%Ǐ.Z�r�{@���b�ht:@��&��zK��D�|�ɫ���w���s��'���MjC~v�h
\����d����9�1���f�/-����b���y�y�J���,����ff�i"�D�`�2���}A�8��=Iw��'���h;���Q�����\��x�On w�n�����4�<���������W�@�P 3��d���m���w�kQfZ�]�N~�����=�1WZ����y�:ڵ�=�<��`_>w�;$@���6_:uΗ%��t�bMH�����<��+0Vp����] l>�5bM|��\�'i��Oں|�j�ҵ���˾1��u���T��q�ע��_ �����h���6Ԝj_��N^�t<��-�����)%f�~VU��X��	l��L3G�[�rMk=��^Zز`��b���elm;�����I�v
0���%�����lZ��X3u�Y�_���^sޯ����a�1�܁��z5g��ˋO��6��vAaZ�S߬v��g7�/�`��JK�o~�إ4I�C.�����7�L�Dif>!���W�Z;�"��Hk}V�&��W`�ML����@����������5M�>��=~��8��%c���H�2��R�}��!@\�����v���R�۸>�>��c�`b����\,C��gֳ�y��r�N��M��qC<���I��1�M-��O�L(� |�.< �j�
��|Q��u�+6�Ã��>�W�Q�< 7;�m�����w�'��������Ε��t�Z��Z�CW�oG�H�
��|��+��ľ����Y�C�b��
 dVX��X����CEC̆A�������c4�8Zh�!	��a����w:�>���������A��q����mO{]] �f{�y����g@�<�>s��V��*�C��4u�{��'&�m�z�A���h.f#�Jn���s�Q ��&��
���5�\��6��Tb���
�3���1��ڲcy�����&��G l��6�%a��zu�۲_݄�{�q>v7���B���R�Th�ؗ�D�����U8+�+@'��1u�7 =��:����C���U�P�8�|d ��.���\�EmI������)�4s��M��m�%�ih�!�^A���COļ>��N;��1���L�jOo��;̑�y�ڏ �] ��䩿��
�O�6M`�2�4���M�"����z>[B\_���u��g��U�N!�)�S�����ZQ p�/�����F�wĻ�N�9��\A���\@��Ց�p.�\h�ħ���jm{3��������Ֆg-���2�	Ыp�7����%y�;>�����Z;8
�*����-�����dzw��5@�v����&.��"��վ��\Y�i�4��G	�;��s�}ʹ�*-IZ���W��uo�O���γ��l���+�� ߵ ���oɔ.E�j�裏nv���D��${[;Ů�r��S�DCd<��0����ϥ�N��
�Fj��) ����1�&w��4V�:<�	����z�p����>�9� m�!OI���2��O�?�����a�R����rş���Mp\W }(}x���7��q� t"���{QnO ��&������ҪeBRT�rƽ銃ФKS�����.�@���be`����&ΛV{�6����lp����1k�^y�G�ΚNis ��\+��uz���9�������L��'�|��̡�ʴ1����W�/�Y6�l����\tG�Z���=� v.Z�#��U�:��)
��<#t��PBm���U��s��z�4������Nu������ƺ����M_R���\�����<ﵪ~��<Y,���ǧ�����d�S�M�yП{�vWH1�]X�5�]�UA`. (��
��3ӻ�޼�w�9T$������mf7�[3���Kڸ�-OϠ���4��7"�����}X��&��}�6�;g=��+��8��K$wɤ�Q$f0f��(>�1�DW���(v���Ch�����W�Yn�᧥��R*JxW# ���5�����w�����\�n���݋�9����ȫ��e,���ڡL�#�@)Y����x�֧:)�R�z�#�B� ��?���t�g���<P���P4�=0�w�Dͷ	͎�xsi��ȕ��7�ح	�%uz�H�j��CW`��m���p}�Ŀu���;�`~��n��`hs9��)_]����y֮R�3�ף��?[��Y*`��{�5����/���0Ơ��A^�&{f�Y�]�M�`)�Jl�����}�7>*�yQ.�ԩJ� ��k �+���eۤ�r�Z;.�b�<��~T.�Gcn	�[��=���hv݃u�1ְl�2g>�ӧ�͜�����M���)l�q%ʏ�^UD�yVC��XG�>=���; �m
���w,4���eZ�"3�}���@�AY�&�5�]�x��#ys[@�}���H��k���D��=�������`����\x����MYj;���D��E 9���U4?*�Y6U�V�Q�ۡ�q����;���r	11��0��N\gP���J�`j0Q�) �h�*$�姣���R�*\eu����G/��]���?k���[��y*�'T��6Y���륗^�qF�� �"3Z���ծ��=z����򗊐��D��I@g�N��?^y啝 �V���3wj�4pi�M>&jf*��+yMPk�/"�k�uޥ��T�E!�_��>,Y��wt�1�s��,��D��_@z!���ݻ��$m�v:�;��ӭ���A8��Tf"c�B1'�� Z86��r��B1z6W݃�/�zs��n��>�T�;�3Q`n) �	�i"�cs�#ڝ?������� m�:@ۂ�2?������w���V'���.�_����x����u�ׯx�� ^e�]�V۸"�ƚyByɤ����U������i��� 4��@�kb	p�Z�sʙ�s�a�kr
�哲�]�)b����襽+`N���X�� x�̶�Q��&@x��Vg�y���u����l�C�o�sH-@蘛��p�k�&��������,sz/|�u	�Y�{��'�Y�P�'����Y-��Q�zf��x?L�̿�A���9�t]IR �x�Z`}ԋ�]�n̛l���Oʄ����:3t[�n&\�
q1�=7�� ��"��}2�;݊Es3��~|9�A�SZ:m�A���$xW�M�y
�1�6��!EM���d���b�TҾ%-
0�M�ʹi��]=/���#�]����4��6sI2���-Q��K���Gy���&c5h�f~ �Z�r^7����]N������h��l��f%Q����V��K��!�.������/2aH�Ӹ�.:�~���:"��!�dR�J���/X7m�����D��+G��v)�v:�����Iy��j����ڶ��f��1�2�}<m�!�K��o ���3�~�V+>�@�\Y��:W���U0�晠8�sU.3�� v{M(MJG}
4��֦h�Q�޽{geZ��^6��<r�/-\����L��LV�q�L��V]u��ټQ`�_�+�!{s}7]�k��fnm�&+uN���	�v&�vr��9���H�Gic�Iҙ��.=�rU=.z^Y@�6^ ������U��S�%A���V����X��9��/��R��5n= �~yQ���J%��d�y�4Wct$}��<�J{$|����Ɂ���k��Js�)4ә���ZzU���\�����YC�(��-07�: ���7m$�	m �O<F�k�K�Q��Ak�����)�0����?���0���0�m-lx��qYX���X>@:�ϰa�.#]�$|O��ޏ��SxޡТ�����h>;���/�y9o`.���ԧBU��S��A������K^��lf���A�2�K(���</D#����Bk��Y�NL���nާ�U�b��PՈ	z	����{��������w��em�M;ϕ��V/�	}���� �'2��EG�.���uMP>�,2o��ɾ]��59�-���ۿ+P�b��>�� z���V[mu�'��8`>�R��� �wvۑ�V�����Oo�jI97K�ND�����T�\��^�%bFVR���}�����J���Cϫ(v,&�R�}���LRo+�ĜtB�^���|G@�+�!�D���^�T�_�{�;�����kضR:��&Ã��ZVn��!C��D��묡[�������K��,7��)8�X�x 0�`"/is�&��1���Ȥ�&�L�*�*iVoj�p��I�kծ���)Px�]����~���u�]c�ҧt[�dǴÑ���Js-4�-��޺�����BǱ���WU�����s�%���v~!��*�W�y�JwNk��L�w5<���a'l��Fǰg{*�:����P ����u�}#%�@�˴����3%$��]ʵvy�%fh0JI�Y3�-�u߲k�3 ���Dҍ\3��y��:�X�i��o��pi2�J�y����u:���^�2�h�7�����gґ�K~�L��#�V����k@Whj���:�.k�E �O�o��~�>���~'�{  w��A����rG�뾎dwiؼ>�,�#n����ޫ�|����w'������,�����o�.i�xMAxI���˵����}�[�@�Q�@�ڀ�J z��?w��y�֕6�?Ӗ�N�5�f���,�v�?���^��s��C�}ξ�c��B(b���ij1�7V���j׃x�v�G���Q���	��@^�v�Zە�\ܦp��I�vp ���<�����!ߺ&�$Ro���l��>�#8u~,�=~f��ۉ[o�uV�����s�a,��XX�'�O�gWs���Ρ���#���+ϖ��"_W�|_�B��n��g��&8�M�jm#���%�Rr�����0੏�B"л`�^��֎֑xQ�UO �.c�u�`�ܧ=��)j�Ef�-�y�y�\6�별,lo�e�f����W��GQ��p��x��1�N�焠� ?�B�G7)I�l4�}�
7E���ɛ�a��.�[�n͜��s���C{>�A&�x�'|�9M�9њn��v�I�<��	,����v����O�"o�x��MY0���e����ԑ�s}'lR�}l0rx��9���!���#F죅�qP����A����?��J��#��G\'=j�(@��b��~RX�r���=m%�������s`�ε��J�{Y���Sc�?wn��sE�#p?O��`\"�P��^\Y���wૅ,ͥ�q�_!B��*L��tJ��GT官m�h�x[Sdq�����������D���_�k�J;w�b��뭝�������6��t���Gh� _}�A�(e���^�4f�����@AaQ��o)/|3���b�al��J�G�O$�m ���G��Z��d�eD���:�)	���s�PL�琧?�#�:Q��(��>��*KW�K�K��B��A�Jv��n���<h*ז���?���!���w���\m{c$��z�s�L��p���Y�ؗ��l) }m9���K�C%�]v�`"ڏBr���|Îl"j�K;W0�����v�mO%Xm�.�B�)�����Z$�ծ�t����&i������~���}�z�������_~���ӷ�u�^�V]4��f,8���O��"��0*��]
sJ��oP�u���[2�v1	G�J��pD��4�D���{�A�@����x�>�[ t����c0��6g��*�q'$]��)k���&GY�]�Y&&�o���:��_g�~S��_�W�3:7V�s/���\�}*�V��tN�)PR�N�x|秒����ĈvMpi�t�^�nd�n��;��3h�u�Nu�����FMڸ5�H��ޖ�m~w:�Ih�����=�h���t�-�b/�#��Cu�}�y^u֖�gK�y4�$|T��Sʵ$|J������"V��$����ͫh*��-d1L��a�����pO��_�����(�q'n/�#^!p��Q|����O�O�s�Hgʌ��Yֹ��#k4K9��:�>�1�wwo��u�������p7IU�*%��/��<��� `e�u��B���'�GC[�Z2Aqh�m1����˶:�I�"����e]5��ȯ�	��f���~��1��O�FG���Bf��d� ��\��R�M�����Ŧ(g`f�J#Ć#��3?
AcC�Xt4��U���ܥu���$޷�}Ė[n�Y���\ހ<�� ��	��l��+���\WD�/����S�b�j�����[�%$�k��D�y��/H���X	œď\�R�KkO|����g4�l�j�9�	~���Y�}�k���x�'�������2v*�BC�P0�����6�q<&�e��TGV��tޟS�$4t�C��v �vc@��5>����]>4�h?b2��?�A&�t&qA�縒J�
�]����E*�T$IU/�w�6��.��6�|�,"� ��#h�K��jQIu8K�^$y��2n%��R s4����톹�x�@�Cځ�Ҽ����5z��"�F�qNO`�XR���)���.kl3��%h0�Q ��%,�;;8�"M4���w�u�@����i�h�J)�vlq����9�U��W ��zX�ƣ��Q_l�w{�irIk�׺�r��蕸 J��C{(�W��}7��󖚢��mi��d�����p��[(z�E� ��t7Л�<Mt����S�4]*V��E�A\'���||��{p��5KMs �@�p��t�'$��sR��b�-fk�T��W�)6Vi�u�@"ُ��}E�<J�l�k^Ȓ�u`>��#ٻ�����7M'&
̇���m���6wN��C��t�7�Vf�����y��VVr5�ا�������?ߔk���)�@8���hoE�d=�4;ÀUr"����]��Ӏ��}�ѧ�f��t�S������Q~,f�F�&��2j�sM�<�sE��y�/�/]�;�BY�6Vr*�&�77���+V���j�>,>��$�	
��^x����&|���܌�UF�f�k���e�3���9��^�S��� �����J�1��B�2��:����`?d��v��=�%n�(�'��4@x�>5��5,����ua�ۊ�����_-��k�eέ�kH��P剋�I���E�/�C<Tox�X8+��k�v���K��{�v��[p���b��&F�P���y7��O�b$��.�j�L�T)�#�Q?M��/��^>�-1�7�E�`/G����}�����7�5��G}tV���f~ Q���3MT�I. ����s<��ɼo�ӿ�s��	3�	lG����ײg��	Pϛ5?Sd���%1�Yz%
$
�90��t��ōԛ�o���h1�KO�i�T�F��5� ]�� �5e�w��>�����m&������qʹζ��vgЯ��Jus���-
��wMs�r(P������w�kI���ƛ��Y�a�W �aj��]�b���\�_��Q���\�l0v�9&����/�p�}"9&��T����v���m��Y��"Xu.6.�)L�;�]
�9�.����o��Z�9%����L7�^oӎ� �_O���x�*g��V�m
(7+؞ �"=+mG�{�&�?�X��X��'�va�<�m��͜?ı@���o�g������txq/�+FS�@��ϬO�[�#�rP���t��B̚i;�3k
-�#���f(�:��	�D���7G���I�8��3�|2>6��NH��z[�T�z�;��I-��8�]��=�#ndM���|g�N�/��&1G��=	���}T��=^8�|�Of=,5{�~�0ϝ� �5S�^ϧ�7n�c
�J��w��1��.:t������f���(��@{^����:d+/�l�Y�ғ%�[>�g��M��,~�@�E���lnR�x��
��M�#����9�ܦc�l
/�U;YZ���aE�;��Ef�Pm�9�_���(J@L��u4)�=�]�E�"I�Q�y���DV�DQ��
sq��յ���LY�Ȗ"9/�V`̤��{���_N0�Xr&� ,�D����.��̮�&m,s�s��4����E����3����{����Beu�hA=�1��b�g1t��wv�:�s�ꫯ�mZh��� n�n(/��sz;N�{?8�=W02 f���I��aeG|Q׈YS��P��Ж+��N��]�o��hv���l�9`����ԖA}rttN�Ӏ�G�����V:��(Pt��O�Z��lL��#̝�am�����Y�Q
�\@���@ ժ%��`��As�����1�N���Φ��gb���H�w�v������hԎ�a;��u�k������� ���w�a�w�}*R�y�g���ͼ����:b_���h�q��$�!5�O&��4��n�P�4H�K�N
�eץ�������V�lm�%0���h�Yo���Ӽg��2�qz��*\�y�a�sh����;���҃~��/��w���� ؽi=�'������}���@�:`�&��r��7�$�v�J��U4���S6>�e17u�QOp�������# ����@8��<��#7衇����g	�U\;)癣�����P�$�~��E�{���Jo
��7����.����#D=�r�quM��%��~�S�^��� `�4)�����q�J�+�[ſ��H� X�Nx�Ѭ��Y��&��0[5u�>�w+.,�e�VE:�k4����(i�,l��ﰊf��Vv��;�^}q�oC�ܮ�oQ!���fJ��t�Å0=LF[GnJC��Bz
��ռN����O#-�ی�P����ù�c��@�)eZy�[������.m�C���&�g���:���s*un��Ett�9Տ���	�^.��'����;K6@�lN��85͂������e���m�f�+�+Q Q�b@�莹�(\��
xmf����r�����)W!<��w�7��k����S�z�Kmx�[�t?WuT[���*��2[���{R��^��wD�B7�1ok�]���-�[�c�(�Κ��	�j�v~���!j=3�ڏ�	b_�#��]I��;()Z�����I�Ш�c��!�����9PNB����E������j�.X�n:!b���y��՞&e�]�� �c��j�t�O=���&�^��<g�<W>{>k	�[uN��r0�=C�w�}�{��S����>����՜F�����L�����S�Tt�Xq��%*������\�e�>;�ޘ�N[]��`��t��� d� h�\��
m��g�WNF�E��ꇁ\�s4�5t�fxK/��m�J�?E�l��<&�u�Z�����YHڹL���L��(�z)ј�m^���L����M� lv*���r���~�s_Dۼ
0��nbK>�X��Oi�[~s}���)���/��/���b�
�Òq&��m�s��b(��]�y�c��Շ(s 9�E/����͟��Y3Y���֛�K��.Z`��O~������j�=���x��N%�eM��_
0���=&��9�/�Ze��q*�b�|�Ηw�1��4sA�Er�%�ie�a~m�( �����J��?�D��я�$5ѝn� 9����D��?�g/�A��d��3N�pe8��X �y�K �e���%�����S��p4��]�A��<l׏wn��Z���`~*���U�
�y
ǜ)�9�^�A~6�{I�Zx������ D�K�]I��^���7�Q��;���_���Z_Zkq�)���rW��t>��p�����P73�q#�W<RZ���L�#�S�s	��U��'�B���j�ho�b�
xz-����;]��zW�G��>+����E�h�;(��{�j��Mۏ$M;7�OZŹ'�|򛅏���S��L�m&��vΥ�;8���#��G��ˈj��U��}��GP�p}�MWjg>w��a.��	��C(x�Ew&;��:wCR�WS��;f�3�6b�e�����,D93 �LLS@�J+��W�>��꩘�(0���F7�U�p-+�����d�#�e�Z�����\[ }sxa'�i}J��u�+��>s׃�9.�혘���r�oC�yk����+���4�LK7ߵ?]��?�Z��w��Pe�c~l������Z���,o�A���!.Ңɩ�^L��������_���߮,��mF�o[��ڹ>{2�}~�|�{<���1�7=묳a�m�y�9K��)hei$�S9�@���R�7������.�R���4��A�lw8	$���]��{�k� 忻����}a�"${�R��b{2�9|f�xQ��2��O@��w*8p� z�5R�szY:�� ���n3s��VJt�O/k���h��t�,*�2^�g�@]�
}͞��+��Z�r�R�F܎��a����~̏m�(�coN�����x�	P5����xk�5�8������߽�m��ijs���$ X��u��>��W Uf��׿��w����� 1I�zy"
�����r59�$Vi��*&#̤+�i�"�l��_�f8G��{�z�"��'!��L��A<��Uѯ�f���@
f�C��6���ە� 8���
��ZD����aÆ���!%�/|������i�V5en��^����}����/�{�+�����{f9�"�S~������ݗ Rո9\5
���D6�)iՁg�9w���>�x�GL��v�i(zp�UW���~(�b�!�+vyV	j�E�X�Ѭ�CH�⨣�ڇ�2ɲ�E6C̵�wW����`w&�J�?��8��2��`(���Zߚ���������q�"����lo�0�N��
����x����M��[�vĹ����x!��_	To��xYR� z��M�.�$��r�F+H�Z��_<P/k��^s�5��!��LGx����H��x���}����"P��se�i~i�� _u �`�&:�|J�;�������no/�'�x��{0ɗф�����wU�D`q�&��;��SOݙ��3�����\��s���
i,�Ih��9�X�O������1h�[ �7�ը���ZP����Hn�w8�2_��$
�>���;U;�I+�KV1i�Z{v-:�6�s�<d�@��a�ֵE�'���f(�M�I
���+=�>�|���T9c�7��"2千}�8����I��:����݈_Z��Ʒ��Zc�Nu�aHb�;��mMZ_/�|���4r�G���_���MѼ�Hud{��$���qE�3�YW\q�H����&��������JN�h�4"�GӀ����a& �� �%钵Zd��� 1m&�oz֋��J1p�[QS����5s���ś�cb��Sr�Q˵��h柡h�FZ�{�8��gvS[D��\e���B4P�ZhP�gS0�ߎ��� �x�+�I9�=������������F�
��m��o�z�5�h�]��KҦ}��p4��B��h�w��N��#i``[����Ƚ5y5�}]4�ۤ#�u�, ]�i�*p�7	��q��!�����!���v�}V�ڴ@;�3�΢u�w���q
bZP0��ݺu������<��o�N�eu#��x,c�J����:Z;��<�I*n�߼\S��h��v��r��ծ���Ej�;���dw	�o�ƕ�Rv���vU�c�)I�CÀ�MatT��\7�q�v��n����վ1�\Z̢0��A�:B�Qx���/���ҢH�-��w��5	4Y$�F�FPHm[2T�x�����iX�w�Gd�r]���zϞ=O� ���<C ����L)ݽ���*p�9��7�s�1��ߍ�����y�Sߊ�Djw"��P�klL[).6�R����R6�%*���/"�vby��~qxX{�xE�2+��\�q���ij�i��?���s�v~TU���18[����4�[Պ�-olűf�e���r�����D�ƶ ��#��!:�B��b&L�IDn?�S�`z���@Z݌IQ�+��ɦ(�&�@�H�� /@g��U��F�Mі�=Y��#=�Ciػ�yR`uh���`�7�����P%��0��c�+��j��g����7���)�+�=�*���;`k,�!~#MZq9�5��H�h�A	� ��l�|n�r�\h�M�!�ۺ�e쟐�;���oFc\��r��.L�W%�[m�����Jْ%�j����5xg�?ލ�ͫ��MU�fs����ז�)�T��ڹk���o��z�w]�3Q��Z�AL��l�v�v�������啉� ^R��8��v�ς��Tu�lҸ�O�̾�xz�9�<��u`��IĢ���"R���R�y��X��B,��h?���]��t܍�\�,��@\��@Xk�U5����c��n�D:�����* �6mFW;����apj�����Og�W��+��k�>��p�ɔ	41J����"��2 �H~��\�
�L�h�;Pl�YZs��s$�h�q�}>�����jx�}��΀ѳ�_dm��l�w���KV�I��h�.~�6,�J�T.6��)��_��k
�M�W��^z�0�b�/(fb_��mw�o� ����^����_�R�Q��!SÉEH��-)�<��I����f.���(>$�#�#�5/,3_����[��p\�Am����r�%-�0s�J���i��s�ATe�v����FfE�K -ގ���_[{w1��];~�Kǀ"��R�:&�����{�f��@���A� ��sm��c��cw���m��N�����e��Avq�Xk��]/����͛��o�ȔS����Yp��/��%9�c<�,*�����.��� �1�H��������n1=[�K�@1S  oA�����|nkaZkϹ�yZV���B���MT(�|{���L�?�eA�A���(:�G��]j�����X$�=���^�9��	�FC �w��ď]�Ӂ�{���5�{��S:�n1�{���� H3Ev�w�&/�I�����0��@��%��~��y�v��0Yzx2�On��v���$0ش�Z�j�l6�]�����,�Sw�a���m�b0�-����Ki�X3�wA�^��E�";8��6��!����5�-Q��(�rЂh�](Lu n��Zc�'Z{��Vţ�����HO�����c�����=����g���jߑ��Uٽan�g�����t��St��4��E݅�����M}q���ճ��)l���qad��ҫb�6@g`z#q�$s� ��+
ُ�dx�	�l�#`jߊA^�E��,�ټ��]�е���L̖����y�M��o�����S#g͜������`紕����c��P��,�?��k�}<�]Ӟ��^��&
�> �6h�{R��,c]��w�c �֞���ŏ�?��U6�:���YQA�-��s^�7��ږ���I�#��<w�P%9���`n��4�ȏ�Wm���K�곃�����u.��32�-�*F�jt��.��v��z�����A�uq�|C���ί����k|��ΜS����s��5s���^%9kQ9�˚��a�c���}f��+Fʚ9 �A%�������(Z-p��X��+��������iw�y��k��鮉�O�'�� �P����Sb].�Q�p��t�?f����ǦPOW�(2=1�w�R[z���ީ�=�����@��W�v� �xt]�E`���:��tco֒�H�Ϊ�O:�7
T�3�;�^E�Lڱ���$����i��8@�\sM{*ʄ.�� `Sr��	�@��ǀ8MzI�.Eh-�~�<�k2����_�9�J�/T�|��'U��(����G i]ځ�P��z�f �'���g+jA�2��H�*
�1w����d�O\Pˮ��bV�] � 8)y���D����f��W��q}�mE�m�;e�v0p܋�����,ֹg1��Vݥ�yΆ����s�U�]/�y�hn��ϼ�ʄW�N�jt4��
�p���Xk��7��z���5��̊L���	�t�3Ky:
�\�ȾM���i���`�exb�E9������i�P�%>�}��4r��s��+��̣(�x`~�"AM�D�D�٢ t/�`GM�=�6"��i�1�\Z� ]�S�=�|4<�<��W�>�"7��֏��N��ߒ;͛��H�K8��'K.����!�Ҝ_�>��9h���Cw
��u�Q^	.��������z�����*8 U��S��)������F6�x�����'H���3�<�7!1A�r�hiٞ,־�w��j6���9^��gk��"���t��E����n��nGr�w#��Upd�v�g�s9�f3�纔
p�R)jr�G:-Q Q P�b1��i��� �����3�K[�ړ m0������7�|���,�P�+�P�v��<ȕ-��⊏ꞔ��-�D����&O���4P��rY�X�St��n^.:�g9�Y�(��j�9J�U����1�kr�?" -p1S���ƜU��Sv�D���)i��;-�fwG�{Y�w�d-@��\x!OQɢ�գ�<���7�����j��m�����#�O&=�6J��KI����R����� �g��⋛��&�r溓��1�W�J37��#q��w�-��n�*����F�M0Sב�Z<N�+� �,�]���L���؇�J�V�Z��ץ��᧰����� u@��+�g=��j�lPwʰ�S�熾��[�*J����*t�%k�?�	�AY�t&����`"N�y>�`|G�rm��%=���b[����\�AD�	ĵ���k
��'|*s=cEk�>|�0�#�Z��8����1�A���8��.�m^�煘���)��|0p�,�ԙ3��\�w��5� ��g���*��i�y�½�޻$f�#�x{8�-�"f�vW\s����%��'l��5R�Q�uY��ȷ��V��v8�������L2�W`��.�����)䌷�\������e��]L�����ۡf�຦���v��[��5ZP.&�klnw0��wt���;8,N�<��6:� �t���)�3���;��)A�'f��\�Ւ��?��Q����!m�:[�7�\�@K����5�&(u��b殐�:>7
Eݻ�{MRC�C��u�u'�\��Z�;�����g�Hp��^��f?U�������+���}��}���z^ﲀ�߾�o~)j/V�>�}�i@_����KC
�^:����n+�x��k�ߡgoܶ}9������^�:f��H���ي��Ԧs	RLRO��	�v�,�������t����h���p\KXm:�T͓&D��G��Eܿ�r5gw"!���&�c~"I�q *N!඙�V���.��b�DZ�����}�t~���R �^���+'����_|�~�O|��X	`&�o�t�I�y��%�X��d�l�H[@Rlb������]3�v��������ЖYg����z`�;�9Ty�Z����g
��"�Ӈ�	x��j�w𜳺E��/z�,eA�z��m���#>-�:߁q�zҳ�lm����ǫ���H�U
�,����]5p �M:�Qf��n�xr2d�dd�O���K.ّ��Gߣ/�5��.2��&�'��6��hvGY"=���*4ػ?��Vpz�K�7Ѯ��8�^�dfSѳ����n�ꠢ'b�����(0�P A�. �KU{�| ��|_ � �i����E�l������z�>��s5��?�c�����x�)<��y��Hk�.=���u�KZ4��J�=Nb��۱T؅G p��.��h�[b]�m���7�5@���֥K���ʹ �~���U1�O��S�X�۠n?�����I��kꏃ�mY�[�� �t��-ZjU�sv۬2@'�����Dfn��\�8�y�m$Ռ>s���â]�ڴ�;�O�s�^y쏱��8�� q
��!��D������~�m�?��õd�1����#&&I��?������]�@�=Z�N�@�( 7��Z �)�&��:��DZ�'~�|o�l�̓e�OSM��i�����9�o��˗��+��o�2�7s�k4w�6�{��'�=B�3�y�q�=q�gT�u{��/�|/��"y5i��_.�����M�$�F|�i���i�oVE'2M��V�l�u@����-�a<�x.������;��� B���&@����2@G"��g!���9F�����>#�*�ҏ��䢋.���}��վ�XXF��Ƌ�Ҟ���d� ���e|�;�JJ�T����fY���mK���L��r [��ڈ�������a���f0WM'
T"PZk�@�=�� �
�9�w{ ��c`lq��D�	ڏk�"�����/���d���V����S^z]bU����2��-�9Pg|�fa�rpj��A��{챳�?��h�[�R����cdxg��ֺx��^�� ��
+��j%�7MB�lw�/�v�`�7�QEtG��($�J�������vg�V��w�s���U�,�E�nq�mW.��L+���Y-��$�s�ucjCKr��۬��4��:G��	֤�=��Cn�~��
/�^��L�5���EC� ��t���NO��L�޽�p��J���pW��N��~
�1��[j������!�K j��yl�#���m�����c�AVZ'Қ���?�.pؕ��c}��.g���0���ϛ ��\�E��w,������.x�t��>bV�8��ߚJ"���m�	5;�;KP�K����1��&~�Ex�8��nB�(Lf�ޕ}.<��n`��
V,
������&�Wa}}�[��@����5`���ꫯ'!�\� :�����58�$��= ��^�z�����;arړ�������M�����}���� �o9��X,�2���	]Y�"3�<�c ��8�\�۬�5s/��"��\v�e�[j��*�SY�M�$
����s�n���u�{	4�%�� k��b��cN׉u&쏵��\�yP�z��QЏ5*�j��������r�)��w6�W�����2bb�-����+�b���*��r�~������2{��?����;�U�7��?���	�@[�����u8[���ov���?/�i�J��ȶ�}GB߉(ڶ��y���L�XL�@��#���2v��1��d�t��#>F�
�q��!�k��.�"�J����M龦�g�E��Tn)�)y}�_Y$O!�^����i$�3���\
X�%��dL��h��ټ���d�p����I �ǰ�̨���>Q`N) �m
�4C�j** Ֆ5�����%��!�=Zw�͙�*�Zǖ�BS��jv�Yx�WQ�wyQ�o~��!pTiI��_vgL�SXcY���(�֚�����\�T{��On� ��;���٥�Yg����)X$j���+3��	�E����s^�������S��da�&�\I�,M{�|�#��4� `�ł]?՝�� }泬J4t����Me�*WW������o�v�m�O?���X�]b�VUxAYJ�tn&��8-H^�^Z�r~js��D�����fw�U�����x�=���|5E����=�|��#x���f�����:���1�R �p3�L����1O%�� ��vĂ
T�Zs�J���ܖJe��[k�43{��EY�mk���M}�c�к��, � ��J�8�{�s��X@�7ĂP����>k��ƺ�,�����&+�k|�A���X��K�'����Z���m~��^�(3<fv���?B�پwU�`���ܥ��#��4��I�������ϳ���u��}Mo�m��wm�	�&�'��3�U�Tx۸���Ū�c�OG�|�b.��s|5�j��k��mn�ޟݶ}�6����ũ�b��B�M�(� ǟؔ ����FY_4�6�bJz>��&F1�`�8�/��l�TՂN�. kQ�����F��yؔu,sxw@�~��e�U0��t�"��ʹ�bp�[T�	��T��ױ��&s���Q��o^�y���cb3o�8��<�~ZG9��b����O���ճL�֌���G@x��I�e�]II��ΐ9���W �ςO�=��׺�$K���:
�,f��ɯo��&Oӌ��m��SV�g�e*�˂��B�����X��q��f|�Ƌ��4�Tf�o�鹋�/U��x�`�t��h��5�'#E�#M�	|SP���`���/���q�Z:�0`�ǗY�W��R�5�+2��f����)hbTZ��<g?c2���e�y�
m�X�>�s�m
`oP��� Y��Y�=�g�}v7�Ns�aS~k�yMa�*�wc�n����qt��4�����5jb�<kM�k7�u�.*`��(����Q��B�~W��M��v����s����A����`�=GZ�I�ߏ�����g�E���I�=0_Z�����Z�[k]��K)��@V�c2~@N����� �̶�~6�:ۧ"(��~e&w�٣���)��	n��
�<OVú�"��g+�ㆠG?�����3:��,�Flw�`��Y��f	������g���k}���:���f6��Դ�����dPT��c����7۳�.���`�v��$��k�=G��?��)���`8i+�]Ҳ)ݢH(@,F{�U{R�!5j}L�&��9k��9먞}�^�^[R2(��eg4���{���s3�H�( DA�:8M��L�p������n�0�5����#�SԦ�T�F}�Q�����7a���(��)B�����������z衳U��E��*�\��������kk��Z����c���f�U|<W~�2>n�leLߡ� �w����x@��q���rKn�6ɭ&���5x��	�b��V���!����ےV�y�	�i�q�^l6����n��4�;��L)^��$y��1w�u��dLo`j?���KyG%���u��v�F���ծN������ȕnS
��ۚ�����Bų��}�D��T�������($�V���3k�1�zy��~��[0�����3-Uo�/���1k�v;����!w_�0a~`��[��.���r����3�F��>�����Q'��sTJ����Z�]`���c����U�ES=������ޤ�)�\��r�%��y ���ĩ��+�ԧhOx��Q��-���k�sS`���J��6t�XZ�t�h"�M���J��؁��S�*�e�|Z;�ئ��@�2����k�-��|O���X�6P�iGϚ3�h�÷�z����z
u�U	�@���#:hq+%E`��&��^b ��^`A�H��Ϫ���fEO6D���Z
��̥E�^Ħ4A;/��Ph&���A0�2����1G��P��Z���5�5��|c����-�������q���Q��¾̀��:����=%<�ڜ �v��cb}n�n���˚��,���h�9��J�̪�r�zv=�ֹwY���E�������Q޵���ڮ���!�!��"�=�Lo�8�������4��>�L#���t\)>������ ���I�D&</�x��5{q�C�+Iԓ����%��`��.��;�X�X�����3�ȍ�J7�o�iAkk�[��s�w�'��}�V[m�j���P�^~���IY��D�a�,�l/FH�D-,?8x��T��:�͚kd��s\sQˍ�i!�)]g��߮��-��f�-<�/�}r_b?�!��(h�/������ʴ��������٬��9��L\ѡ�B�0u9��W��\��Z�7p�>ȝg���b-xD-E��ֹ��~������ چ
�����]��zOb��Y����D�!,K�1�m�V���X9��ch�M}T]�V*��t]),L��^��0�p�%8M\i�����+��<Qt}���w������D��K��ݴ��	q�7.Gt��$�I�;9ye�m�w1�rw�L��Ϫ� I� C� ]��%Dk�ki�.k�^:���g4[{F ���h��--֑�:z����v�9(��Z��'�cF .4�G��<����b��w*��ϩn�'6{/��"1��N���{���s��`>���s �� �>H+��ٚ�����DK��L��\�E�)Y[t�6偞�mA�+�ZL���>��V�2�����1�m�����˄�ݦ�\��޽\�v�v�w���<"��%dK�p�O���sGuJ�&i��GӜ́j���.��""��7��`��	��f�\��&r7��V��W@�J�������	v�|g�Ȓ���Js���Z�e&[[w�.�9�2�� �[�]�!��'�����sc�J����5f#?p �����k�}4`��h	,\����s曖�+	D<zv����G��O��>�A���G3?���5���^j��y�s���PDw��~�Z�s-�Y�G���tQ�m/����cP��p�bt��|��>���mc�1x�����K������3(7�ϑ��hݠ����ɽA��ۋMG�����[����y��Z���?����*�=�fsd*��1y뭷Z����CW6���Q���-���g$`G��N�uPt�IU�)��G
��t#�q9j��:[�s���4	~ˀ\�Y���:f��]7^7Zgc���Ϊ�.~6�����\4��#�ǵi�9����
_�>
 ��� 9󛸛�cO��.�[K68X�����*�IH��0'�a1E����Or܀"�[�s�����`g���%��C�0	��Ÿ6�c�q� ��xF���m������o�����g)�zY0�UI��h�U�K�hX�� H���<6{����=�Z���;1��"ׄ)4���d�6,)*�iz�R<f+L}���/�[���O�.����L���j-F�2����ɶ �૯�z_��! yGi{2��$+�*�ѺsDz\?Z�*���K0N��Pm!@�/��ԦA؁NǙ�r��k9
Q��uQ ��Z�7X��r5(b] .�H�����ڽ��$���a��FE����g����� ��򕜚�
p.�j�'�V�G=/�˪�a����?���_�?�J��q詂2euܣ�4�Z���Kyρ0�2�>�k��Y�{��v�[�6�26��ƨ��IY���;{&-2���h�d��B�5f*��n�(UO����8����n���A���qt��o�v��p:7���1����n���55I�}k� K��|�M�V@��%��H#�y8�B��a6��4���%m�L�L��Y:2�h*������0�ը=�
�Q{+�� �xҚ%Ժݸ�u��9�2kmV��G��-x��.?�@���"k�;[�N��e������S���U˞E��%lX3W4;�@����rzV�Q��]�V�E��k^0M�e}���8'�F���(.�W�)c����V�l���6���6���Ns5�%��Ε�^@�^�?�/�Ƌڒw\���˻&2���@
�٘4�ҰhR;���6]!�d���'�����λ��ڿ�7�Ғ��dI}�>
`BoA
���@����2���P���9f@.�|�@���M�	��Hu���2�Ƚ>�&�h�)���G���ba�@�~Y�����F����m���j�O�P܍�[��"�X�5ew���-��jϮ�Ͽ�vj���G`�I�劎:{Q,O����坹���=�-��,���1�g����2"�W� ��HS{��}���qC�Zfr��Q���ǩ��r�es�U,Nk�\�����lv��B��敾� =�Jt�����.���vk��l�����?3��T�B�&��raa������|o�����`�;ծ�L�v��\��6�	�T3�$Ч%��R�dO�9Q̄��~�֩-���l�/��Bm:Fȥ�L��5�y4��#����� ��b<�AԚYṾ���-���b:z=�nW@(����4���[�p�
�(x�zk�<O��!�~sEfUV$H��*����4W�� !�C��Q}^�͕jQ6�3�xi��̌�́��u��ll@��[P�{$O=�<3@��M�m��a�oϵ]=5��L�E�ߺ�@�~E�h~8������ H3�J�Z`��[� ="��`�E�Y80f�Ė3�ٮ�\U���|ULx[Ø�$��d\����F�a~���"�*z�o�5E�^����0��F�O�^�u�Su�֝1��k�U�4��Y��r�C���5c�1��z\cꇅ��߼^-�;��@&�n�� �)[s�:��� \(��s�5Q���/
.~V+~fL�P��3����V޼<��WA�:Y����lf���.1����JM#�5��em�����?�����U�RPSk�qm��B�~x>�:#�2?���]�`�x��9]}���c`���P,Yw@���
��Ǣ��A�ȠM�@�W% �r
�<���o�����V������keA�kکNBSֵ~��a�=�Yh�:}�y��>�S��H�g��R�<�s�j�^�[��Ї|�]`N�c�z�b�b�^w~���0P��l�o�\~rL���b;�����7[բ���v���4LL�^�6�Gm+���^yk>jl8
�����l�3p[۳5Pm��`!A�@�6����˛�{�Z���h��zm[Pw��#�#��+ N�\U HqNgs\��ڀ����e=�wS��-5��������Q�/�w�_�{�U^�S��k͒�!� "T:�3!��Lf Zh %�:�T��A�>./��O��Rv\�q�Fd�Z<���边/��b;�7?Ƽ��s��~5-xOT-z1L,�u�v~�j _�-��0�Vh����N�W�S4�iN���_��2�l\/^ьiPS���\)�.�i@4pG�UԬ�x#��ZǲX��)�~�M��j.;�Ց�~k�qݺ_�	"���[�rf�f��,�Ԫ�:m
P��#q��A[��|'���&.y k��-���@X�f����3����u��h���~��תiZ��m ��4 ?zYFA�T�/|n݈ ����~�̎��V�lArfP.t�FQRո�����ŕ� �D$0����~2}ւ/� <X>7�О^�6��1(4��LOz�:L��m�ݶ%)j�q)X03�����.���?Ƅ������cy����c����D�`�;f��a������Te>Tir ��ģ�K��L�:�
��odQ�7��l���6��je�$�^����'�S�x�nd�Q��sx-��������m`�|��Zh��zz��~��5$t�]}^��{+e�>��[�mx��;�MѪBH�}��%P95-� ؝��ȕ"͜ ٬��w�M����+D}_���E�@��\[���Sv��
�!�̲;�y�|�uKX�4��=�*5gMm�/�!	�"^�&X������پ=��K�9
ׁpfqQj�t��,�y��謽8X�<���_mi���Ѻ���%�{
3=�hS~����uL��k���>K� �����-G�y�L��tC�n1�+����V\UP �=���KH4��kP���[4���uO�+MJ@n�����^G��u��*x_��p�9�}��s���#�D�d0�VDYJ0	��B����Ӛ1��_Ѻ�ٝ(@��\�nw�h)�zw;�J�>�Z�<�H-bjʄ{W���u����a��;�<G;�UӴ.�}��,m���B�yr.4MC؜%�#ȌUQ0���gT~����NH_[��E���|�* �g��G1GjJ����hv��-���Qh��$�I�y���wuOn���g�U��qh\�ʒ�(( w%����7}���/���-Qt,�{���4$�m�x�����R�d�U%0��I{�5���L����JQ���fp����/��W ��7�H	ȭ��T���}�t�h�z-�G-:����0+���*��ֹ��泥���p��W۵*~�W&��m0�W�vLpb�s�9� �tgƬ�+�IH��ha�{�;5M�)[A�i����Η%EZ�[@�',uO!��v��IxY#��,΍ܼ^&l���tm�2�u��Zk��j�#��u�.s�Zr\�h*�A����	Ы����9���Z/�(`԰�0�"��Gf%tn\�LBn��j�T��0�Ɣv�?�j.���}mӚ�E���#�vM��T�`�P{h�������G:�5��-3Y#�e~S�kT[��I�A?Eip�%��<
�vm��u[^cZ�r����o;�C���V|5���Ľ.�����g5��Y�
yE!X����.o�#����p%,I��GcEyd���R��q�� ��d쀂���� 'p�IXc�u�x]���3�DW�f߹�Ⓗ���c?g��6+�z4�����=Ξ�������<�,K,%�b	��h���&�� �	�0>��H���9���S �G����M"����/v3zi33'K���[�y�.�U.���p+*E�����-|����6�-QG ��Jtg��T�t��E�Y[�zIJ�|0��C@,-���^�4b}v0�օփ��k�LP]�t&	�>k�~k�j�ך	�4F��o�v�h.���i�B -��؏�ng�+O[��3�#�&*�>�/���5�gS	\	[*�#���8���c�9��[o��U���q`뱞[�:k���5.��6���{C�f�f��^�B�t_Y꬝��F{��������x�Ɗp��w�-P�����W����c�͗}`��;6A����N<�֯�:ͷ�]��9�A�����vd/|ny �E��^��̧��#z��.L�Z���^JQCb�-L}�[J��5�Wɜ�y鍊L�tN�R�-K�L�?�R_�U~X1u�"3��;�'�Sk��%ל�$3�qĴ�M�^QX��k_y4�Kk��=jR�j�G���m�=�m4�p!�FKZy~��P~f`^��G�I��3�+CV�*_��x��g�=鬳�Z���.:��Z𨯶t�7SҘ9�G .���D'�f����^�|沒��袛ݒ�=OT�����jC�Y�:��	��4��OϹ\��T(P��%V�u��1���ʫ{8�B�������*�{�Y���O��'0��H���و5U/��k�s ����3�Ȍ|N�F����ɷ3��������%�>0��<�_I��Ŭg4- ��H��-��r��>�D/��~�I���h\�S(�0Eo22���'�q3�T�MsDf_��-�ڄ�����6����e0����ӎ`��q�sV-�ն5zߧ���g.l�pH��̄���c��>]�@Z��r,���K۔B���v�]s�5�������r�u%=������E�y,�#��ޢ�ֽ�Q�� �
�k\\�AtjWZ��a�|�i���ɴ�p7fZ�-�9M3�4���Pm���~�������y�]�E#�݃��U9���T��spb����2' 裵hb
�&o�q��'�Ma�qY�+�-j�q�A��Ǡ7����%솵~�-`���H�\Ҵ�zɣXe�{)�4�}ш9"�|t�����v�Rj�,4����Bs���E{`+ڵ�5�5��^����Q�%"Pf�Zm��;�M�Q3�}�V�i�`j�l@�����dM��5:3M�Ϧ��L�^1�t�o��2z���
i΀�k �s��l����$07O�f.��n�������-0�8��g�r���KtQ
�����s� � �Z��깊��z_h�΁~V��|�k�y���Aɩp�2��̹�=���AN�ڌ�j(U-��>�է���6ߓv*��f&3��ق4OgȞٚ���u��Pd8^l�&Ġ��^ͪ���G{�;�O/-n1
�j��S��E��?������~X�K��:
`����.�;
ӑ�{��vʎbh�� 119��UhD&z�T��S��9g�e�k��S3�i�i�}��M�^W�g��ڰך]g^�����]H�x��NF��@=��#������&0��ͺ�Z�8����?�y���B�?��G�K9o]4�¹~7X�.�h+�W)W���/���\j#�h)+�-0W��j��p�k�Qr�=��+�ѳ防�fs��M4��R4��C�ƀ~�����������1XG�?�؋>t�h���yU�hS�>�c '�!EM���΁<q������P���k��Һ��j}|�;a�[O&xĨ�B$�~
4�i�Ѫ�[j��) ���4��S���e�]��Y�hz�����u����jL	\q[��z1Hy�۲%�&�)SEit�{=��)Q�m��a� ����(`[�6��v�dT"���t�������i��x�W�A���:�}��k�ǈ}h����#�E_q�����=�.ˇ\)�fטh�2�k,T�U���H;�[��5E/m����.���*_B/�y�\|����1X�cE�cm>��-��-:צM�@���������qW����Z�
/�_B���V	���h���p�*���d�E^�`
k*��h�l�7�:,�.$U����7�Ƽ�Ќ[ڹM�ꋟWR>�ϱ���GT4[�V�̚�d�Oe���޳g�,�M�J�S�uS��J����02�ʇ5rG?�Z������}��)W���K��z�\��!�Z���?Gs���x�f�B_|4�������|�Sa�}7_qj��*YA8��iv*.�/���~ �^��CC�������beG��{��`��&�����M��lll���\�h�5��s��0n`WŒ�9�X@Î ]A�c���G[I-5�E? }s�97�(�@{���}�;5V]�'����/�"�UHX���K�*t�3�ƌ�ь��&�(Q��[^�t�[
}sn�Id"z'@������!0��]�C��s���ob�H�S��5�\��_JibWw_��\<DcM��L����q�dڢ��*^�t'3:��}t����w�����ڱ�(�υ���+j�33����nK��(x�I?Z�
��򄏙	��Ͳ��I����aM����O�O/����O>��+0�nA��ծ]f��(��-��5���.5$>�`��$~f��!�v�@��H��y��+�~{���l��Cu�ٹ�|o%��!�K!O��y�.>���B�j��� 6�����|���}R��D��P���q	�Pe����g�<nA������B3�h�17/j�DfP(�{��cG>^;���T���P�|uiHf$Z��5���5���rq?�?m�RcQ�M2��1U�2���̀\ں
�P$��*������Z��"*(Ӝv��4?� e�A�`g�>���P# z]�w,�=����P���h	(����9jy����	#1p��Pƀ�͵&c �L�p����~>�ģ�>zw
�\(�V/K��2�v��x�@Z&vi�6ǣqO���]��
�|��4�ظ��x��0*ѫ��|.&D����r�;��EM��9�7�O]r�W����T(��1ט�]��n�00�"�f��@������_�L�w�g�B{W��y�*t-�e$�/Đ�H�}�摲��c�P\�85)�Ny��<��"o�⫒\to_��~H�Y�vK�b�b�ꯅ-f"[_�M�e</N�y���O�OŬ�,��WsCE]�^{팡����;lƶ���i_�R��� +�hĹgyZ��7X
��h<ׂCa@�ǳ�`0�p�gր����4�?�?V
,�O���%`i��-����C=��Ac
ǜp��˹}u��m�ְ�G/���\8oN��0ߏ�T~��{�}`ފ��59��~��rQD���=�Q������|�nF�[ײ���q��ӎ�٩~�qkhѳ"<�p�G�߸��9�8�g~kG�������*��8�Jm�[$ؗpZ,1 G��Aрh�{Ayx�9J\�EZ"���������+����.w�Q/� ��Z���ū�Q^>�/W:����tϪ� &�����bl2��X�ʻ
 �!*�\/̫�����Iְ���L�
�ӵ��G���o��u�B���(x}^<Zx���\؇�Qc�`��}nEF�<�Ŀ�g�Z��ptT,�bt�hYۮ��:� �_�.{r�!Wɾ/ �E�7y�4]Cc%_����w�o{w�W>i��w?os��7���G�FM_	p��Ѹ��T,7wb���w���T�f�y�js��m�
������|m�pD:es߁���k�@n��V ��AU]���轪�	fPë���Z���%2���|m��D�ѩ#�,^�tJ��#d��5�_�ɖ n+|f�,��-�[H��4�4���؅�T�Q ���w��C�� Y��汢���j��I!��'�y#m�9�S���9[��������c��- fnw�ܶ�Y��`!"
��r_�l���}�}���`���������}�٧��m`����~����:m(����D��1�8J+���k\���?�`~؞{�y��-?��Žo���ϼ��Qr�`�k��6[dS��݁.MU�#�-y�=���K8���B�lT8X�́o�ߋ�uuV`��5�1\}(�����W���I ���^u�����#$�h������o��&��c-���EIM�禠fH��*sd�*�@?�I���^2%I��5��F��?AK����Y�fz͛�O���m1�Uj�K;xIsW��]Ƅ�)Z���2�\y������;���*H!!��{�"�l��:؆�c��f�ݱ��;b�]�4P���B�������+��%_Bʗ�����s�>��������μ�R�[��h���P�x��ì`�fUW� 
���~U���������0T��=����s�#��E]�������O��8�o}�㿹^yb�b�z�$��3����JR�H~���~���2������� ٭���M�9��C��[�L'��<S��]�׌_��*�᥾;Pz�U�F�h�ڞU����6�oʆ̻�����$�̤^�᫣�f��x�߳$$�ƨ�C�	&~�U���h�L��qWn3V��y����G��1���Җ��|_<�G�%.�?���vβKܨ�`}�~`�o��<������vB��뀡1WA��s��`L��h�[�- �����[Oi�Z�ì��-¹�;l��`�nW�M9��1L)�
E����� ��.u�+'���7vɈ��G&|���>���<`�U��t���)8V��89��3��2?��?�_�����~8���6]���*�Ҧ�2KY�)����<O3PB�BJQ��
^x'!�x��4"+��^�"t<m^��y��xgUB��D)^���.�;�K �_GZ	)[��5gYI&o��܀����9L�K�@7[�L�"H&���_$nw�|c��_�5�vv�J}����Nh&�_�.?EF�2�,e�3�x������s�\J��	-A�����^�癰��=��k�R;��������y��RϫU�e����♷��A@=�{���@���V�{�o��z��C�qs=�j�G�-oyK���&|��ߟx扗�Ћ!�,K�
���ìW������m�Z��������~��h�m��e������ٷ��e5n^���J�He�$6��.��%~��C��ݛc|131/�+�ቺ�%kG�&k�����%謹���ӷ�Y2z���))C(�|']�\�����a��'Z�	^[�¥xK�ђUO{� ꋤ�/1�}���K�o�����0�ᖛ�2��//��/��F׽n,=�c�޸�R&hhAw5s�W-!շL��kuo����*x�k<@[��as�Z���*d��
��Q]�B����~Z7_ 7����U�����h���)?�m�5*��2��p|?C#C{��9x�>��=��O|����>��O�Fh�e��n*j��"�k�+�|�P�N@�',W�0K斋.�j]�l����]2�cp��o�?���
�(� �I����[��t���g$�m��u�[��D ]�3��Gv-��+H�I�N�sh'	�Z���Y}�-�k3����m0��g�Ͻ�zDXl�r��75e�O�߾ʰZ�$��pY�*@���	�R��qd6�D�"p�#��S��\�	T��xZ�_�:�[�4�ݴ��,����Z�}�z�Vyu���ţ���,�=G�?�E�����w�U6/�Į��X7]0�+^�U��Ї>�y>�YAo��3ۖ��%-[�f�8k�O��MM�/��u�r�f߉��E�<Vkޗs=����ͱ�]���=c��g>�-S�t%Ƨ�~Z�+�I����!w3
S'�����y�?�f�vO(�s,t?��HT�}�m//�-1@��)!�M�~�N��X��{���J �f�<�Q�����x�����$�D�0��v�ʽ4�����VU��)|g9��4��,��r1��-��K�c-���ˀ�K�����t�Z��w��]��z<�.<[r�r�j���5��om��(�1�B�s������]��{\䉩�ް8h�5�P��$����O]hX�X9�л�|��Yǃ%���fZ܉��0O�ue�ɋĺ�Û����:�_�����l������X�+�i����ʁ���N!��N֪/7�0����Ҏ�7�X����뱢�^P@�Mj���|�(<V��Ĉxm'3�����"	�.+�k��(1�C�j�K!�a��EÍ<��~g�}���e�wg� ��--�9qa<���e�X�票�&dɾ �`Z2��[-�}��oıh��.���u�. �Ir;w����Z�Z�Z�����|Y|�Jr@a���׀e��_'����Xh �oQ�FѪ���D�ȵ�����k�u�QZ <@ÿ��#� ���9��c��g�X���
渳'�yGߺT*�b֚ۖ�r�q������{
�o���%/y��d�w��Ge�C=�5��i�g?���_7���}l�q���v���}�M�ÈY�,�-I��m�ح���Q���6ty[���T�7UA�w���!S/���1_\yBy_���ik杞���]i�`=_��N���)��	b[;B���0!� D��Z�Z4j��k�K� .=�*Kg�w����ŭr} }���D���2��K�Ӷ�;�aZ�n�<���V\����b������O���K,���d�h���*
������Я��L�ը@�ޯ<���O\��ꦮ�:���@��N���v�mV����cU�>���s���:A �������L�����?���v �0%�vd;�A9�򭡙��lqi�w�-%�}Ģ�կ~�9��Wn�f<W���k̃�+s-W�]���e��_.�w�>�����_��_�ڋ���:���X�T����	=��)T�|,v��%x/X>R�a65~�r| �v0C���xNP@6���w����(�KO2<�Ak��~601ֈ!Z\��0���`��Y�3�{=/�)� ��1�k�]���+S7��mAr���:������t5{��Ț�h�2�Vבh�w�a�u�� �jΏ~���ɮ� �ߴ��X�F��K8�(�ǫ�2@<q+�������v����G;�ߟ$�U�=��<��Ҡ��a5w�DY�x�#:�ݻ:�N"��YJ�mKWϩ�H2g��� �B�]����nB�/f�̳pϯf�m۹/�3�*c�Α9���|���y/�����'P0�u0{��SӧxO�����ܖQ�B�xLe�K�Pd(�=}`��Aᥫ������O�D�uP��u�dy݅ქ��}��� .� ���~f�nH�9n�t:�o���m����Wq�H�`�E���@����C��u��������A����"?��m��I3���G
�l<�}�_�[}j���9J�O �-uc�5Ku���F,����*s�\�9�������(3���n�+4&��fw�+���׻$-B�{gy�t���2P6���MX��?��0��~��ݛ��";~��|�+�G��Wb�k�c0p͏�6H��s�s`�}��~�4w/_X�^��yo���+��$(��tL�1�����W�  �CIDATc:6Q���R�����G���/|�V\M~���ͻ���l���r��v��Ȓ8�Z6�����'�beҷ���DQ�%�ٞg�4�B[��:n����G8��H�����3<��^��]�Dں.[���� �},�Gr�1�c�zfX�{��~v��k�>�食0�]h�G`��cA���]�)@��t�$~���������_t�u�W����qG+��-���X�*cq�W����-�� ��T�* �ky4�!���YA�z�=�I�}E }���5yP07���8l�������O�Q�_�r�\��20�5^�����=ѥnya(���/~��(g/el֋�D��27q.�:۶�?������g<��d2,������v�o�"=#�v�<����	�J�M��s7����:��r�+��)�s��	�����h/�k��^�׫�L8��w��ۉ��-m5@_�b�?�J2Z�Sc���k�"Ld���g�z��^w5
�7��ԧ^B}�`�Ŭ+SM:�=VB+ܛx�F���%c}6,�]�<ظ��h�Ս�5إ�4�� |ʕ4�>���p�mLa��}�x*�Y{!�p��1.��X�*�E���$���;��ݷ��Y��j�Z}��uΏG ��̋��OQL���( �	��g�^��I��&���pŀ ������
�=i�����4��˱
��|�5�g�gB)�������7��F�3�+1��<52�R���g9�i��á��ۓ+�'�sb�P�_���-��#�M��%� ^�ll�$��{z�mo���} 
�?Xv�9���$�ۆ���6Ź���M?�}l;�9	��A9{c�'�5޲`Y��^*�$Яb���ʇ� � �,Ѯ���̓���G�vj!�v�A����W3!`;):��N��s���c�Mf��q۬#3&v������]4�[H��)3O�r�b���a �}�oc�:?���OD����Iܓ��g�����S�����/�f)W7v�L@��T@�(����W�P��pH��+ }����Ir�2wOs-s�n��s���,t\���}��$�Ƃ7^����8��OsYn(gkr�!��B����� ����)�|!��'���'`t�Xh2^�Ai��Sb2^QNS/!Kt��ӄ;������em�~6J����ٴ�t\���7F�����at�c�&��m�9�b@QF����c�}�9ꨣ>C.�w%|l����5^�o��� ݎ��_��E�u�5C=��j��~��wrݿ  wv`���vhN6�c�n2!mnL}֑Kr�|�5���0�C��e�$3%�6��L�ڿ��Y����v ��K��U�����(Xr �����7�o'G��2��g�j)����=X�х���p�X���ў��}�;����[����0T��~��n�̀}���Q�R�s�������oYJ�ڞ��/ϳH[�����&���i�]�0_��iOg��70[D�s]�ʓ(�m���x�p�n�N�EI]������o��I�;J`�Ю���\�X���L��R�c�0��������7��~��>�1+��鞯����&d��ȁ�v;����͌�Gȿ�caxz�_�T�8��X��3(O��V'��#M�	:�M��6t��^���n�h�NF��K�6'�L��o00�t��O�����:��d�T���D����ݕ�l����&�+a�o��[���z��[=��<wo�i/�!�X&`բ�5-�f����y�\s�����꺯�6���o_Q��:������rϚ#ӷ��wWʕ�v��n\2ݝ��I��|������aY��=A�6��X,��z�up����!�jK���ر��$X��\�7�)Z����ל�����#�y�xSm/
Y���,K̸�_@��T��T��|H�^��HJ|�{cvk�=x�z��E?�����?�
]U(a�u��gc�}���
�,�|��� �l�pི ����ӄ�d��X��՜�h�]�(x$i�s�ԑ	�`ߏ%(�6O@'�i4��u�&K9�)��&
������H��Ҧk���S �����ӟ�<A���v,�z�DM�
of�R��/�[�iCP��*	I2���m7�%�n�;�����Ô�aJF���#��}�J�t�cil&���J��=B?^�$�%�5�ƒ��gd�߄��9a�w�������8����� �+a�q�Z��ر��E���� 󷲣�����ϕ �4��z6* WϘ����Y���lډ��}�L��!�2�ǃ����V*��5r[���$��\,���K7s������F{?�_t=Y�����1��I.+���%kp�X��/�4_A�I+�;x�0ކU��vB�M׌Wvc\x�@K;���	4�����X�����˚�ꎲ ��.�[t��ZZ��ó��8��?��?�E�m	m��X� ��gb�
�+G��A6M^0�&ˆ͌:��w=����o����w�׶�e�g�~��Ґ~�8yΏ �K۶=�ߺ�u�����cuE���+5ޑ�y���ϣ&ĵ�w(�����5��L���X��J"���$��<{��͞=��L�����n��^Ƚ)��F��T�%�=c�Vwx.|�����Q*�^��(�k�Ӈ��^̳r^�Q��q������&�d��L�w�����7��~KЙS�Uu��0h�s	��bN=LQ��T��f
��H�-g�%#�Ʒ�*'�$�39nhV�ր���m<U�¤�(��. �����]����v�ԬM�M����i��BC(L�(���,�̲�$ae%��[]�պQ@&�9�1����G=�;��N��d)UW��o�����w`���]��ʪ�v�� {�뒥�7n�(:q�۾�	ia�\�<�zL�9�p���h&<��ynY������0߈��WRy!rhFA�\�ob��7���`�.�~����}<��B��e�Ȼ��
���{噾���Ǜ9�_��X�wr�V�����=���7��~�;�zl3_�rw,5朻Iꋧ���lp'���)�\��[��|�YO>�I�i�L�	XI�R*�9(
�0J4龠HU.�k&�RQPΖ�4�l����h��R�'0�ۨ ؇h���EPɀ��N�>�.J�������7�OFrۓ�������cM$	(Kt�5�`�=ٺ����>�m��N>W4AK�H��F"�2�2x'PG���;+8��o l��2��p��>�s�}�¼ҢEڔf�[Rτ�W�"�y��3�T%��q�绰̏�k���I巹��l�7�����y+������qIm��A֙�I�����]�5��Q�=��F��mVkD.��y2JfdvUЪ2Y?ې{̯̵����ᛪb����Xs(�C��i�c������Y:-/m}2k���٬50�u�?��E�~�T��"t�`��U'S� ��Y�T�ۈk������˽��k�e+$�mA2�0��$�E�L2TL�Y����g�>Q�`�轿+ޖn� ���>�1�����_������p�sJX��Y��Q�ǊX���W��eø��%(���n��h��'�wc�ۉ�v���n��$�Vz��Yc���rղ��*��>/,���~�u�<�:�s��I��y�	ui���(A��7na,�����D�w��5�9yس���×�����O8V���E�z����M��e~9��ģ��o26#%��^��:��
"m+�V �'R�Y�a}�+���Y�9I��ܮ
��Ԡ�����\������6����İ�R�g���e	���ӕɍڛ��w�.W�,U@hWa@�h�0I:�nG�W:��In4����;`��5cIgr*\����غֺL�k^&�i��}�b.0���@���YFJ�*�c�a���3��O���n
X�	�<�E_��շ<���
��K���q���KrMw�� V�9�I{� .�u˚N�}
浸z���	��;x�����mb'���mUI������ϝŮ�*��*@+�����C�j��+�Y�}~��{����Q|��	&��|�bzV��֨H^C��6Ʉ����&4�8�Ɔ�x����(L�F�{r%�E�`�
p��������	�ϰ��rW����sc��߮�9��TEp���z����bY=���w��a\�Ak��L�^�Г�Q��xϔ�Y��{�>�����o���@�Of�N��&�:�`��F�M0Q.��{:��ҵ0C�'�7��&��08Qu�	�
H�����O@K?��:�}X�܄���W\5��S����q��k�>��Ϣ��� �c��Y�n�HL�1���V�bWM��#JZ �~%���Uq���e,���x-<r!���d���e@/�B�\Bi�=�<���i(�7a��L��	���/:���NM�	�t5��OzW��Xz�Q�0��>@<?����f~�_����?�ֹ`��x���5�d�'䖱�xx�5ɰ'C��	[|����xa�?�����
�'8�q���#������eg�f�&7��ڗ��V�7�̓�����
��T@�&���̌a���)��r����e5�-̥a�~ }5JȺ^�%UQ����Y	�m�	�c*26?����K�B���%-!���*���D��%5(�0c�2E2�c��=�w�E0D�Ta`]c�K��A�Na@�a���s��q�����|��U��/�]��VHf�2 �9�����}�V��7l�ؕ��*W����9y)��
��_-�_�;�y#��,�Sq�F|�x@�b���$\�JBL�x9}%,�f��0�9-tJVNx����Y麣�+4�L�ꉲQo<�U�(G���N�Cb���I��X*�eEK��U���wD�[�0�݁�v${���oGC��C>��O���o}�C�������yvM�=�r'��(��'��G�`~�X�����l�7��OJ��Q��0h#3���}��/��|�r�K���{����eγQ�.f��_�}�<Xs\��;v���w3xf�(ޝ�����*�C�!�D'��p�QS֪vRQ'��%�t�[���x��&>Dx�I2�2H�G�Y`׭�R!2�wŚ{2IR�`i_@l��o-�h���%VM��OG٘k}�r���1 �I(\�3N�0n;�J��t�eC,�u�$	�D8U�1��*��k\<
aV
x�b�NG�� �;x��'<�	�Q�xL��/«p4}�������RI7r��M�����.���Ё{�g~7�[)������0wk�~hW~�⺤)
����r���+ p.jU3���c��{X_~������]�����~����ܚ�ۀ����FAo���R���I����܂�DC.N���^�����1��!��D��9e�P�E��h��.q�kx�@��͜��1��c<�v�T�遲%��?��o�,KǗ*�3�+B`�cb���8��1ƹ�J�:�kݒ4'��}9�d��o_�<L���
]�hha��X��k�b/,�uRԣZ
��$�@Z�Xd3���^��GeM93ӷ|����xj<�k= |&媉����[B3����X�#�>�3��"�3) s!V��	���\�SH�Y�]����L�����?ї��#k-��'JB7�*;�q��)�,���n�:��r�W+g~<����7�	Wk.`+��4��=�W�=�{� ��s^�����i�`hR*�d.��P�ތ�xPM�����\����.o �"o>��{�t�ױFޮ���:��e�TV��^���(�#a�g�]�\�&����A�b����xw"�#���-U����}�'Yڸ�$8.U@�Qh	ں��ҵ\\Fb��2-�2��q�q"F@��k��V��*� �M��#y�I�ZG��q�v4.�Č��`������;�' ��� .щ(X�a�����?��Ό����2���%#=�Aުq׀C��c��P#$h�*����D���%T���r>occ�{������(�D�x�ϣ%�W��;gW�	�*؅��.�\�a�
�ӷ��c�p�f䚾�0�̈́����ҕ�s�~�5��ˎ쏲�%i��	̿����OHP*�)��g>�������ǳ�:W�d#��y��������ǒ��0,w	p�x��2СK2��.�3�P�<+�D1���є����+��?�s2(�Q��%u	sg��x@�*�ݾj�%���?7�C��s�X��x?o��`��� Hl-o--]�îpK\]��z1�h�;�[7c����,��AЇ���ֲ�,`�U����z�(ew"�E[��E��xIֶv>c� �?V뮌��L��y��^�� JM�I[<7Ս�����|���Uh���b��N��	�����v	�E����������*�.�4�;j�w�DM�rϖ�q?Wwvق����}�ZZ����\Z�9���%O9�I����J�k5�a�D��6��������	l�1�I0������b�?zmn?�G�2�:���J�6e���S��[���W�|7pZDS`�7����Z5�px)2�zW2#C��]_)�DI�+���5���e~��kF#!ҙ��9����O�<�M�"<�g�(z�a,n� }�|;�n�Hh'�nw�ԌS���>u�ղ|��st�	�
@�WWy\-}�I\%	6&$���W�r�f���昉�u�������y�f�y���XȚ���'̱�{�󞇡�m�p݀���U{w��&�ld�&�����5	���+��f��=�p����O��IF�bg��(����_QJW���!�Y�"y[��B�Y��Y-�������}��p���Q-2�+y盯��3懲>�mK:8�,�U��}�����y�s�Q�5L���|e�/|�o����NkEy���k6�Qf��7@�W��7Q���o}�[���6u;�m�M�'�U@�0��Jf����S嫾U]b�s{�
�(\3Y�y��@�U�xV�4c�=��{���lc̵ے|�x��{'����צ�s0�΢�y����#K�B��Vͺ3.	o���n-�w�csF8	q�u�h�浨ո�����a�$De����X�
 ��nO�[��>�\�	0M!��6c����]>�1]Z��{���ߙ����6�H����jL���F��q����$���",��GY� ����: ���������.g�K��W��y(�^��������_w��]��m�$y0
H r��5�`>��uNU ���5Q�3�Su�ץP	g���O	V���0�?��'?��$	�:6$�=���w�o��G&��WR��=y(E��+#���Ǣ������c�B�����T�a�:�5���Y�*��n�ʫ�[U0�b�.Y�m+�<ZWqʓPg;��^�O
��@��B��ET)�Yt'�W�٩<�]p��=;O�w���)����/U@g n�-��Ī�������:����~�u��ƾ�š��;�w��!���8{u5��W�lϺ.L��ov����X�r.� �+��r�\�0�������8
�:(C����|���j����{�h�Q�⒫����eIY $�xkCU$�1>��v q"��~���4��*�%-1�����$o�*��БGS�TKR^�RE(�����z_���?�R�B�*E�^ǥ��v<^?��i#������̧�yf<�MP���|([�BfUj�?��z��v��1�d6�
����٦v�,u`�;������/����5BS���*��g�������ވ��y���G��q���k�c73n���y3��ݘMyR((��g��'d�x���L\3��nW1h�����C����������Q����ǯ�
��E���!��w���UL�ݘZ���R~���;َ��]�]�n5]��ZOL�Z���Dq�łS����V&ܷ���t�3p����$0M��e ŵX��o�xB�ӡ���4~o�?������L�ՠ� ��X�%֏�V�q<�'Ge��f\��V�|�1�m�
@�<��㰈�[�x�J��ǅ�����?���?�Y~�0�J��0���A����
���1L����@_�:f�����"��q�g.;��XF�����cQ;�S�3��J�����/��U�6$��@v�{��F�ŝYz%f�4���H��)9o~�K_�բ�/� �UݔE�d.���a<5������(p����N�d�<�}o&�r�ƃ�ح(l��[�M�\�������<_���J���r�6@�=������i�^Xb�0�Rt;D�-L�h�KwM��������s�t��jO�����TPF;O,���2�I�$,V����G;\�Ԏֆ�����J�L�tbq� 0��}=���0j���>OF]��'B�L�i�tU dU�{ޫ1����;���+�׶d$
���n��*�3^�_ǸZ�~/Z�\ED�9'.��O�n�Ou�	��Ō�9X_ǐM�+��ȍ��%�|[�����7��t��D�?F����R��*��N���旪|ź�P���o,9��/��/���Ix���7|&��9�W<^�G���?�q�5�����S���kY�z���c
b�r�*B�ȵ漯뛱�~�ʂ�����EM�e�=�
���5�"����o9'
tU(��vj|�o����^�k6�C�$V�^�u���8n��ɟ��l����CP�*��Q`����1��%��&�F�В��e��6�k��V]�Nn�A�Jw)�1	r���. ��54Z؞맓\K?��0_��$uYM���
�M�͍���0׮��?�,�q��0ō��܈�2����?f���L޳�~����6ι�g�0��~�µ��.\��q�p&�D'+4���nI8	Z�B_W���
@��6�d����n���<�4>��l��*4Z%���w&���>Յ���U����C��3Y"P�%��s�V�#����S�+���K�
,����⚤T'\�L�GB���'b,fDь=���_}ָ�g���%Է����[�aW���E@��1�)�_�<��s�<�ۍ��xOޅ�����
����ͪ�'A��l��ȳ���Tv$g��P�˲�w<�iO[�:B��~�sY1��A���
�u��>W������+��(�[J��]ya.e���}և���������K[0��܉Q��ӯ*�*���9/�o[���>7�ٙ��]���h�$�!<�2����1�Ii�fƻ�+����T+/�	sO}�S'���RhS�P�dj[��cm&�^-�X(�1�����\=KcL�sY���3��ush�6�V��㶀|�=0����5��سy�����DB����u� ܓy�L���;���V�r�A�5��St>'s��W��Oe�]����R��8"���N�$u<l#�*��Q�UP�*,�>V\q����ү@@��w���_�/��/�r�cB4+�m��,�{�=\6S��4���E��#Y��q��9�i؜��J�0U�6c%�ZR�^��
@��c�XEE:a�xTº�y_�<�&��/zы�i1#��$f�>\�����lGY�P���}S��s��;�}��Ǐ<�Ol��dB�)���@�XF>����0��h�����Ivo�G ��ȿ뽆͊6���+ɑ�'d�x	�[s�mN��������/[ү��$U����tr�,l�S<�C���m�Z� �L��ceEXG88�V�sI+i%�*`zN^�c8��c�x����	l�Е��^2��>qI�(����UR�
0jq��=?1Ĵ3 �I�y�!� ~O�����p�*����RpW��V���of�JZ��w�t����5��`W��j�Q�B�juU7k���+����g���Uy���o���ݹ$K�	+��X��4u-ռ�@�4'���d�ߟ�A�q9
���ː�sx%�z�X��1�M�R�S{2&�2�?o��`�Җ{E���mG��m����%~e/�[���fS������7K�~A!�Q�Q�Y������	w�o��Ҡe.���.�%�FZ�?`~��	,�Cx�[~YҼ�7nShԭA���3�J��c��;<��
��� �p�2��_�&;W��^��J�`�5�*
~�=��O�˽�L�R[eV���T����^�mI�]�v��R��
��B:�=�}t�*B�#r�#4ʀO��ظ��\�o<�r��� �N����x߭a��w2i���x�m#V|����;��
�\�>���+U�k�N�(3}��2����}� �6�Y;\A�j����s�Ϫt��<W�$��H�f��A7�%h�g�O�[�U��r�+_����e$��V8������}�Y�����������E�"��B�4�<�����ơi孾�^��/�2�" �^7�O���~��1��3�sY�	����{Y�}�FF�2vA�+�y$�� ��y��40o&�����VVvLTq� 8�u��e5��Ÿ�v{Ab�+�1��[�?_3V�j�L��^W%2�>��$����Y�
93�2���S��u5ҢhD�2c�2Q�?�.��s&��?�5�u���9���ӻQ�Q���f��:�9���E^�F��Ij��R���!ݓ'�tRW2V7���3E;s�W�p���vUx%�.�:�l�~f���k: &�@PV��th[����s#���{�) ^�q�	(i+�����*#�Gt��_��> ?˱,����ul~2n�	+��S�4���G��g�z ��Ec<'�c�A��e�*d��(e�I0��N��V���X-� zf��y�)�Ԍy�5�y��e�H���/��X�_"��sl;O�� �bބR�$ڙ&Mj�!I��0ʼ�4����I�|�+_��?4�� �j��Mb�h�3��>p�/��&cj{9���C�آa�Pw'��Pv��^_�vR�m4��ܩ�0��y�U%����130:��v�q��qi[�!�n�<��0��Z|��Q�{�:�d��m��\�Z�����ս�@���T�@��TF�����a� z�+�G(fU��6r��Np���0e�n�xi;"`R'B��X���"�~�D�ڪ�G+NLn���i�����Ō�)�1x�AV�,���������gu�Q� @����~�: ��������o�ȫ@�2E�󭳀k�{�0L ��[��j�9Unڏ�X�yM���s��@�k=�dQLr����>ت���?�e����j5I�b�C9d_���	�g�T�U/��8�o>�o�V?cO�7��Y3���5�AGv���94��V�P�}�����򯞧�%?��g���N�檀��Ȼ��s���\���'%d�q��b1o�����Ƹ��,U@7�A13 Z��jT>&�1�/���.��YJ@�Z?�k6�s�Z�4��c
D��N�� o?byN���xa����cU��X涯�RS�[k�(���8@��F��4�O�0qe��0�	2��LȪ�T�;��x3�Ws�|����x�����x	m�#t���&EMV"Wc�g�?�ܮ����ŀ`����W����H[��$O�Gwi��Y%0'P�j�r����tE���Z3����OQ�tī'*<��K�qNiE3�b����'���矅;uT�d���?��?�p�Kho��.vc���(�%-c�/�\Ox����b󣖊]�{~���
��e̫28,�R��"_�M�om�o���m�p�z�|�X��U���*c���Teb�E��yI���u�� geK��58w\�ї*��-H��"��_���վ!�ad���������j���EQP()��f��d�1u�]����_�_�ˣ
�0B <1�ξ��������/%M�o�o�ĩ@Z��y���Ӱ�db�"�sTK�>C��"�����y_�/v#�������B�����b�2��R�ڼ��>�	�|�%<�F�x����&�Z�>�W ��_��\���0����pUO`�VW�����K�x���#��VLd��,E��W�@�/��݉�j��9��;����O>�Y��!�<��s��'>�wc�=��b�*�zӲC�pD�z��_}�ǈ��L�y�/���S3���T�<L�/"�"g*OE���~UNнwr��,��,��c�TŴoyW9&�����Q�y>�-{��x{7�{�V�Q����9�	>-�
�Jp,׫��ϣ(��z衷q�k8�Z-������$���8u��u�η�l,s-d�0�5/�f鋃N?O�zk[p����&��o_3����o��[�!c9�D8�x����  r,2$�!��x&�@�����+�Å�������"ȯ�Z���'=�e�G�̮pS(j��'��Udr� l*O�>
�w����x"����8E�jy"8nD� 0�����/���M-��}�{�)��I �	d�O���4�t��P�^�{ƶ�W"̪R��3�_u��5��O�}P��*x�'d���/���Z[NaU��>�g| �W�� ��G\�*E*�h���y��3H��^��S`�n��,�r��[{:t�67��9�9����6����J�Ȫ�0�wB��(l����NՀ�@�Temέr����xF�:7�x�"�i{]�p[p�i�q����.A����.٥Xu[:Hh�SyOd�^A��g���:�����0d,�T��U`3�.Pk��Ll�vd.<��$��#h/d���"4���!�5�O;�܏�mD��X��r�މ}O�3[��@�a�$�i�Lu��x{��j��I�I���5m�1�9\��aܮ�W�>�ԟ��P��$�4���r#L�lF��Yvv ��nLtZL�Xrr
��LO!a�<J�<fq!@�X�?���/�2��"? ��f�r�W��(�ѭܠ�YW���X�׭�p�f�1����Q�*�d��h�9䛸���H^���|�aϕ*� �]\�7��������ZǎW��m}��u���$���4&��]�"�;WSG���o�dI�y���O���T!uS��J��(��WeqX���m��>��"N�z ���LwR����*"�s�������,�����Hb�J�}��aud�������ڥ��(��� |"4%8�w-�X�a�����?���򗿴�\��Y�&��.���lK��0�Zwm�	sn��w��肾m
�&�zŽ�$�yǼ���=������;dϻ��T>W!ib=�؎�w�)�Ԥ��W�����5�S��b�e$��?����]Gq�E��N�
,�fw��5΍w[��&�7 ��"�/`�Nt��/w?o\R7�]ʖY������a�ޏ�z�Dy�G��6 <#��3n*yɄ� 0�EA�+BM�K�.h{6��%ɀ_����UlT�#��<�{�Iq���� ��+]�nx,�.�>�+|P�����o~FQ���o����Ŗs���W&���^��S����d�|� �n+L�-]r�9���<��`-�x-�ca����%,��v�s�«S���,rF~����b�Te�Z��C^�gϜ���A1�6s�
�R/���ク�\��a���LQ4r�~;}o����aۙ��"��+�Q���d\�Q�s�:�&�5�0�:~�A��+����<�"�K|����gT���Uk�w�Aʧ�YIN׻Ę�}0Ʈ�]!bL}�G�d��t��el�9�W0S�X]�u
�#9��NE�Z}2��*����ڌ�����H�������Vl��{e��q�|[�rE>;Ņ�V</?;�{���6e�Nα��߳	���z��<�-\wϥ�}�IK�/�<�[����(4nex����+ஓ�p}��6'k_��-�b|֯�\Q���.�$�*��eGa��E������5�Y����eW+�����\�K��̵S�?��X�;�E:%T�\k]/S�'U�ν3�PM�Q�g <s2 ��eURb����D��'Y��}��w��Fy����������8�Ei�(ZD�`)�"�{�k��>({1޲/����}��׎�M�`���J8-�<�+c^�`\�1"���W��� ���k�v@��/���7ᣓPRw`�� �e�d�@V%!�D��k�P�*�à�^����U�84�AK�ז:����vǲ*<��R�b=��8��7݋�/�o¢����*!s}��=��9��y�J��[��oR��"�W�6����bݷ���s	i~o?�\`2mOAi�xLD`���(|N�W�ߖe�C[��r��vu=����o~�w4��ֺ�$�� �&����R�[,���{��X@wZ;�V>o�M�{ܖ5\���� ���q?����~shݭ��K���y&^�
�4��I���⾡�yX�@h}>9�5�Cye�Nj��������9���JW_�m?;%Ծ��ɄO������sT/U܋ì�X'�z}�2�.Y�6X�y������mo��������I(|Ʉ����%�u���gb����$��G��Ei���'|.5
/l�ȝ�(��DA��(��G<O��y9��G���d��s���ci7�o[����Y�}�s/c��i���SF�p�%#�+�������ԾE������j��g>&��X)�U�^����I>�B3ڑ6~[������zJB΁�O�:�Ӯ*��hd�0��v-v����S�Kk����l�q'E�?�U����3\�Z�˭�;_,�p�M�_�1�el?A%j3�|�$x9�InG��+=I`5^-�� � �o׵/�E�E���G?���]���n���E�ux��;����r�[��RLWk���u�W!��
j�U��9�߄�<���c�H��7�������ʿA}��� Z@��I��sl��o~�	������� n�\�<�Lښ���ӷ��1hx��/q���<i)��rqK�)�A��A���!��=���U�w��V��-Mx0
qQo�u���9x7���N�󚄽ҷ�bQ�����w�a�{������5��u���rW��n����s���L���8ӣ!UM+�� C���⊜k�y��g�2}=�W/c�佮m��W�,�e,�0C�.�P�h��vW�(p�|7�n�x�_A������c���w1�q�mK�3ġ��|��� �͘>��*��/��jvz���.�TO�Lu?W�� �F��υw�ěs( }:���(�����x]�(��;+���>ʻX�]^H��OI���<s�Z�Z-���2���j6���,�E�ޟ(3�fS����O,���/�F���Wzj��x?�Ӣ�zO��kQ���B�A�h��۞����N�̃5��:m��;<��>(Vp����^1���/J�y; z'K��+�G�sF��w�Iȇ��+�7I�̵҅9�2��]1
&aȍ��;K�%��A���a�$"�Hq�mK֒�ಹ �vX�{!8�����A�zL�`�[Qk�W��d��a�f�зIr����؍Y"��g�_�"q=�3K��ۉ֮�w�&1�0N�h�F���7�1�����d����q�o����y�&���o����Sh~A���<������G�)nu���,*C��qc�Z���ٝ������{��?c!�e&VZ��� �5��Y̯����%<d�k�klH�|��C�]"�u�ۖ^��3��ٷ<u���{�x&��������;�o\�<[��,� V�<��_ �^�>@���}�OUy������ 0��'n�}���ȱ��6����i2�+�s�GY��=lt��r�oZ����lO�%����5�����p��p��V�>�C�Or} }=��1l`p����6���)��6���0�����(��+�&NW����i�]pX۳>��XLO����<�`U-7K�Ƴ�#�m���z��`�숰Z��ސ�d��c�&>����5���}K5�P�R�>���/@����7�q���E��6<u4|�֞�ea�l¯���M�[7�^7���Nv�c>����W,4ȹq�J3s.��H��?�����h���i���]�ڃ�xޅ�@�5�`�U���.N�j
�xP�o̏ D�.�d^�%i�`B��61w��E>����am��L�/
t@5
pdq��w����?��~5�ܥ٘E�	H���[����i��~}��3U9�2��pO�T�s�l��[`�z���]ofu�m%l\�I:D�%F��Լx�Moz�iX�"�_`����μ'��ZW����Xc�U�|V&R 11�E�}��H
c\D�����CV�)$���M5u�8ξ��r�k�W��v� �H�z8|�`@@�^����Lt'`2d3���_��X���TK<�'�CK|���x���0��гH���v����� r<�	0���0�-E��8�A.�Ya1���Ҁ|�9�}��~����P���?����|����[x�6����my1�sC��u��VN��lun����S1᙮`}E���žh�2 �-�݅9��3�t�w0�M͵�1���jy~^���U���jx�3�P��r�g�θܳ:��ԇ��3�+�W`O?r���(5ʄ,���xp���v����#`\X踩od��_ �cI�"Ϡe�!�$���;�%<�\CE9��O������Uh~��I7Vpx���n�<�A~�xc>��ʰ[��=�f'��@&�L��L&ȅ�czK`^�3_A��"��v���֨ 6 _0ۈI�w�����f�^��1�q��B���$��[IrK�W�-O �����In�PD/D��~P=�L�Ś�
�]O����:(6{
�.[3A�el��Ef��}��dx8@A^�㉈p�\��v�r�C��������d���+6�����l�*\��p]WR�H��$�E�J{b����J���}�%i?�#�Lm�3~f���;����W@�xųS-�|�\��n���r��P��hV�?W��J�	'�A�������ӒЙGհ��z��0�"ǫw F@���ȟ1(#��fƹ?Oc=. ]�`���5��ubE���N,�Ɏ�mݍ��	�!����������&�^Π�ő��Z]��F�G��]�}w0V�QW��-y��`Y�1�kh�R��)p�߰�OA���{ ���®G;��G�ŗY�x`Vg|WG!� ߉��G�n��Ѕ�N�G�T�`�^'���1����;�ߙ�ȫ%L� Z`7�?P(�5�⺗ rK,!��'P��=�����N�⻸�k�rw_���3/WUJ}�����:�]���~V�Ϩ��qJ��N��Qْ��;R$楌ٓi{�(��`�FQR��yo�`�tK�������#KT��aq=3V�4W�T+��G��G��W"��$V�m�w,� om�̹9��\���s��z����(o�_k��s> ]y������*�^����r��B��`{��tBA��07��]��s�L���*��D�	�m7���פ��5JL�����Kn���� '�0��.C�Ð�
���z���^!�+���u:��c���>tv�������P���x1�?���7��bY�{�s��f�bnkϿ: �����xwz�;ޱ�f�u��1������wu!��N2K�l�c�j��-�	�vߢ;gA�� �b9\�x�%f�$w��~<A��������~�[jk'yҦ~��+��?t���?S��CX�Z�
-��m�������g^�b;Iĳ_�c��V@
�Y5�����GA9�X�g�`���w���k�[F/��>��GUl�#�a;o�/|՟O�����������	���\�N��r�s�!5�[sB�aU��y��V?���W�Z�1����.^D�Q�g��F�7���'`uV�Ÿ�a]��T�Z��i���d��9�?���.K���ծ� ��-[�BQ*"�b�p��4�Uez ,��tyݺ��&��E�7r��L��ic6Z�L��_򒗜I����ˡ�-��R��07���n����v��S�LL㙦�9���|S���,�3tނ�^��u�L��M4�j�{J�! �m
��'Q^��TU Ě��N\��־���g����aT$;��W.(�-���9��h�Sr6��Nl��?<�z5�T-�B�i�t����T��HD\ (�����c�x{�����_�ϳo�Rz��ފR���aIڟ��}������y�	�� ��0K�h�aک`\�XϾ+>�/k<����xh��[�ms%��D_�E|U<��6�k��W��x��@;���%����5bD��c�1�)ל���o����c6;1����`b�W�Z$Q��UX�a�'��MH<Z����I���]��q�����:�<��X�aD��c�K�0W���2�2��yq�V&�m���q�i<�>�e)Z�3�w6�op�&�Xo�*p����1���XF3��u|���JpV��3�ĶF�����a)�;��*���]��T���+�|+ѯ��dbM�ʚ�VF0LF0L��4ъw �j$�M���V$'nI���V��Nƻ]S:�echQA[�D�4��<��.<��o]��V�|�g�Z#��9�w��_ ��#��B���f��w���(������)�^��*7U�\��ß��������dԐ�n��7���Y�L����|P	o$�J��mbS��"�vǥ!��&�O�p_8^�����s�mWýZ�QȒgQ�̡\S��߼\�u>z]d_5��:�n�s�0ZΡ�O�8��=FT_���Z~x�:�M#.��y�:'"�ʨ�������#���@� ���@�W a�hL!�D��������\�@�΀L彮K����E�����u�}���x	����M\H��n�Ez]����A�
�%VT�{0�V�O��n߲�{�K8�]�V��[9�V��[���y
�-�"��o�������9W]�S ����\��<�=��W�ޫ�̹�g]�n���7n��#��U��1��Ex8�>s����-�L�d�Ɲ�� �Kp��Ir���ů`��{�9/� �
��+ɞ/d�]�>��D���X�Q�"�
�K�� �g����0�^(3��?��U��^��
������-��n�.��d�;��|�<���q�C���^K���6fu���ܩz����4禫՚��N��#�6��6��[P���!"�s�E^??
ydI�W��*s�O娹&S~�9�WU�>M4���(>+ad��r٩x��P���q�d_�vv1��������%,���>�<�'�n�qe���G�^p�K�mP����p���q���B!#;Mه�f����a���M� W4�0u�3i��Ћ�".�0r�p&�$ oR��`M&q�N�+�F[�'K��H��������93��/9�;JK��+P}����W�h|;�s�k�MlC��%��Ofm�L���E����/���7��9XƏgl7��84�c���U �����wX������x�ʇ
&��UX���Io�Gq�'�r�@:|^��eT��S�$������r�)vH[�+��\��e<6R�s0���2}˽�}���󼄻*`V%<J�����қx��`�1��W�w&Cw|�,�JCU*����]�iT8���c���yS��EΡx<O~�ۻ%�B]�� �?!��^��A��C�
Z�Xe��;|2Y���"��igA�$���[�R i�[�Z�n̂�v5�{�������g0�3 �u�O�Z����[^�"��f (�y߀ue��j�6Z�U0�c�g��͔$���IV����稼x�� bmU�Nf�Rی�m���	m��#�#��ϙ�Q�2i�0�yL<�U�����clO4���]�W����wa���p��~*��?37�y��':^��UQ�̗*��;��[��o����]�я~t(��w������^|�l�x�F��*J�ڽg��4�j|;?䧁U~#V�QX�bܱX_�&�c�"�
ي�E�	Q�E˼��	U�y]ߣV�U=�)�#�PA32�soH����Xח�g� s�����(��O��z�����*�k97�)s�6k�] ]^�s�y� t�����ƕ�N���}�k?a]�S�3�E���Z�!��vߖ��[.�3�9t���@�2�`�˻���&�G��t�A��Ɔ�H�O�`�)1��3�fO����b%��c =}�G� _�j���_/J�����2��o�]�\�_����G;���s*@W��*�a��
��=E`�,T�J,����y�8��� ��N��������0R�:֫R2���y�{^���so�z>"���P/�/���B�#��|���#Z퍒��R �,U{1���(�q�����|��N?+�;.��Q�Og.}�����0c��_�l�/m����x��b�R�y�C�j�GQ��z�~U�;wQ�a��|_�_	_m�"�jH��y�M~�?��*?�7@Y���D����~z��PI��$��oL�ەs�:�b\���W���Ѡ �%������C��xO��xܘ��^�_x�o=V���t_p��x� Џ�u��m�I�nV� �qб��/�����{'+�2W 9}�XuSܪEa�5��k���LҚ�W����w�j�Ղ�{���������>S������o�G˯�>A��Ap�s �?��=��	�$w�9$3&e��5� ,��;��u�ڷ�s!}�@UG\��ͧ�X˗^��W�7��laz�G�pͺ�y1���ۻ�3S�s �k���3�]�b���k��n`L~C�����W����Mc�q햃�A0�}�[�j�We�Z��Ѣ��(�y�ii/�(~�0���T�;����l�9�ѷ��;���&C�|�'����ڣȳ�W�<��>��Q��=�x��wص��z�:��%X�v��B"Vi /�������M������2Gnfu[ܻ�����3�_��s��`�E�wb�o`'�k`�g�Ɂ�[ޱVd5�X��-ȣ�E�f��WӸ����$��Y�=�ʳ�$��cu4� ��3�� �� }�:��=}Ȥ�sdѯ���5�� \.`���8�9��,���ͺб�d�,�-~��=�K_��s��y~Hswyξ呱�Ɂu3���,�P����Rh�]#�n*��������'6�׮� �c#/'V�5���=���N���R���C\[W�0���q:�4�^͕�Y�s�SV�DdBU����iU�#��qR墏	o]�"~w��"�y;ޤ�bL�jB���	���	H_�Cd�ߕ���~'��{�L���W�����6۲([1_��ܥ�H;� 0��@�"�e?�ȍ��_��dqKP,�mHj;�eg�绕� ��eZ#�a��L�I�7�a�h�-[/$���߀G� @}��� ��g�F�..�C��Up�ܷb+���*�VF�����smګ�Dh���+�Te#4�{�m�~�������P�	��p�,�m��u�����2��Y Y.*�Qhg��h��EH<���1�][C,Qp3'�:v�'��?S��/~�O��1wV����׽�u�%�dxkK��Z�
��b���0+,�$��G��]���k֕ �)�,,�^�E���9��3 ���Z�(pt������[=�"}c�?�k���r��F$r/��+�uޅa�*�*>K<F	���m��
�UN�R��xW�Ɣ�&/$��@>��� ��zЇn�3�@��R�7�K!�|~G�LEk{,;�}��N�ߌ�a�;S�7Vh��a�A\�JJ�ͫM␗�!x/	K��e���隔aL��Z	�z/LA+�Z칟mT�t�H��V`�x������0|7L�`W-���VK��(��'sڬ�d�3����񹎷 ��+ܘ�\�� �3]�
H��m{~~�>��Sx2J�C(q�2]��ƦU��@��9�GBO������X|�eh�ƺ9��d�R�����X�ϴ��'(Դĳ�i����uN���"�2���;+��?��S�j\��㿤����E��x�X��!u�V��k�7���z�j��`���a�#|ފh��T����>�qQ��QJ����I��ek\I��2g�d�,'�'d*-"�{r��vO����C)ޖ�N_�cٿ߸��� ��2�ߡ���`�.~0��H!���������Z�n�
:a(ێe�w�u��¼
��r��S��t��[q��Kf�4���ݥN��PP�qO�B�/�E)���{r�Da�j�Œ�g?Y$���m&T�i?�����Э���dJ;=���߳��u<��L�kt���]b:��3��g2�̆���d���,�Ito�5�3.�Ȕݟ1�>��㔼�2ޔ���+{��w]��I<��wOĵx���2ڋd�W�X����u`.�&�Ww��@�Y�+E%�U*�p�/���^��,�_�v�)�\ڒ�t/��鰥����Vl�A�ܾ�� Å����ў��F VքGvFn���j8x
A���&�B��rV]t�ԍ�k����o�R�wBȰ5����~�=��־��P��[����}�$ڄi�p%f֪˜d�?���g<�y�8���Z�j�'�Pq�U���y��p<�C��k����֥�a��Q�Č�ó�]7e�T�S��c��y��"}Z����� ��y[إ[�T'X�T�<��+6;Lk�����_=��sq�-��8͍�-]{=4��g5�}`s�|�W
� ��"ߧ����|[��~��_=�q���sL�����Z"�8c0�S���u|��_���W���e)����(��J�pO�f-�.��ʃ򟿽w���]�	���1�W�	�#���b�O���"��P9�� �h�!��=riRU���LT�K�/�����0e��(�}�!
�@ނ"9�*d�,��ńv��d�WyW����zI��I��@�]
�A����&˹Bju�����i����J�6,e֛�T�w�-��ʾ�,ۣ�mK@�k&���#K� ��<
��Xw�Zu\c��Y��L�
Xa8��+Ӯ�������_���߉�<��_��~?�L?+(�|��u�D+tB�0��a�X��+���8@x=���x$V����i���0Ѻ��sM>׆��A�݀���{:fU�6���߭� ���o?W�M?�\Aw-/�:=���'MM&�m��V�z󖐵8�uL� ���6�U��Y�o�����<�}^��;����?��>��UV�_W��y\��J�'	9E�V(�r|t
��/�2��x�+N&�n.�e5�����g;��ox%s�a�c�o�Q�����Oy�$�;}��^cIaBJǑ1�Yʶ��>�\1��N\*0y����&TW�qv(���x������ju{,s������{�w� �F-Ђ���g?��'��v7���:��]�H�]rm��ٖ����ZW�Z<�Z#��7e:
��B�@�<��(m�>����h�_$q?�pk�/q��.�q�8g5�����G����њ5�
�<;�h�6�/�l�l����+Gx�� nΫ�8�O�	_@{��Pژ(���G��9���I��KL �ҏk��~��LΛ5��au� -V�:��M��Y_�]��x	ܔa�z5����=0�%['���brXv}5)�f����Q4�!#@=����m��@٘��$�-I���	k����~c�@�1#!���%�-��B1�k  /b<����Y��?�<�{��3��> ��h�Y\�
o�@5�-Kв�<�n����~ݾ���O~����f��EO��ZȂ5����<�lt�^�he%M,�Ęã�#����TP��ב/Z��T�1�p2��Z�q�\����G������<�a%)�nҕk�\i��B�m�r�V^mH��"_�{�[]b�:<��р��
-�� /1cQ�l �.d�DR�Y��jz ҝXHg1��]4�@F�5�`o=p�/PA��}�mo{�i���@ߟ�u�v��3��D�++���2)8og�X�O��v���>�����8�*XL��;������ ��>`�p\��g�we,��x�#��Յ^���@��f�S'�A�M��~G������v
Y�;��~ �Z4[F`�R�E��;y2��$k:����Bq;��0?�_�*?���R_{��cr_>Y�㺮�R	hz����~zg�Z)���F;�\yE9[哼�|<��,��~��X���1��R�Lx�u�]a�Ѷ�QȽ�WM��QVLP��s���]�%V�c���ٝI������u���Q˟�&�k@���[���'!�#�,��U.�D&�e���Z�d���j4����&����*��d2Iܜ�w=����z������*m�{��B?_��k�&r��-���g>�`��Mq��w��'�p¡X]�{�S�z��d�v��)@�gCǽ�� Dv�w7v�טc�_FXDѫ�^u����8P�����=���=�#�������i(��q��b)�3_���.eZ�提M�	B�2~~K���$*�c��wS!��#���N�=���d�2�<�lZc'�~��B�F*k�9rM�Kre�Q��+��ڟ�'�w�˅����U����]������F�p#.���u�{}�{������(�e�C9�D�;���d��1{s5w�k@�a�NE{�B��]�z���LX��۳#�+�NΡ������
إQ���b�ɲ2ݚ$J��},BLs&��O��g��q�}�g�\4�0c��Znt��-^��c�?����&	��H7|{�
P=p��;��xx>ޝ]����V_�=K�6�8As3�O���=刿Cq���Tyb�މ����we�ܧ��ӓ8���#ɣr?�yy.	�)��_�6�ײ�X���~�~��7k��ua!(���ٸ��y��1vI��J�C�O*{9pK�T�9��e�5�%"�eld��r�!�yZ�$_^���$��^=�`�y�j#J�w</����pxr�MZ�-P���޷��f�.x�5�b��f�Z.ɸt��Xh�.a�w��a	��9��n�� �"���{�a�kԫ`�Me��v0m����pC� 1o+f�K��5��2��g�>=�} ���YW�m�đ�!��q�Y����l�F��~��_8��NVai!�}�d!(@�@��a�z׻���ֵ�I�-�������Œ�~?����*���B)���"�b%���W���O6߄9�=�51���˹�;E3"�j���7V�	J�����u��?>��d���`�dqS �nȴ�RH@O$����ȡ�vO�()�����+x&��^��[Y ���c7#��k^���9^�E��>��g�[��}��9�f����.�(,����(>ջ��b��٣����q����b�=�i�~�����BS$^��0V����&�2�Ų��i��~�0��΁�v�&Y��I�K�f"�[�X*�zM4K��e���"���͗c1큋���]�=F��9�3�g2n���R�=�@?E�o���矻�Ck��S��k�X=����qd��:�{[�QkE���ǹg«���>��c�k���Y�9}�W��Oȵȹ~ŬވE���+�!��Z8R�8=�<w�OX��闽�eg}�ӟnC��S �v������k��6�[+6a�jPTE4�i��G�Y�1R�����5���n�U��H�m�)˰�S���H;���нN�aT��*(W0���-��x��2���=�B����io]�5�uLe�K�{=�[�P��F���K���KD����_�ꍿ��//g���b�Դ�E,����^1n�:���2�$]�����ŋb�V�E;_{��_�w���'}`M��
�5�"Z����sGv� ��������y�3�y���kkc8�k��;��B+�>�*]��*�",��w�6B�����X��PގƻsY����luս�'0�6���p�~��2�#Y~�g<\�,ܦWQ�
�|�	Oxl-;.�xn<x�)�%��]�'���֦<�����F �*��
ȧ�i/
A�V�'K�sw�}u_���Z��6��7�L.�5V�D�oŠ��2��24���>A�W<����J=⌊s��tpb7�f__Zf�@g]�Ŭ��_�� �:
�0W�8
���F��w�˱��O"�\qf��S�)�����P�M|�lA��%	���0��?������E���݋��2�VH�@��[zaV��yy�����ۙ��c_�җ~��8N��2�{/��W ��d��N�۳᯽�+�!.���yx5VP�6Bf LoA0����at�wÓ���ow��&@�`,�`m���[�^A�`f��$T�O���A��MXN''�<��*����[o���k�.�%g#`��w���,'��v��<>�w2 ��x��Vd3��\�N����[�|lL�@��^�$�������WV���>�d�zmU�ߞ�`I.�����Yn����%�Zf ]��c�Q ��򞕘O\�ח�M��'� t����K��Yi$��%r��Kа:@��kl'�M]+hc��v0�yQ�� ���7����`���~��=g$�N��t�ue����u]��'��!�~" �9<!ƾH��EM���ޞup���?-|�mۀr =Ja���VxW0�P4�JXG'�&u��-�14u6�D�>��o��?�bw���<�����P�Y~���X�QRcQ����t�߃G�E|�������C���`�a�;nQ��zΊe_��M.�&y2n�X�}>.!��g�Qb���oA�]�\6�(���'6�gI�Q�����ၼ���0���h��^\c��{�*K����_��?�}I(��Y:�'`�	9WkЍ��I,�kY��!��#}`��a0A8Y�2��h,�z�W��K��� yWx��
0�gv�dꬿ�V���8�菁񾇋h�l6Al��}�k�e��?�������3�(�T�m����-�|}��?Y���J�\��g�����r�%l�o|�����'�~%}�A��n�v&�J�xN"���w@�f�п����k(_?��ڍ�|�;���G�B�B4;£�U�P��,+�?)F�z͞�_�Ң[�g @��/�����)�_�G�>-"
���B���Miru�Z9��#�d�A�mT��Ia�Ί��7|<P�y,x�*Ii����f=�׸�Y��kf�О6��%���w�Z=�H��&9W��!��~��_�_]�b�;�|�#6��o��ޒ��J�s���%�ȓ��E��]C:1�0R,���^��w�q�ĵ�k;�~�P����ݳ���j?#�� ʰ�q�g'6Zq7���ޘ����y�o�����F)��A4����|'ô�
Ͽ!��,�zފ?���g�Ӱ�.��/���^���<�exa������d̀x����r�|��{�}(<}$V��&�Q�f;��}�Z"<��^���&14���	�?�?��l6����K�Π�z+@t`pb�72�?@8�2���e��c��M��s�='�t9��:C����k�k�,�2c�
k��WgX����xۑoUL��_��L�����ϥ�k�$�e.&I/�v�:_��x��yY���o��.Ua��e��=����V��K$�o��[�a��3�k#���z2��VAc>a���}�s7��%/���-���"������j�2�ד��%�����W�i�u�8�-oy�Y�x_�`�n�70���Tk&Fe�0h�>�I��/ޔ�M��>�x��Xe_f����������5��0��������(��sh�~�b�X��1F��{�&y�A����l��gX�B��بe5
v�""a�l��Y+ɚ�q���!��d�W����}ޜ�Y�v<@~0�ޏ$��F�lq�oks�R�%��ӵ�߇a�<�e���;�|�*�Et�j�צBgǫ(���.��\��w�������L�T����u�8O�[�}g|�1����GP��걒�v.G����k��U��s�M�?z�jU:�}��5��>՘�KCV/=���)aZ�ŗ�I@g�B������#�M* `K|B�I�܇HD{7��ߒ�xB�$\��;Jr� ��I��2)��d����	ce��=���_�?�5���&����+��m��(�c�U�,1��V9o3�c3�܃����/�����s���n�	�6`���P��EHX�pz��Ǹ�i�2�c���x���Mx�N!~�+ �0��}'0�e	�����f��+(Kβ�<VM<6��#��k�/}�3�ɘw��?�я.,[��
�L��c�D^���O\ğq�1�ce�.q�5��v����4��с�V�
���<�8�#�n���aK��l����d8��b�?lAH�입�>k�r�smC=̅^Cds�˹}�μ�g���TWL����1�6A�Y�k���}�t����lx�3|��q��c�&�]�(P; 2�~�d?Hr�'��0ٙ��:(��ObE��m�<��G.	@s��E/҂�0`��?��ϯe�<Fr?�Vε��yE!�wb<�� ��Lȍ��y8��&V��d9�CB�<�5-������X�0Ė�to����
�<�n��9�<��Ō ��Zx.�5���-�sI@�e�⡬'?��\�,��~��%w��
��b���TH�W�-5�Aȇ)�o�'r�^���SU���x�֯�@@�oȀ�ോ��7���{��	���#�SWY.�m�B"o���o��h��mW��	�� ��K���?�~g,	�.�F6��@�brI�+M*0���*�W�O?*�����>��`��0�1���F�dD9�PG�;�}-�:5VS\��l. �����~7��t�"׫5�i�y'4��u��*��X�U�#����:���_�{g ��<�^�i�d���hb��Ŕ����:PV�C3_���y��Y[������#�q6n���_�t1_�ү��,g�����C9�n���N��X#��������ӻ9�x;m���:�mcH��p�g:���Y�πg��=7A LK�Gދb�������^���%�k�]�õ��2�Ӈ�=�=�Y��V�'�p��]]���t�U��}�߁�����Џ�8�V~0�n�y�~�^�ܕ~�K~s72-��z�*����)	;e�D	����mQ��sӓ����w�B��R)E��������y@�֓�YWЗ���3j�;5,�����R^=\Q������YE✫f��:(J��v�]��e�B�H��- �'pEoĠ>�eK�KS�:����)��Mu�^��t�k	��LX���Xu�p�%
�>/��|�P:���q����n���
@�tQp⊷��#B\��o�"�@ѝ'Q�Xv���p���o��ʁ�)Ȳ%�d����m��F�������$���k̭�8�q>�wۘ��r��ǽ�g,�-)��|�ǘ���֐g<�ORb䂱��Z���������b�%N�'x���wc�gl�K�5܉��92}�����;y�[���{���[}��&���[����k�C3	��y7�����&�n�{��l�70�T���;i��;8~��
�[d���9�՝�k)R ��:��4�AY���덊�����J �7�Ŭ��
���ZY����o[�?����������q��f-	\�R�+���
��9\��]-��������_��(�{��|�j Џ�����N�T��<��^�L���s%q�wAX��K�Z��h�ٝ�߮�ԝ�H�~�x�h_<4��(T�L��E�X 7��R�:�-�A�O2�	:9�>�3��N�`��L@����c�H�K�X�@����a�>��9��L��7h��B�e�z�n�`�6�*؟Ug�����٦� E&&c�U���Q ��s����x=�x�2���#&�f,A� �>�k�ۆ���p�ʽ��I�g
W$�.�'X�����Gq�_�y�#���;#�8�n���x#V�Uhs��r��_�>t����m����O�w;��w@�;9~;mx��QY����G�z���[~�B�܆�p}����d<_����o�.ۖm�.�x�mz�F����ALv�
�E5��V; �z�q�|'O3w]x��YUQAM���H�/���S9�p#�O`G~��qzߏ�
�C+��(�$�l?�S�O���:�+�W�=ϓ�"'����Ď:�������DAZ��Ɯ��(x`�t�@��It{#`$�?Z��@�"|��RM�lD��<c=j�&���y��d�hܫ&}��t�G=�[׾4^�FM��0�U?�_
�ž�}�ɪK8��q�h�I�Rp�= �v��Jσ ��b�����o���b���{�+��3�Z���E�z_,��y�i�[Q'y,�h�ᗪ���0J+i,�O�w��gq7	��'C�ˀ�ִ�|�X.Q��>1�(�q�G!��7���8vcu
<�#� A��S�	d���^���n�!_�s�Y�N�`���DX�}@��:�v&� �]�g=r���0�7��Fi�|�&J����7oA^K_e�vw�m�����[}���VVx��� �E����7��/Kc~.�7�Vzm:hB���
�Q��px3�+����s�*zF#k��g�t�4�Y$KQ�����{�s��͇ѿ�w#|�s3���X�BT^��@�Z�(���`��\� }a&Y�g�����k��>A��>=�CDqYf�A��<c=���؁n'@a����Fs.��&mD!��i�ą���S����$���$�߉_�̈́�TfK�����g�� Mb��@l*��	m�a8����]v �Ԋհ1�:ڌ�z$n���mx��x�5�1�&���;���	���1$-Ɓr3�8�K~^Kq��X�1�V�B11HA��:9��#H"x�  ���g]���X�#�a�5V�$ѭ�����ȵ�*��US��>Qbr���6=�{�a����s�SA�ȱ��\�C�	�Ծ{<���o�!�y_	�NM�7��x���s�C[�k%�Kn����B�l���O U@��g,2n���QCA��xi�ۆ1ye+|kLy������7�����Fxjj��G�x��M��x���1��\��|�8z�.��	�o�rduѓ�$�,z���?�O��%H��{�Pk�$����c%Y_؄�u�; ����;�=��k�����J�.�Av/֎��� ��(��@@��ټ�X��^\C��c�rCƂ��܏}c,,�.�{.9'��5��%�v"V��Č�FJ,|<(Z��Y��#�Ȟ��3��ҷ�����U���(@>����;A��3f��)��ډ�^;�t����ȳJ!ɗQ2��݁ �J=�xt�:����;3���V f>�b4/���Sr�>�a��9��Զ���o���߷�����K�~�+�k*�1�ݺ�~'��5�������V��&a�ܨD��ݞ�� ����?R�2ᘌ��k�=�^��$6�>8f6�o��,JZ������3��	{}�����DI�ﾒ[��\Y�|M�r��Ӫ��B
Mﱅ���Amk�t�U�z�?>��O�
P���b��%�9�&#�e\�n��$�unA�.��O� ��/�X{\��Ȋ$Y=��U�H��[\�����9E�2�way�˘�!<��Z���#2q�"�GurD������3`hc���V���"qn�3���X=/�y(E�/h�����4�!�u���g,�u�:&�i� *`Śh�Ϫ�W�Z�ս�� ��������M�X�Q�|.��M�_rVc��{�����Yţ�o�;q25���p2�(� ��$�_���M���p��[�W��N�&L�F��ޫ���+��W�}��W�̤<ܼ��/��6 �)�����9𙀗oI�#�_�Q4���ݧw�_�����ぬ�>�ۢ~~d����g!6R���G�ʇ��=ϓ9R�/��6j8ɶ�	͒9�����
��
�,��r�R�egP��UX���~? �&���P�j�j��/�i�S"cyVQ��i��6; ���>���������I��Y�`�_������&�|c��x��L��f�13Ew�Z��H�5}cun�V�����q������ޗZ�|��C�d:���&��6vO�v5��qـ�Z.�7Ev�M�:�޻��=�T����s^����� ��S�G��ߡy�� r#ןI���I�<��-V���F+�Ⱥ�}��hܿ�X�b~��;��^���0��z��@��1�}�l�� 4Y�"Va,���
�Η��<Gb��8�>��Ǒ'P���4�9ཋ�E��$�e�WgS�(�un�Oa�b9�<w��g�<��(ʁ�����z�����_��_���㊼�e;�SmP�#�#�ðI������.��lM,�.f�o�T|�7����;�����{Q_O8�r�G�?	g{7��� �Dc]q7��Ʈ@ͼh,�$_ �m\�@z �����*PC��k��/B9�+��~M�j��i��; �;c�J��KV������IY�g���@=��9�:�+(��p�����������1�H�X7��T
q��j�������퀆�i-�=i�u�#��u<?�_���&���r��U0���V�����*���#��ï��=z
����3�nLc����۸J�\�1���b���%��@d�H%��~&ף����^;�_-ۀ��Q#�d8V't��]�񻭪E�b-�l�q�aQ��~�sź�i��u�eL~�-��\�n>o�Coϻ>s�A����K=A��$��5��=��ĮNc���XzI���(q!E&w�?�R&BN��_	az ��`�O�c��Kd^��-��Ջ|;q{\�����AnM�Q�N�V�ܣ�W���nd���]/s��C�ǣD�`��ң�#X��%���Ȝ�:ߌ�g@�iQ&�[�8#\��N�{{���zb����՘	> ��L� {�n�y-�4v�����3	[��w�kLC��:��z}��W���#�&��a�G����6��Tǫx�E�G�VYU��y;��P�_�j��J���;�WP=Ϛ�*��n&���z��s��4��p���3/G/ }��i�Gz�N>�����A���yUzg��K�ֹ�g�^��E?��R�	��w��λ���Py��k�j�����+?W��K��|�x�
�T<�� c%��D6AZ�݁y��h��װ��&�V4�G`�
`�*#_Ml�V����w�Ok���F���u�x��ĵe,������7t�b�?��¤���n�
B2��I,: W��j��]�"]��lr�td�!�M��(�r�������[�!�1�0��q��=���c-���V�0+��"��&�笟����~]��l����+�q��CJY����g3>��1~^�
� ^��/����}���~U*���:n���?��1/k�
־���:�
*����C_/��H�҃q��^�`���ʹ3��of�n�n����}� �J���sfb�]��rBt�.u��-��-V��	�G��%r������!B<����nQ��3Z�Z�aXR��
��#�ؼ�xN��M�[�_\����1|��HWe���%y��xrs�a�~�~�1xh�����v��u_�=��}�>��O���͸A��U�QjcW�.�8`TAa"�x�k�ݠ��mL�}����[����OL�����i,q��~�l�=�5�����d�?	W�S��75)0V{�6���-`gFXFxe�&5���L�չ����Q�����q�e2U���2Rg�%��յX-=�#�5=R����?�H�2��i{۽Z���V?�MS.`��X���ۡGc�a�XA~����Y����T � �W�u�y�y_i�DT�wL�QL�Y�3����l*�����Nv����YS����>�o��&��fλ�snaܠb���Z����g��ڜ���R��^�k���m���NW^�~�����-�\�@��z����̭S��0�gb�}O��(�Bø߽�9��.��&����yOY�~����"��k��Y��s�ʜ(�����k>2(
�穠�+�7���J����ԃOl	=\�� },�� �P|�B�Ț>K�e��e�V��9�X�VM����=k�@5�Zpw� [���l��ӈ� ���{�r��W_dk0��w.٥f����g��D6l�y�uå�Z֨ 3���S�qR�ݒM��:�bq�5�\��Ѣ����X왘H�=�T p���� A�.���}�n���C�����D�3�A[g� ���?�[ ��Ox�.?��C�7<�=�`qͽ�^�s��:�&}�97�['�f�#����y���[���������x���q�oBg���w�r��k�y��w?�ibl9e�Uޫ����c�[E3�so���z3�ρ�n��U�����s��
.7W 3�w������ ���Y$EYh�.�q�?�:V^����J{�=�D��\򷠮�H�Mν�g<s����'�%�z�2 ���fÿ�x�3g�xA;�9�R��j�%Nl����Hk� �]J�T��X}w������X��3��3^��%�g� �c`��U d� F�5�\@'��� �ڛ�;�!(O!)���
��B��G,�4�\�W��t#�g�ld6�By|��7Xr+ �+�}�}L+pO����5؆<�'➜,3����>[��{!C�3�3��g��.��G�GІ�} ����X�P�
@�� �5�Zx�����(vާj��#��\M��S���賖�i�"� �]z���܎w�Mk�o]�3"�G��y4�vݼ�Z�� �{�Y��SF;���$Mu
���d�f���<๱�����w�>��6�+��T��{���2mY�r$q+�pVH�f�)o��m�jo�~�r�̀�dt��|���[$�X<D�0ϟK��c݆~%$1��]��$�&zL��m	h��s�"A}a�e,����ͅ2?}�wdN�
 �w�b��e-y�ǐp�TT����$��|���
���@!t����g��y��9�9@�(y2.�ױ���H�x	� c�J&����q�:��Y�vu�LP3�� P�0U(n�����z��j��+���g^jL �Ƹ�n9&��]�K]s|ꎳ���X��~+2�&r���m��y�)~j������-���2���2���o�N���z�UW4��a� �������[:��Zؙ���
 ����i_��;2�c}��o �#�wjnAmO�W�}w1���Q���G=�׾��Xˀjv�f���Z�6&���R-���9V�Z���=��k3F�\�Qt+�Th^��X��#ΰ>���
��n���S?��|��$�)������j��ߙ����>k�wF��X@���.��=u��o_���>�ek��g��I�(�㢬UO��G��<�c���S`Q���>Vo\�|c�H�(�ҖFݒ_����4�c�-��7����	�W,�v�
�OՃؗAyF���|��!���g�[������^����M��M�{s�D�Ư��:����݌f�?�gb��� zĢ��O̸/(�v�	�9oM���\�K�hS�ۄ+��u���ݐ�O���*A]��m��v�9��
�>�N8Λ�*Tf�[g��k�^�$�}����}���Gک1�>��w�Lr���I��1�Z{��9V-�������{xNܳ\w5���[����	�}�s���Ozo�t�ע8��m�8�=���7}P�X��	��q�4�u��Wݵ�n3_<������ޯ?건�`�RJ(�~	8� @��+�̫�w�U�g�)����_�O��͹��$�$iE9N*�����g�<:R����r�Jx��ȁE�O���K!�w@�K��.$Ȯ��5�ת��
Yͣ�
r>�4��O<\u<�[�Zes0�)���b���RL�d��ӗ.��Xǋ��Yr�"'b���r%�;yU9��̢<>�mk*�]��^;Xu-�\l
Me����^�@=�s�����Wqÿ�x�q�l����*��=[�!B0z�9潣V �{[�a�{T�T cfBţF�)���T�9mT��k�} ��\�3�{�*�+��Q*r^�<y��4��Z����sСiȪB�1��*�+�6�q�����X	'3;����#�pK����W#��T�zC����/�u�a �}��24��V�A���s��:6?��]�p�)}����2�
�5&z��Χ̡()��e딿�����h@"�'1��Qr���x����c�g��@��9t���yA�?�<��j�h}�hl�s�ڍ���ޟƊ�u�Ϛ����r�J�`�[�Y	Ε>Ɍ�+�\k���8(e���䵶4p������t�yE�z#k��Bb>O�6����s�mϕ/�x��7.�?�A?~��c�0�7@P�,O����f���;k�_��dwd'�Zi�|�
2a2�2B+��*�r,�&طJ*0V���j��a
E���A�������	HdBT�ǾUm8�=�+-���ĪJH�;n¸�#h*�k*���}K]�]7a���=8���_ �G��%/�����ܭ>�����ã�V ��h׏F�J�>���~�Y��*O�x�\��X�7�6�;�*�Z��=�ې�)�֓��y��_Ϝ�:���ol�bM]l�噓���V�ngݯ*
��'���2��(@���y�r�Xh���P��Μ7x����s����ᯭ೭�b�,�!#7���+1&�wa%��B��sD�7��;��������m1*w̴\����Q��Kb�։y�{g���xF|��L�h��x�q�c�R��K^#�����M(�gR��;ȇoB��|1����z`k����4��Lb��`��]����$�Ia�.��V{���0�Vp�nk�"8:d#H���}K�
��,��K��?������)m�<�]��Lګ�xՖ#PC� Jh�WX"H��Ve"B9n�X�N`'�
�����Y9�N��>�?��MU�:Nf�[�v����t��{N�5����i�3��Bc,�5�3�yg����:t˃��OD�r(�t�z�5U	3g�z�>�ϫU��bR�����:O`���0tV������K��']�LF��B��x%�m[��U���,$�>�vy����m�.[3��26��
�����\޿�Z�DM�(2��]@��[:�}&QZz�yn��x�	_Τ��2�� hc.���}Pg��.��A�|�]�� ]��*�=_�>ṁG��-�۶��xeo��sǣX�H�b���F��p�k��_�F�X���<��Z�[3ȫ;akFk��F`EÏ;��ć�_@���rqɥ��� g�V�'��^T�0 ��
�}�fq���v�^A>�=�XW�Ѡ+`���o��:������T:V�@���
N�A�˚�P��җ���X�&�����w��G���솔s=�q��9�a���]�l�2�,߀[�j�a]CL���,dr�Tp>�QƠm�a���m4��v��b�eay����j{���΅յ<����V�4��WT�ׄ
������9o݀�,�A�}�+�T��Z�9n|˛�	��#����w�3��%qI�W�}�D�pߛ8w��h�h��5�}[@k�Ÿ��¶
scU�r
@(��N�̗H-�q6�����Q&
q�U�|y�qTAW�g�.(�(&H��G?����m;I�K������;��W.�ǫ�|TB�h����W\7�����Sp��վi
P�I�L�L� y�0@ڪ�[Qr�
�h�i+¨o9Wp���B��%
G_�G�fMG�VP�q�T��[���%�1��1�ڏL�>`�*�+7}����N�L�Ҝ�������Q �D\����������
L�[9�f��ꗒ�{)�{	�ȋ �+�Y��ۿ�o���9�c�a�n_yɘ �V��m��V���S�7����|�x��+x��zDbI�nS�J|v�`&�e�R��I��d<2��_����Q��y�c��r`ᎬnkY	�)S����m^CY>��+/$��*�UOB��K����~K��������<��c������K$�k��f�������8�Uy����,��qt�;~Q@�����'�J�F�<�=l���K'+�	����y>hY,������� �L_$�������_N�ţu{�bw�:SlBf�K"����a��}`T%����p�[=�A��¶
��0v����s��$S�[��}N�Z��/]�!p�F@*�|ؤ�3�~�{,�к��+ˌ�trB~z\�m"�`�u�ե<藅��r�{]˾���*s���]����]X���ܮ�V��?v�]ǎs�|e
�|w�R�H�<O_A�{�y*�(�S)֒��q�_��.����R,-beU�*��~���Ô���A����� ����c�Z�2�Zie�k<'�5�}#ϲ�����u�D<P��{{��Yi�	�{��䡥c�K�4�A�Q��p�����UI���Ѭ%w��#��Ǭ�&����S����o���Ϩ��ҍ���p��K����vfq����}q�� H;Nf�ƍ�\&ȺV&�8B�a�>0UA�$��˹
�
���q�	���wKWa�>&�/ <�1Z}�N&�J��nWߺ�̊U Z�w��������LN���j��.���e����� .�XX�� ����`Bͻ&�x�,ê ����z}�k�1w�������䓀L�>�Z����۲��(��0�\��.�M�X���@8�S&�*j*g�.V��U�� i����q,�^��MUv��*��e�-}�2��v��n�q�&/�f���J���'3���%[?=�>����x��$n纹��{��P
 �'2�C��y�iH�l��̹���N�����)��Z�Q̪[��r*i��sΝ?lK��4�����:�#�`�]\�W����ܕI���$�+���NP=V{�j5�f7���׷.#�*��f��aVY��+ʾDکn^]j���|�e+oer\^K��*@�b �bܭW���0�:<�� �~X2[���?�,��$�$���U �gh��54��3JNm���F�aE�*��j莓�Kα�eM?�x�^��CU΢�EX{�`�^,�����P(�@��Q���f�����0������zd�g�]�dF�|��E�B��tMf�����g��m��fWP���lu�G{��/��Q:�T�����Ϭ�G�u2F�7ϡun����*	�A�ĝ[���b��L�g�.�|%ocڰ^y���!�-���~0|�	4�"Ƃ��{a�tZ7����xW"c�8��Иy�U���ʫ��I�?���������Y���_�GWۡ苀�t�Q���_���6��G����fhFƪ���=�g@��{��a��q[V�e�!������o����>[�0�Lκ��n,1s5��
��,�k n�P�d��ı�y�I���d�w�$m��j3k�3�֨B։�p��iߪ�@��x�a�z<.P?���}�Z�NZ�� ���	�͉�%H�J�J��W���8T���s$����ʊ�+q�$�E��X�T��{�u�D��+
�NYT��֊4���/�3���?i��.~�����r��?��WN+��g�s��K=�[�7n�$Cٖ�V1�X<k��Y�r<M	�e�e��M%�(�Y2�ei���@��*m�{��\�p΢��<H���nF�}����+�ȶ��丕���z�ȃ�+��1r.	�ʈxْ�(�b�ma׎�Tj5R4��at�HJ�.�x5@_j���W��������*�]0���ud
�V��&S2e�\�@b�~�{uk'~W����Ե��C��u����:ny-��*�R���}�o����,���"���:���cq�`�a歱J�bBl��k"�df�Sg�U ˉk�lq1W��V�=�� )�Ӯ+�����U�k�������8��q��}0�����_������8��q��}P�}� T���zuR�Vc��Z��{W��(�!	�e4֋`����T�zE���,g��F�گ�+O���_�j���y�`*/��zj�z���<�cQD��Z|���{�9�W��z�}б��^���%��1�58P����/"Q�\7��Ȱď��_A�5��o�a<߷a�?�w몏�Tޜc����N��"�_*�9��)����>�яv�'�8�\�� �� }Y�<�<68yn��a�?+uGdD�?�#�cQ&n��g@�	K�}���M_��>��3XG ln#�YZ�N�_�~NE���{	L[�����nX� ��aJmw5�S}s�D�!�O��!�&�+�U��{���5���U`���O�:n>���bbv�ͼ'q���:���0�g[���=W\�(UoI�Si��ސX�u\�3U%�Ve�6�5[�UoM|��Ԇ޽�O��s౨�ρ�M��J�	���H��Sp���U٨�ZA�>��$.�<�#Оo�(e^@�)+�����2�
��P��b�PH�0QX#��q� mD)D�8R����>��/�]��-?,+�c�X�����3�}��k ���UNs��1ҕ�����j(���o�R�s�EX��]g� ��9�Z�{Y�ɥ�K��,�ELn6�p?v�!����7�f��� �Ib�)L�����բ�n�
t�r��*e>�+T���[�t��5�ـSW�sV���ګ��{}]��F����>D��=����yuW������}*`�r� x\�� ,p����0��&�q��*r�Y哱Ƨ�{:p����@�����MZ�s�(O~&�!�!��ϑ~��9�k�.�s�0#�����whS��>��-K�-|��xsb�
A���������N8��~z�y�w$|�҂����C�$8z�K���>�S~�=��fæN�v�|g�����"e�~<b��}}�U���$V���ֱ�O�u�?�ƍ���֠/�،�s���(k�ah=�����V���Fz뵋G���ͯ��>y��T�}Cv*���\��8��pS�%�j�������?�d���g��x%�̓`�ɂ�@��+�ZZ�,��t�Z��+F���"�]g�L,���+p���Z��\7̅�S���hi+n��)����{�ӟX��S:��
�m�&�o�x� �3q��ː�EY�Y}����� 6��ކ1���&��B�gl�z'��)B< ��X\���;jU���Jǀ}���`�B�a���褸J���;2a��V�	�
�$%/W���ya�7��Gv��XV$(x��V���Y��\Gu��f.�O8�S��Oނ��Zg]��<El��Q�2V�f8�}e�TK>�}x���o��w���q��3N�27!;&��.���qW�_�J%yֱ׭n�J�c�xy��혫��'u�Gt�yS���q�����#���cK5~��?����1�O�͸��l�`����o�V�����?�0P�*��[���>�[��޷������*�R�����d6�E[. .`2��I�S,�3x_��w���sX��B�-�x"�oRpu&�4�ʫ����"��%�MG�:��g��6�2�Uy��ɔ��EY�S`��45�0�T�{M�l8���vjh ��7,=Ly���`���K=�'��`c���K6�ȳ�:M���z�g�|;������J�(^��F�t�Z�\���}�|�K$0�'�l��������BC���	�Gܽ��o����F�c9�d��0��Z@�Bx�5�k8�ɕе��ƎW�.�^����}����ِ�73���sO}�[1&.�	��̯�����\\9oes�� 쯁	�� F��բ*����Xk �.ZϭVz~�>�Զ"l��+�
�a�
�j)F`Wk�*I>�S���r���5����,,�?޿�/#vyKT�*�%�k\���-�UxOb��l���>c�����ƌ�z��:���ӡ�j�𻽦����d�tۯcR��@,�~�<���S��a�����9l,��������3�P�J����ec��UV0�3����h
F�.i#��U.��1K�F�nTϔ�n�OwaKƲnԌ����l�ʀƽ+<}8�$�V�9�P�����<*H̃� �qY%n~�o���Wc\�xl��)�o"i�G��5�0S�qr,���8�?O�}�G2~���7����KK�� }	�8���������_Blww,���e}�]�]ݮv�/���G�D���*�b�WA+&ǆY�9V���-䬖f@�zb�q{�y+�j��L��IV;� ~6 ~5�t����*�-k���5��짙@�{���ފ��%�=�X�Y*UI�d3'�=�Z��_�(��;l�B���f�����U1�>	��s��(qUA���_�ў%�_�.A8n�X��W�V�c`-�d��z��R[��jx�{&֭b`���3�\��	��qʜȚ�,[��2!�w��0�|�a�n"��|��;��̱sɪ���6QֱUu����H��A��^Oa��t��3i�F���ѝ�`��m��gѹc���Pߌ��0�cq�n��ЪIfnj?D��!�k'­
�jG�ŭ�cQ�5^��j�U�!mT0��۠p������2@�|4���x�r�3���Ї.����<�Mu74���x�lb��f-\�[����$����k���l�
J��
��W��bF���������amUk>}��p�g�*q�y���?/W{����,��dMA�g�*�-K�2%��s
k��m�٦�o*�y�����|M�$m��q�x��Q� ��V���I��}�A4����c��H��������{�X�������&�1�����pY9=:�/��$���]@W!`|�$�1�n-�S����H�`�%�
]��>��#?�0��z̳�6���(�0Y��$�ۮZE�Ӌjr^�U@F0) �8-iX�JG`E��^U=��JVp�H��}�~9 ~6��dbP�G�=���x�R��l��l<4�S���|��g|7�R���U�J�w�8雥j��G�o��{��z���h��0}�?�L���ũ���Ū$���}��{�/�Y��3���Jc�T�d=ݮ�@���eMZ�
rۉ��q���<5%j��̽(g΅$ҥ�}��s�������]���v�0
� Tvc{;�C3q���c.8)0cY�Q��d�X��I-|�k���a�\!�ݒ��K��C��>�8a�`�-1��XsOG��Ƹ]&�
����W�VP���f���#�5)٩�)�&+8�z?m�k�I�J,|`��vv&�}Z�y�s �?�z&�ڽ��۲������$[0��6�&�c���GM���_P�DY˘.,A�
�v����c�1�����ͥ��?�G;�zW�4��r�XX�5���5�*�)4���mP��"��̓X��HDю/����(��>�$=��~7����>9W���w����N}��f��n�����x�^�V�K����x.t�J+�LwϋB喱�~��,�-d;y<��oǗp�Y���E �����z��a��n�pX�>A��L�o�Ex�hW�<`�'�X���'�)�� � �u��`�9N`ދqY�x��d�;o����u�]�H��_���o��o~�!<2�<�B|  `��i��o����Vf<���uL�Q���i^����5ì�a�ͯ��G���y������ݷֳk^ʶ�RNx¾%^��ҵ��f.�6�;���^'`�\)���u�v��X�Y��WH�s�\�c�'�N���u��8�� г+k������^'���X'Y�5�&F�Tu͋pN
�Z�^{��G�T���K[k� ��%6~�!�,ʦ��6�����f�̬^�d��I�zo���kF5& L��ޓa�c-��X�����s���N��6���v#����B�yW�y��o��s� ��y϶2�����)��
 8��� ����?�^��F� ~@�u���V��3���%�r'x������,}�� s����Eqނ޿ǳ#��˞%u
�$�-m_���|H>C��$��u���0��j�����*�� @��X�q��$�ѹ�9�v���o�4�,�EA�����޳�Y̛M�9�y��E�k���.�k�K�x#y�D�n�i�'��N��$��/Ijߋ{�e=��}�f�d���Eo&�4�@0���z���V>�)7�?7	X�s�3Z�5�j]�}�6�n=�r�w�-�q;��J��7��z��7ؖV���ͬ�l���bLɣP���Fm��$�r2 ��g>���H��Ĉk�u^m���������ro2�[K����n��\����2 ̮��U	�,���Խ^�n�|��|��X�^��u˺��V���;!����L�7H��[x�}{-"
@S�����蘚�nr�� XSS�K~S�3i.�LI�u<�O@7Ɏ񿋱����K�Ы�"��.z�A֒����!6�r�IZ�W@���L��}��'���Ͳ^�u/��c�U��ƃ>��T��'��jZ�q�����+�v뱺��e��y�h`� �F�#�(������S�IdKJ�~��Vj�ۆU�;찑���	O�@��U��u���ۏ aj.J�gI���s�v'��"� cu��,���#����X�0ɼ�)+��I�u9������1�XΑ��� �v��	��uxq�"��i�>FB-����B�Y����ͣ�X�� (���I==@ӏ���\�xQ�r^`>���KQ@gÝ �@���+Vz�6q��*��=��H����~�=�,�=@PO��&/�[��=Hx�>}gk��m����/B�3���-	�Z��=E��m-ޕ�^�]��16�7W�d��L��ķ�眃e~�ǻy2�K �%j 5@_��ҚjX fw��
�/F���7,���.`��5Y��Ò���c��G� ����qaK-���O��'�u�̖{M&��R,&�U��
q�<�5�q��U�~�fy���mC+>��m�����1���W@_���K���{h�C�롱�;E,c�<��>���g=:�~yL3�i��cg��ńX�H��3X~{9���E�\� ^ǡ��̕���I
 x� 4n3�G����M��w�U�>��������
��������S&��F+YVK9	�IV��><qn���]�����νU(l#n}�M=	�Q*�nO_�Q��=��s6/�Xj�硔�o\�U>]�1qW0�0	���gsΥ��y�֩d�A����3��n�qi�>Fh�5
�
 |n�ڭV�R+\`��^�ڷ�ꞟ���}kt~�,�2��$��ڗ�|q{�.����&Oa\�Z��W�6��2 ���&�G5�7�����mZXD�?��<�@�Li�kv���<�_�*��i;��.C��s�~Ox��D��K�G���,_���� ��$C��W �~_��,5|~�� }~j���n�o�B7�W-�+}4׶�0�.�%��c��� TO��kT++�)ܒX��)����be��ZHDa��6��=	n�|�N�؎�'����w�G$�k3NY���T\��%5&���`��@���Kk0~[�$36�����g=���S�Ư�L�i�~_�����27'�B���^�#��
�����ǒ(�w�/a���T�{��mS���%i�V��f��G�s�Xޱ�Sބ)��yNb���6l_N�JE,��>��=����O�6JY�������W���0�|�a���w.c���
���,O[� ������&' �ـ��,�z���Z���u-P��;�l��y�a	v���ã ��X�F�a�����Vr�Tq3~�˽����N��,��J�X��`�+	v�|wM�o-��5%d]�dB^�ӎW �߾�e�}ЧPР��5����O��q���<=��i4۳�'(��}�N��\n�z�jq�$�G����5n4+���s~~��30����������A�艛皸ѵ�=O���X�q�ǅ�D�����6N.����8��$���=�_���f�|����}��A���;͏F�x�@(� ��B��2H2l��}%Kh�	$Z�&� +8���Y��xGs�W+?��Y��V���oo^.�a��N���Z�� ���N9�$��nO�8����r@-o�v�>�y��ԥ���R���O�V)[��.[��V�V-��ٺ��(� })�ݶQ��P�8�լ{��|�$r	8n!����
£�w4P��-�\-�$֥��� ����G��TE n�[��D� �m'�\��N���n��+�����M�x����Z�u�V�9z]��<.�xb���	d�<��m��I}�����qG;^)� ��C��2H��Z�N�?B@HJ���-��n���m@)��>���R��h}��-� |ߊ�+�,�XܹG���~?lCPu̟���=�� ����5?��b<�#��ݼ�$��X��7Eg���5)��gb���K<^�x���k�d:e!����=ګQ`Lh�>&2���X}+���%1�:�ڬ���Z�n0�- S�\pO1?��-����O�c� s���tP�������P��$��d��ϵ�~����S��E��\8����s���r�ߥY*��m��T��Ş�k���;~�>�z�er�����g�M���g��0�k����5#Zo�@����(����-V��Y2�&qtA,n�j�J��:��
�qS���W
�@Nv��Re-������
��}_�j��w�
]�&�x��]�ybܺ��9��}{,J���䤜n��$�Wn�H$^/��)����C��{,�\�b2I��ظ��<��e�=[���/��[6
,

`^����d��� !�'v�eQ5Q.@��g^��R��Q_�EP��߱��2��ޯ�~�̣Ԙ}��Y���Zɂ�ۗ�U�N �y���[0����U���߳L��}�ڙ3g����
V���}�"H�Q���~z�]V������\�b�,�m4@_��=��K�Pg���G!����<*X��� ߷����?���]�e_���SMH�Q���F_͑bX.�3*������Z_�:�;s�UdrٖH�����jfRΒ�Ǝf�}�o|}����~���@̰G�ã����-[���=v��Y[��ϩ�M�~��O��Z��mg�E�J���y˼tɱ�VH��m{��ae
��}D�����~U ���g
Ĕ@aשE.̜8(��?�b���g������p,��z�oVjB���D�J�%5Dq���ׇt�Q�J�A���8��t�n��>^�,�;�zS@����!��H���H�D��m�����l-����ع�]�m�����7x�}_�v7��'�R\�2.��Y���6$�j�Z�z���:���Ӎ3�s��J�F�c���%������縴Z�_�'�O�뭍�d�5G]�T�8��F�0��ɺ�׀��hx���_V��5�+ٓ�>/�;�DK��1�B1&>�NO�y]/ ���3�
��G���G'u��ӻ�O�����N��z��Q����BO���Ϲ���M����t�ɏ�Xa��W�M��]F�*;@b�q����In�˄pׅ��T^
C���)�U9t�CFx�!�SK�� )M+��������D���˥�N ��}���먌�j6�}��٪�Haak4�C�/�A��_��5�G��G1���#s�X]+�9���2տ~Ƨ�H6�t��\e��.��^�G?s���l��ْ+�=M6U&�o�~���4h�!ߺ���8���o��Е�nyr/l�B3MO�����nQ�r8]��x�D��Ȫ��"�-4O���S����w�5Bb߱�>E�[���ӆ�J6t�MK��%�����5�wl���-��6�di�1��ހ�6��#D��Y4�
5��th���گZ8~0�{W�TrT⑦ׇ:M�K��$rp
�7��,%v�9Q����L��Ʒ<L_�OH,B�(�>��\�p6V\>*��S���Z&rX}d%�$l!%���'`m�iW�bA��M/���-���z���UⳲ���H�0
�1/$�}����d�(>?^p�q���Y��d�����S�����d�R�w��+Ho�@u�'�>�Q3{ś͋��I��,&��>�pY�}�ڿ��У7��hP d�����A��^��L\lE���z����<�@-j�vn0�{�Ld�`���7�c����+{.���X�ޤ��C�*Ub`!�Q�!�#�M�[���;j��_����n��ј�����С���؜����;�y\y�@�!Z�^[b�K��,8p�
`��P�05A�`��-_/U��8���	o�5i�a�2� �h7���i�U�R�����K�
I��GK�ŻEQ�o�5�A�|�f���$L�����l:�-��a1M�݃~� ��_Y�Q}��e�(.��P�k����z��%W�����u���V�#ca�kQ�hs/$/S��Ib�+�W.ǻ��}���g{�Kf���=m�vdc��rQ/�b��u�b0v�j���fl�;+G�ln�<A=�$�|tdˈ�6:⯬)�-������_���j=�[=�ƫ������ZJHt��s<֋Ǩ󞙋ޙ�+NP����Nc�p�Ac+��04��`��-E�O��O?�����.�ߤ
������.�L�����9����PK   �cW䬂'�G �U /   images/fc51afbd-40d4-4045-8777-933d8523ba7c.png��WT���==t� Rҍ�(���� �%C#!*
�J+�(�t+5���9<���Z��O|�뷳�9뎽���{�/t��H��   ���ç    �@��=AVI�  �*�UTt5TT�>��n� @��w���t���MRa�:a��'�8fīN��N{�̷Uy���J��OJ�m�EL'�6<��&����m�����t=rww�'0|>,w>�?/��
���á��,��x�8��)�� C3�iS�m�ccKN�äѽ���&w����DD��HEF����BF��k���JѺ���/�ȩ��A�1/>ܟ&/1��*�J��2s�&`�_>W� F�E���_���tw�m�zr�f$9Yح�R	�1�+����G$���п���#LuNc�d<�������k�lT�����L��k�m��o��$��qr�m�Ox"�<�����v��������,5�ܥ�>>����,$1h|���Y�($�UyB^%�����rh)�w{�~}�����9i�%�;>�h��0�������S�ux^�!9:�9��xY��P��K�\��xL}�3�>��GY{�T���}a^�D ��(�g�@��g�4�O�gL��}��?"��c	ߛ�b��'������62O*�h�����Lf̤�a��7`H����}�0��R�y�ؽ0]}dqYXC�45��@����� &��I��~`B����m�z�Kz^�!����b5�`����!>��Q6��ʰ�h^�x�	����x�W<b˺�o\*�����ӈ�����[�V�i�AD�x����ծg�d������^"̄��er���/�P�G�H��Rks8aj> 1�6�Dψ�61�����7�O'�1F� �eu�|&a[T�I%����da,�kE���cۣ�6��~rWR-t
ɸ��:�tzi:�$�^�^j�����T�I����!��,[���_2n��3<gy��@B6���r�KF��0�.qu���Q�n�JSm�YS���<au|c����m(��9�A��f��%�H+�"&�!~�9q��O�T_��_H �&�V\
&L�F�}�~���YH��O�W/_	�k��({F,/�'�Yͳϓǉ������M��X�+�k�S�fD��姇�_�V��5�3��[x�QSW�ȁ_�`X_�X�$T%(�q~��V����7������_�	�uMK}t�&��5�P��,�Q��_��7�Ș蠾:zQ'YV�T.���x}\��Iω�UMVYV�n���~���~�M���8��B�Ȗ얛A���+�SrFq�6�F.�� IEW1�[�		ig)W�ieWS��)TE�����Q�+�s�.�Á���fN����a!Ռyj���Qï�Tf̤���
Y����I���t�����+���O�O���W!'r�j����$D$���L���qqf$s$�)'�L��e��֚"����{"8k[J���ſ�4�㛑�[<y��}p@`��w�����7%xn��^���{�P6�5P����d�x�)�/_밦���f��L�b�L����������܋iZ�C�f<s~sa��Q;D;���_f��w�w�et�oX��ɴ=������.|0��=�v2����������7K_{��&�U�Y<��t�T�����`��9�=�=�=�������Fy�#v���i����>�?.;�r�<�:e�ή����:�-�X�'T�k^�_f=T���Ց^��.\��&�v�6�����������oj���~��O��������s����}�����َJYv�j��c|T����I�����{��/k���Έx8�A��99�m�������[�2Aԃ�p?��xzl�W��
���_��(�¦�@�P�P���Af�#YV�!��Q\�U��̎������Q��Pu(I��~���b|g���%�_���Ё�����H��i���oKI^�>۞�LnM�;8_O�ۍ3�02�|/[��)�X{3(��c�:ǈ��l�� i����o�f>�v~�������f﮽�OV��'d�[�|��D�F,��\̦o[����|�}7���;�rc����J5YM�xx�x���*�'��w�ٗ�8>r8���﹖G<���R�� 0䰑�?�tn�h\x�b�
��\����v�t���b�+��@�s�j-��?�~^I�,���6|6�Z��`� P��:�=�]���ۣ.l�L�߻���2� �}��C�R��J��V�2��'�J���{��jJ?���
?��[t�.<���j�2*o�;�?��< ����ԓ{|�߶?��_ck	�u��$ڰ'WU�n�����?߅	;��Hg�'�W,7��8�<��/���3�7t�ޔ^���C-��ܸ�n���J˴�s��K�n��\��7̓��j6yv��+��;''�o��7K���� k���w����m�c�uW��������F���-is��y��߳��ۃ��f�׋~�!�Z[�ZB��:y�)N�;���N��	�ȏ�lX�ɗ(
E��c��M�w���ʇ����T;c��"���}G�A:���2q��$|e���%�������/���Μ.�Z�͌��yN�O���嬶6��yͳ/���{����3]�rD4�@�.�+������Q͎�Ύ2���Q�+ ��A	�V�$�g��@�n2�y�_�sa���\0\���	(��B�0,��3a��E���O6W��L�����6Ȱݨp�\��J�W�X��N;vG����s  �x�4���!��h��@�����>��!����΄D[c��/�TTEcN�/pc&�����tr�����(k�Oԛ���띐܁��fq:z�=���a�����ِ�Ӫ�"�����������?������t�6���t�(�Wմ�(Y�q�eXݼ�e�Ѵ������;�������mc��m#ˠ����u;���dᙂi��{s���������05b~%����t��D�^�^�Go��e����F�*���K������~ˈ���9� �6��p�y��oT���`C\.]��`�*4b7x�2�[�~6�QQ;,KW]?�ʨ���h��o�tn5]�t���Q�oB���`��?Y�V�F����a�Qo��E5�!w��q^�Őgx��H�Y�n�a��[ƈ�U��w���Z6
�9n�� ���8����ذ�(&�=2i�X�W��w��n��v���Z=�6��Iv=��}H*���"�F��G���3�?�QI������Gv/\I�Ǖ���]��Z�������B���cI�A iF�<X�P9���5"{]��-�[�q���C��/ k0N�n�E�H���v�Fe�E1.+N_͝C}:��)�^,�y� %՘˙O��HC3�.|	�|�2�RX�w_�(�����������Lg�j����ve��k<�󋱜��u+{���V,��<~�-�'�xp�!j�ФwƝWSg��Akg<���t�}{�������}:�U�q�!��m�g6����(�Ι|���t�sy�`P�K/L�e�T�~~M����}����P,sی��P�t�}0�A
7�y���7��k��/�76},��-� �a���3�{?!��gOˏ��e�_,�RJ:�R��nO��3��oT�w����]��<+veo����+  �,��fY�W
����V��6��X?�F"���D����ǔu��d1P������Z�?J��2s�W���Q��M�R�M����>��^=�����[Mp��FD�Gv�T�T�a���E���=Հ��{�ؚ��p�Hr�s�����'�(�K�ƏX����p ��	3F(�ܧ��H�,�(�	�p�$���?ݱN��xNO��v�@C�={�Z�P�X�N��[-]%?�Q��*���N�yrislG�(�|9S�s  ���d�L�v��n�[4ͺ��4�y����`�cB�-����Xс�M�3�/�˲����a�6X���������b�4��'vc2<�������!����9�*��ѧ^*���t��˪���[B���t-#�MB�(���t��������usC�f�n�BB����Nvj�����~��I��*?{��J�Qj��(�ܲK�	n8z�0sY��_�C������Ot���\_j(�QW��γ�c�7L�Х��d��7I�j�}�Y�k�_�1���$�!��sk\xޙ��Lp�u/x�������v�����w�V��=�z4���?�_��;4k�<�⛊elNpM6�7�����ͻNo��+�8߭6�~���ӭ*4�	&����6�e�m�^�i��Z�ё�X�N%�RE���: �9s@9���D=E�_徱Oۏ��>���8|�����JV%��A�o�Ra�?��̊v����T1�2�3�c
-���Ln�T � �f��Q��Lh���X��>brW&��W��Iھ��uV7_e��^u%�~Z�zR�眪p&�I��m���c�g_��zv-��b����U������JO���Nܩ�7e_�Rc�Mκ���O���A_j؎�5�<#y7�iTip��P��vD��z�N���ev��Vi;�P�{|�^��b�%��29���͠���M��i�Ҏ��d���q�h~�o�P�(E��R���Ҏ���"n�(8s�׆�|Kl��S�T+	��sNZ�@��!-�2xu]%- �)�%��g��;��L�O�wi�m�#�_M�êgAg�c��l�#�[�vfj�g�"���N%��h:��D�c���$�7.�_�w����#�r������#������}J�C�>掰Ys�e�+���U���� �QR�W;	�tW�v�%Aw߁��^��ˆ=��:�k^1��v#2�7W�f�K�v������*Sc&��`��B��M�펁lY����)]����\�F�D�]>��R��:�s�p���E�����(����3���l<��m�<m�����K� ��ƕ�
�0�tM(�Sh�"2R���b�4x��"yJ�?��t�[�"	�"�u1��W�;]�Ӑ<��P�:y'�״�Hb�~�Ece��;���4��W�6ذ�[�y�N���Ý�Őu����eb+�?����RQ\N޲�=W�Ł �� ��$0��D2��^g�C����'�O��$��d�ַ�UZÝ�������&�W��bf�m�/�������f�45܀to ���5���t����>>&}i�u/�O.�q�&�?H�s��P|�ùC�t�t�9!4�f�{��.5�a��TA�$�E ��x)��:i�B��+y�-D�Z�QQ%x�y�����v$[���i/Ozi�9�W�3R�
t~%�"�2�=�"��\cNp�7E<����	g���Ġ���6�&d���J�����Ήa�F�����v߅�(i[0�k����煢� z1O43p煷,e=L����H�qX�� �J�0��؁�j����J<�+��4r��R����,^G�<��MЭ����7d ��'�����5��T��q��q��\�_��+�$���*��9w�	O�}H����KP#�w�����v��IAio�U��t��Ha/xw1~/_�/  ����{��}�[k����̥c݉�0�F!pdԓR=��B6��=���Tg���&�B�h8��J
1�r���M�z��K� �7N�.�|��o&8���b$�w��ϋ-�y�C�7���R�4��	�@��(��8j�g�񖟒$�ҖT[�z1c��²n;;[�sX�7���{<U~�O��ŏ��9 (! �=[%�@=D��Bim Hr����hL��݋���"��OE_fi�+?�vv��T>�T����H�oj	�4�|m�����/'g5�&A#]@}'�����hSdܗ��F`#E3X�Z3l
��4@�C�!�O3��h�!��9;�*D_�
`Sh����DU/���r&ôG�a �`�1�Zx-�� �0��}���3��_����=��
�ا���W�
����c�J�uM����S��)i��|Sy��bI����fh(K��X;�[$����^@g���<	���4�`Փ����',����IKz/F{|꒒ڙ�(ę��.�Xq�˧!�"��n�܃���UV�?��~eO�jG~� ����=*#_���Sc��t�2��]1���f��{�ԋ�n8W���
��B�/O��lǯ>���ju��\�&I��5�D^�,m��<��!��]��{�HV~� X"���zU�P/Ǔ8j�>���Y�J�^��OG��{��s�/�Ú��c4�x����+��0K=z�fos*�|A*�Xٺز�X�z�.��$%��n�<=��,��ы_wӮV׳T���ȸ's�쏼������a0��Չ|��x���8���$�����%*ͥ�O�*Ƶ LZc�v��(���	�V���,x�EVj�N��[�����Z�)=c�[��F�o��m��Ց��I��"��@M��
B/�&7���5�XΤ<��H�K}#�[su�R�(5%A�Z^;ȡ���+�jQI��=a}zW $�&�	$[��^ۦ�Ͽ̉T�N� "��9�(�m�>���v���K^�s��zO���M�X[�!oαuN�d��~���y�Ҝ�ϵ���u�w�kE��[�m�d��P2��n���bt�Ze�X�c5���8΂pGf���u���e�Ԡ�2��E�W��@ �J�C�:���ߓ�<�/�/����������d�_/�خMp ��J�4'p$ё
�烞��dډ��i�x�ĽT�f��rbW�a�WƘL�	���f)ڞ��jh�a��ܰ����Ё�����=�˿t��C���E�2ķ%�j_y"��GP��1U���T�'�b�e����v���-0���0�%����嘧b��y|���9o�C��Ah�$Q܅͡����Nb�r]c�Wl47��_�f.
�SEw#/=��9�tPs�&�A2����Mk1^*/�����v�m�W��xo�\��x�y�z��1����EV�_|��Q�W����X/�;�w�w��QU{4�"qpV>�������hg[۽��W�ĸ��x�f�m�#���X��� ��M���)?�~���!1M��A�jt�Y�֓oŸ�m7C_�&���D$ͮ�"��KF� /R8:h,��O 9(�
G9�׹+*�3Q�Q������cy�(��#S���p&�{P2K��q��ăزPy]u��#ƍ��aN�K��� �iZ��c�M�O�aºZ*H%d��=��*iSo2$�ܣ�ۡ�����f,uc�LA؞��H$p��w����Iߨ�C�I�f�wa�j���zo�?(�o}����ӐГ�h&̐ �Y\v��L{�,�*��z�^��8��2���-��>
�8��1�7��14r}��E���g%!L���L<�hp�lL���~lC�U���"�����"DlO��y�`Y��H��H(�f�ޝ�}d�5!n����8�W_n��:�jIy`����a�|�`ޙ�Ix��#:+��B��S�u1�j�+E21��F�P3��yĻ��hE[�|a"�Up���Ԯ�?bC�l[k楻��z���ȸ:�;����;�Z���)f7����	�����ք�E����ŨM\�H�L�����<��w�����鋣I�����������IO/H�qY��qFѫ.Y��xңI���.�b�'���MQ�3~��7}`X7|,�u;V�c�WIMׂ�ƏAoH`��ʒ�;\�n(��n�0}7B!���C2+Ѽ$���^�أ�i����P�R���������g�?y�.-��y�'���f��ȑ��R�xpQ����[I^,z2���0Z�{����  �/K<f�w92/Y(���X��ś>���I�dl>��A݄��닌��u߯Ļ�`��Q�9�f�z��SW�Ou���0��fK��qXz~�����dR�鶝���	���i�J�)x�WG=� ���ԒY�<�I�U��Uy4kШ���GX������(�.x��Oy�X��>P�~4�GF��R""� B���Ww��.�w0�KOf�8��{���'�2mx�"<�	�`���^a�Nr>M�H�т�u#�1�"��\�� s5�0�r�&�B
9�&��Ѧ����3�7��9��2 q��P�֮f�ޚ8#bWb�!��X�C���t
;�|qw��QB�TW�,�J[���~��y��6W5SE�>�EkB8����	��=ݚ���T���t+%�|�;��2FI(@����#�ۇ��j�1/���C��"���/���ױD���aN����W�dF���W�߷X	���P!v>�6D���b/���T�Fb�/����|�����N�:�5ş�r�<�Vc�d�ʻw�ch��ZO� �hh�܃d;��^�����WF�)�U��.7WZ�������R�<;o7�d#z:�T�Q��"zڒW��]s;�K٭k/F��F�l��Ns�"�Nx��d[�;�le��*��y�!=_��˥�.��2;�|>#�e/a<NF8��4���79Z�jp�.��g;������j���u/ Kq�cM�#@�I��n�63�8�ƈ x�G3;�t���!vteL%.;Ï�-�+]�T�#>�Q������{-��� F�&���<�I��A w',�YUu�(~B��>X+�S�����a?��-�Y:�2 s��'�#� 0���T���v>�
�g����lt'�D��V5�ܧcq(�G�Q��e����_b���;��$*#�G�A����;�M{%��h	q �����T��Bgxbש���)L�
��������O�$!P�pۜQG��d��ͪ1��]���o,l�s�)���l��x��z��X��D� �k'�DNL�j?ʏ�$ȗ�ه��-Q�V�ّ2�_Ǥg)o��A_�H2O<�RݿN����ګ:�����Y��\� ����ܐ�w6Mo�:w��R�o�x����i��A���a������Q�V�*r�b#l(��4Z2�s �,�2��U!��F&�s=��V����kZ~�tF�+p�e�L��#�9�$�Q�R��с+����N�>2ApZ����w�@�������)�W����v��=�nVK���}����r�������-J���c�
�e���N��ʺa�E�(ՙ��Yt��y�t(�v1��B ���K��.,�1;	�v�N=bָ�v���)N*�6����IB�@b��L��8R�%�
��ϫK��4;.����' ӢF�Y �K��]A��:���<���?ұ�~��^�Ev���}����T���%�l���_��/�[�i�r*
��m�8�|e0s��?cљvL��q4b5h.����ߊ[�e�oM��Q܀O{z1>z.��R4�`)��ADT3��N>�`��1�� �>خ$Ăc>����)���Ԝ�q�	`x�a${��z�y#��fY貑���5�N�˽y ��^o�{~���VR.rn� �HFF0"�E9��D.<0�\c�*c@Ux���c&@B��:y�s����v{�d��M*���20�m0�Z�v�5�j�+����VJ�8;��u��vk���#P*3ժ�7�;��}��y������p�q�J�I���;F5�U%��d:FT&�_rT;%�Sd���ab���}�R H������3� "��	4<��o@�*�p�H���H��͒�t���1�* L�¦;���>�Y��z@���ݺ�/F�,* ؔ�gM"T���!�8�ӟ/G��󭷝n��x��Bb��=
�+÷&t��?2�>�8~-'\A8���%у���N(�ا�Y����H[
�y�PR(e���&��6��5N"�ڭ�3� �1��-�Ʊ^u�q	ԯ�S�,7���4���nA�s"�A��)E�L����)A|'"t���X�p����`�;d��c>�]��h/��t���s�UJ���
s�~Z�|��ˌR�#i������ۻ�B���v�H�H&>G ���w@IW�E�Ig�P%�gs���Ԍ�)%�������n�`�3oG~�w��8})�@� lS�_6��t"OR�e��.p�p8�Pݵ�r�LF�,y!0Y	G��'�/�I 
U��$�6�ġ�u�x(IW�� � �3�>��%��>��ni��h�b @;�X{F?��w���~ř*����%YW�Nd`������>ų/)� [�* �8�-����{|zqZڳ����W�x+R��.�����"O�7�%�����aǳY�]����-��)׺W"��>�E�%���jJW�3��}�m1f����9��x�/%,�K�-b{sqw����[�"n��ɘ��ǧc�$[eH���~��Z!�m�*��qOh��V �M|��VX�|��.�gr�
w�wwiA1�j�qx������� ��e��Xo�f:]��kd6�x������^1��[�'��U���a�P�Y��h9r��x+^�|��K��X�? �#�L�c5:A]\xѐ��V5��A;��/�P��g�sss�s&�yT+|�R�15�����[��"���{�jB���9!,�/�=�'����N�����'z۲53�t�T�c#*���>�6G_5'9k������ ��<�ݝiz�3����#5��'�-���]�{*H�ŹgzLl�=�&RQT`\s\�y��9�E�X���Az�B.-���22���!�x���f�b8@��@��#$s3��]b�J[�����ܺ�0���}�{ow��u{�O�DP�Ľ(4���=t���Ō/<o�&={4lր�d�)y��!��=��c���q���_dw^f���s��	�Y<��+�K�~�VB�
�<���˵y�nE�������p?�. ���p@����[�
v�W�:�5��vxBRy/
�JK�<��+g�aD&��������U�K��T�D����k�y����S�a`��K��.��'��k^�t�U��Gx��m���J���͠���eŔ�[�f)�H*}��"@$�-v�{K�	z)���j����j�t+�r��)�R��s/K	%v��;�9�?Ib-m?f��m��p4��0��|?QI���iX+�EJ���5���
�Ha'�׍C��%�@�A��!��3�}.}@%K�נh�f���`�Q�Ք,���{w!��}۔�7|��D��p�l��
H�	gA2��v�Jh���^�1-�g�/DC�GF�P��x�=��F��5|�U!��!�%}�s��:lA��Joe�u�N3��~�y��ZkA�A˓B�va�������XYy�,���10=���ͬJD�è�M�%��k��ԟ�R�k��W���?��p�ݜ7�ɖNi���Oy?wJa0�  c�"���n&�A��zӄ��#&��#L���Z���Zg��u{��V]�ߔ2�W�OcQ�����5����]9��v]վ$'+�n�4�o�����ۼu�����6��Q(�SӓU�,�w46��A�cĖQc�l�[�a��L�Y=�K�#��Ѫ�N�bL�QyS,�n��d?�9��T�w�@?6�F�$O>@����74QCf�ru,}j�Rd@}�?62�l���ij�xp�r����ui��ҽz���l.oW	i�R�@�je����;�� �M�uk����<�SL��!{���JT�E:���#�{��1cd&Y��U��Xw|C�)�5zV#��N��
V/S�9�7�i��N���@�=@��f(֗hSƹ����R�^W�{
Q`}K)������^�� �m雹��W.���� ���o�j���� :�-��}��(��п�j,~�������M���ӥF>�ţ�I��ͧ3II]U{����j��=��������%��7v�(Ŧ)�Y;��������b> !��3rym[*"�az���|Y��m.?����HBP��)]��~"A{jT��'���8�����=r�/:h���8H�~�	yYL�����KۊW��^aЈx��Nq7�!�ҁ��uHwp.�u����_��!h��"#Ը�Tk���1
�;���l�y�Hc�{��(��>�kͽ{��	�t�E
g��]�|�wZ�;��TC8l�'��.��6  ���|-��T��P��b����=D�B�ќ�8FK^�6!�f�9��7�S�˯���=�-��)��v�<���$<~O��c�ҟ�q�1z�j�����QP�S3��������������/K�<㗆/�.�?��J`Z(f8��ls�' F4H��8d��T��I��!_��Ȉ8��ެ~L7�B�D�!ʑ!T�+ժI�jO[^�=��!�!����oS�n��l ���k%���c�Ht�ѠG����a�����wK����o�M#�M�m�9TO��N���{N�	v���[�ڃKO�5�7@�	[�p����1k�4�ܸ���WOF'�Q6}�K&@2>����������$���0�qsKo�tnu"�P�j
�EE�����:��)�9�o�]�����48u+g�ʸ���eI�R��q}T#�|c��e���h|���6��;��#��Q0RE�4�^��-w>�jx:�CT�HNV~F��x�����CF�������HX��Gc�����p�*��j<���Wt��`��my
g�zp'�n0�W�`c��`��{��iv��P�"���!eIPč2﫥���k\�ON�w�WɅ������$.��>���g�G�X]cO�p\�Y���_�+���(T��2\ʣ(���FVF�z��Cn�,7
�MΪ��`Ĺ#h��3�8�ID�;��T��{������4mF����Jk
�y&Xt{�l�rB��ls�S?w\ l�H�9F��/	Hr��$��G1鈦�f��"B��
���Rڷ-��_H͂X�RE��	��� �J�(��b�|!�J9�g�����oπ��6���jt1/K��.V Y�*�Zg��³!�N��~ �{SŊ2���^>o�ȹ,W���ƍ[�s���e��D6�#�_mj���ߐ&<��ٰ=.�|����,�B��YN��~�Ê��7]
g5�,�)I�E\X��b�+k��9����e�����1)4�a{��w���doa�&T���mίG-0�u�����ʕ.M
dr{f��At��K���KZ�ݳ6��[�	`ݨY�U���O�Ka]-)���"t��Ef�Y�(�&'X,����݌ܹu��Z��ȟ7��[���p��UُL%��	0CE�ۥC║!�켿* �aU���(�8ZP�d�w+d�x}�^�cTO�� ������O���ϰ|B[M ��i��I@R8���|]e'Su�V���A$��@(\7�Ԡ� a��P�Y�л��y.)6 �!��ҕ(OK?!,����6��(��D����͵C�)n���@��s�=��b�T�Đ%��a�]EI6kuE���Z]US�H�kZ��(Q⨘,���Ugf�DU���U���O�g��)(�y�:�7X���Zx3�vPG��d͵$w� ��Wc����׺k=�l�wV��2��d����:��{�-'@���}��)U��{��($3x?95o֧B��gR2!"Y�I z�"{�F�EZ	����R���?�	�O��0�Ҹ�RI�X�������	��4����M���n��`��R���K煫t�^�"�.�¸u�Ϙ6~d��fws�u�H$�0���Y<~��,��ȴcv=x�1�ɤ�4r=����H��C������o���B����g��&�x�T�[�{���i�q���n�B�8#���/"����<���~��V�����GO��������������N�<o����%��"L��N�(���
�o\��ݧ���2�ȳ&K��/����i*������V����/���Ĵ W��n�������S� ��4"󁘺/71�ޓ.M����C2
ؘC�g�^W�4g4/�M�[�2�S�����>cu�ږ�4ȗZ$�~m� �NEp;���G��SVl._�7 ��iI��L��L�{�~	��8�H�&����$+�^m҆���ƈ���=�R�YAgg\��"�&�眍�<�D�?���4�F{���R�������	U_��TP��ST�s%�q�r����MKra�D�y:y�1�I�|i���������1�R����R{T�b0��Fѥf4*<��w8����;��޵ t/r ��S�N����_���e5�x[�&:��*�ng���c�r��r�-js�mu��	難; l��[�Ͼ�!W̒۴t��&4�m�ε���*�������D&o?n��?���Z'h<-����wk۸�ޙ͝�j4<۳���Z#��Vw�N/���s}A�μ�O$u[����H'�<Ʃ�Ռ��+�l#�K�T�۫��mJ@_"��q� ��
�ﰻ�:mP	��=�	��f��Ђ@�L����T�w��J�.�?�4of�&H���B�P}:�@#��r��*���" �MOYw1�8�AȐ���mk��Ν�G$W@-��$�������D�Z:���]��MR�N��@	�֚ �*�Q�cٓBw4�-�͉�`_RF?k�P�_9߿��ψ?9��t�������^����E�=:���i�R�������|���	���8��
D�H;0"ҲR�N���ѓH.�{G�/⦯��M�i��y������+	�9��g�Z�~�� S��W]Zp>����?+�n�4�P	���:�W�Aˁ�����f����4�Y�\��*;�I��M�H v��1}��eL6�c���S�x� ���y�Į���=<�O�D�@����}a���Bx��c��z4�m  ��3l�l���X��p �w��	"���J1��To-)��*ƭ�(��#*\.0��f�i�������
�OrA�v:�Bz�^ˎ����Ǘ^ڗ���Y�6��06)�$��];`)X�e��Ԇ���Ò��?��9jԅ�,�P�i�����	CgY���+߫�h��А X�󸍣��<��_�e!�/�q�,�jҟ`C�|���A*�-`?�la+D 	�N�]�	�N�_[�l�ȔT�I���\CTN�i��	k����c��2�9��P�����r� -����z_I��JM
���Q�M%FHC�r~�Cmb�o,C�s~~�m3���W<\�zq�T�O�n��(���u���N��겟����g��NT�.�W��:X���Ŝ;P;�Z��@�9t��7ۥQ��fl��Z2�M|�k��m�IE���E��?��hx��I�qM8mvX�J��N@& u��xm%�c),�֩3�q�;����Gµ�OxJ�Ҝx����l���a��_�֒كF�7#vn^�;>i/T���r�B�y�:��cG, �k�+�y9�9�Ɯw�O!�*j^3��a�΃��IT���u| �/����vw�7V?��i�wu�| �THiNʅ!2�^#�8��l�^\�)��3�n�BW$��U��:w������W�̠���w�/*���//R��K ҝ%C*Œ� �@�\H�I�p����#�l|<���i\-n�>
E��|�SV�޺+�E�7mX_�
3cu��3���JQ�q�Š��,�h|4	��╟��Lq����g�^e[��U������8B��Ȋ"���l�<o��#�����Qm)��/a�7=bm�ף��x�rp���P�D'coC��� ���ƅ�8�p��Y4ճ�S'am,9}�m]O8m���̓otf��G/���<���Q{"�[=U1o۸�i�hĲQl�rs�c��j�҈���-h�.G�֬����f��i��I(i�T)���޽8t `X�A	s�f�%`���zn&���򟉢�n�7���{u�O)�i�pr:���d˅ߪwgG`o	�o��i��j�jjD�j� ݱ�������*�	�� m�Fq�<WVFV}�ʒ1�������i�Ta�����_��T�74�_]r�l�hn�}���` �ǝ�m"���pt~Mvmx���EBj4(1@QJ@z�4#�a�RJD���;6@@�SJ@�.��{����w�s_�s��K[Ԋ��H� ��D�EW��?g�<�5��ж_��R�3?��2.� ��Xўy�yb~#^�K�"7�%^&���dod:�%�:���Z4���}ocA�v�@��o���s`)$�7%i~�+�*�eXc����O�-P~Pk�un�"~�8nn�t���𱴴��: S\c�+�E{�$g�m��[0���~�}TL̞��a��)�}�Z�;{�~$v��h�^!T�7�Y����A�]���彼`���i@AX�1�t�y��I�w�m~�R������-��֯����X�P���(����w�F1^�kY�r^�.���~�-���2�����s,��K���3���H�T��=�g�����ai�߱��3�����c�M�U;���O�e#:X{��Dyjp��L�"��^��-��U>9�s&�c���	n6���M��?i��`f��r��SY�؃0����B�,V(�1ʏ�UG�<��z*H�M,��a�,ۊF�b�E�\��=y�	g �������ިA�ȱ3�`@�?���g{uuD"��|�h��`z���L/I�$��2�Yf�NjY�Ȟ�-gH��}2^Ƌ��X�i��K�e@�ʜ��X�?j�_n��0Wa0�B��Ǐ�HJ�Vm�*�:7��\r�kk������)&. @X��o��5�����D�������՟��z�o~�As�ͳ�䛒&c	��j�(�1�� ;��Է���_��Ń�tNϾ1�͐�D�0g���l7".K�[~����[:l����R�����J'!v�ɖL�L������$5�n��%�:g��ʒ;R������<�%Q>&�����%�����3�b� Is~�B���];�w$@قU����ؐ�;�3��ܧw,�Y�x����9�PxWMv`���##�x�����a����uN����<����Xdr6 &jh�;��6�:,�G��z����Ycd@�	�ox��c/Yj�'�����$����'��!3z�˽t�K�*��I�����	�}��Q�#!�6�vX�-q2�)��Y�q^���G��̪@H6u(`�j�~�����s�]�Z�6�.��[j��۝\���	�^3�a7���T����$L�V�-��N���l�U���jG|�0J���,u��9��M%�V�������{��E�!<�"���CX�=��^��|��+����-��H9��ހ�������$� �W2�OQĄ�-�o�J	��+)�$G�E��,-��I�\t͔�e㱝5d�V�;lͦ����M���Z�3t_#�B����
��]���[x-,j��"@Q��OR[���ώ'O�b5�V���`��8�߈@H�af�� �Nt�5�|?B`����� իv��(]��\�$�	Cc&�E�ƍ�Ғ�t��e��nM	O$J���U�s��K�?��g��Ͱ(�g(O�u$��W��|�n�?��%�%L*����BW�����#�����s��{3$�g���CO����%�g%����%��1��׷G-���{��	�(�|"���- |���ɗ~�K�4������ܐp��j�j�X�ų���;�bo��x��kG-�R3~��H�g��;��)�Nn�~�7e"b��	���5�M5�|�CR�AHKW�(��	?J,�n�"���>�D�*��i��y5��M�YJ �x��P��l�&��E��z�2�S�y��RW��yӂ?m��G;���'�ž�(�a7�E�$�_�0���F�3X9���|u/���/�ų��*n���7�t���J��p �륱�s:�����A�$>B�Yt������=���&��n�ϣ��!M��Ya8���t]����x� ׎��.�Ȩ(���X��UHv3]6��<=��?3��R��H4����E���p���F���'�v;�\Z<1�47g��;�����:G<��O�ㅞy���{f~��n�V�9}}�baV���)�Ia)s��:$�ᕔ�u�סz�����3ޠ&�ÈJ|S3֦�6%�-Yu��Y1�˲n���W�c��-x/�u�u�;�����aq��!�� q�N%0��	a�>,�(�a�������=��)��w͉�� ���ј�3�`��_p[jed�wyfhwI�>�o]J}yӎS�**O>E�ά����[�l5���?�ur��b�^e���#�7"{(WR��[i3/PVTWn#9�d�ј�Ίi�Q�L����̌�փ���E��H>����^a�����������? �t7)T�L�f/`�GON�a����.�r�$d�,��˛���sƏ�)�;��:�'�X�IY�%L@���Q�Vm>��\)�PKݨ2�<x]3U��BQ�mt7��ݍ$:;��C�d��	!,��*%��,�!�QU�tu��+����I��֗�!��2B|�厄J�+o����I���J�1��]�=�F�����\'3ڟ͆�ޛ*i����Xi�������u?�EFZm��) �q(A�(��u�P�,Z��&oέ�5 X��t�^�@��4��O���c���2�<�D��G��2����ݽ��2���fz�+��$���lv
�/�o�*;eϫn�p$��R�K��6|��	q��8���M�[ʆ����n�n���1�o��@�w�j>�Ec��]&��w�a%��r�vܔ%�C����w��G��V$��k� u�'Lt�� �3S�B���@�޾m-ȔWl���I�0���A��� f��}'�p-w��t����Յ�!w���	O���e� ��ɼ�J�!��$�,�{H;8�?��~:�6x��YE�c�x�_w+"�w����mw v����w�;%69Wk�G���Tm��3�S_���p���wK�u&9]�W��LB���������q�0w��GZ��4�q#v�@�)H' �{�X��vh����	�Di���������!�v��F��~<��Ԓlػ��F4�C�anJS5q��h�Hf��">D�H:�Ў��}����s`�.f���cWi�+����@�ǚ+�)���k|Yˬ#�;.��һ�(l�T��X��%�k�k�}�}I�0+O!�e�\xm�u���N%2��s�)݊,Kf:be��{s:Wr`���Ci9m�T �����(����A�w���
�x���;Q�4�s��i�s�&�M�q�Ѝ�T���~N�����wN��p��"��M��K���yi��D�U�����2#V��7���Fy��Tf��Q�*��3?�vf�y���� X�1� hzHw[���K���Q_q� M8�: *�F�N���=���%��t_�F���u/�N�y�/�0�4�f��L���l�Y$�!��ua��o[KX:	�%��]�_�<�2�O�Z4v�i��6>c��af	H���(�����!I��}��\��O��Y�o!�a#��k�Z�
%�����^�FW���q���7�a��"�Q�O)���LU �e@�H�D�7���xv\�/�t~������6���s~ٜJ`�|�H�?fb��hm��-a~�S�!�F�&5al��lI���jM唻���a�����&t0�	�� 44�+}�!k'�q�������ֆa�g?~^,]���:)��^.�?K�Oh7%�s����V����d�fFҼ�\2��;����� �	�g����#�i����
]C� J�a#���,t(�\�;`ؒ��O+��ޖқҦs��Byٍ���.���8�~��m�Sh7v6�eU��Z$n�r�,%����:*�����@U��2�b�4`���z�,�&������W`C�4:�?�8yx�7$��
_�%���*/~�m:�#�P�p� f�s2�A��n��Yc�>F��܍�v�n�.Z�5S~���v�����,S�zʟs�!C��醋>_�$G������\�vMN(yל�i�]�?g=e�#������P�rQ"��xA�z��Z���|�Q��J�����}���;����	�)5����/��ԇp�����4�T?8y�0I�tR.ԻĬ���`hx�lq1S���msbZS��:�8z�aP����`ɶ+���3�.��9|1,]zgz����~����@����n�
-�M?���Q�}�|����� i�Ԋ�;|�{���м�4��x %)�}[��J�"���mhv�RE߯�3ha[���s�iGs���|]?�.С�˚�@�g�Ӽ�3�?�T,��\̰��!בּa�n�I:6+�ԗ_Q�����gςo8��kv`�G��*�8^Ie�
6��ȭ�������@~Vѵ7��=ε�!�e�� ����RO�mJ�ʋ� ���2P��W����E��8k����ʇ��IfuyC�bjqS�Z�,n��~1i!n�1/7ߑ��`�k"we��*��(C��l��������-0h52�ŉ!��l)�%�A���;!�T1��5�{:��aI��|f�DqJ#��FG���rxLKh��k���y��A�*5l�u��n���===߽^ȕ�>T�.�5�qصٞ1��y���K 7ߊ�hɤt"i���r�>&�A�2*̋;��"�� �$��#��'���٫���]Bz� �c�(�~3��q:6��=i��G/�>�G����cj�Ȱ�t[��!��앗r�4w�a��!�^ug"��o�GÙ%S��[=�Ϻ����/���I�D��LL���ԫ��2��$&]��֍&C�����?U3ܽt��3Ap�>̽U|C+�oK�n|)Px�bȖ��C�s�l����kV�}HƸ��T< �S�y�G*|��U�j]$誉Ӊ����X6�| �LO{�>|p�����荭
�Ә��4\U�͊�b$րS�� ������y͓�bk$jJWJ��c�^c)m�n
���미���O�7f3a���2H\'�~Ef���ڸ��`��mh��<`S��G?�ZrW�H�&��]�{7&�8y�?�h�N�V��r*O����\B�����T0�j6l;l6���[�$�b)]�g��iV�����8��XO��c�N�+�ciK�C��J[�o	Sb��7���a�.�.b�J@�dZ�Ŭ� ���L[+$�y��B�*zṷ�z���z�>���m��D`%�\l���x�
�z_�^aV�^�z3�K�������v8I*LʯIi��$�B�ǿf���]v�xu!���r���z�-�^�����>�5��y��>f��k���"�8�y�:�2ZO��r� �w{IT�^1�w����4�hcO1oi9�lj��9�g	@�.�wCc�T�.�.[�@������6�K񹣶�J�_	��$��V	�i�6��-������]^�4���*��҂�1�s=}�B$Rp"�Ǖ�D4?ك���S	��fQ��h�OC��wz���2=�8�#��r�0�n�af�-f�T�+�d�#Ֆ��*�x��D���g��~]zҰ�ka�v|M�L����_�SAl��5'�e�N9��\��MTs����O9#���fp�~��x:˰h=����hL����؂��=�wE�&��u26���l���>�[(_�p�'2�nWt{-���\�a���D�3�OQdD��
��%�Briݴ�|�j u2���~T�cS2Þ���M�rv�pXXްs�z12M�t�M��+�4�&�w�80uV'�fY���;����]R4�G�x=\��xLC���H�3�M��uvX�-T6<���iL�����$84��_n�$�_eI����� =)��T�\<R�-�,�K����ᐁ"m}�v�������O��=�Yv�t�__>,V�J�N(���F�7]�3f0+%p�,��\T$�;��N�?z�3�r�"�No����.)���������WK66��K��,��{BTw~�9�K��1��r��S�|�>�=t�g�g ���xƱ�����df{.rS���s՛¬�6~Vy5s�E4�EX�FoE��_6��YG�T�|&�q��}� Jq�1�I��w��ew�@@��l1�@����}��7e8/���d����_�������9����L�k�(��N�y^�z��*׍;�uZ+w�U9�Ϳ���G����������孌4.�EV�,���+�_��]��$k�~���Ց��Ro�g�V�+FQ�L�_6��~��*��Z��G�B�2���g$$��7~��8lH,��&^�k\��T+���k4�?������kuг\	�`]m��g7���1I�<��  7�)2�RZ_���ʻ�Z�ۓ6W6��x�P�aő���&�ekZ�Z�ݪ{頉��|ńtE{��
�p����`]|)xW�N1�B악��ǃ�7ũY���}�K.e�^�5ئc޿��R��:Z�����ئ�7����Z���Y
���.�ˤ�*���샶��%jm�ǖaE�N5�� ��%��H�D��zH�E������̝?Gp:���r���b�v�M� ~�3]��F�i�Іg�3�o*�$z��؈�JY�wU���G�C@V�� ����@3���Vg0�0R�B; �[��ݯ�lq�l�M�=���(gX�g��ɲ&�w]��h��dI��cq�ޱ���cg�O	�DO����k#O׎���{����v���8�z�6���m��|@�f�| 8����u���"=�fC�W�Y�?���P���֥*;s�ߢ��õ�_�2�'LزG\]BM=u��^�: <��hL�0�մ���D�i�Q�����������,��u�?[�O�*�ILj��|�HJ��s)�k��T;%�q�vxT�f�P��;*��m����+��9�¬d�yt�t������R�B��-Q��Z�L��U�rx��W�G��<-<� �|�%�x��HS?��,�[�� �y�p.[��Y�5����ዱ���>?H�:�Ož��Is����
3��pXl-������������X��c`��X�3R���rFX�D��Wͼ,��y�S���(g���<�*��hw���sf��L���y
�H:�|�Go��%z �ᤋ>�"(�z����ғ����S�o���#Z3�.�"Z=���_/���Y���-3�{�&���!*Ӥ��Q"���Kh��l�ѿ?����qu���}9�̏^XX����~�O:�j������D�8<����5�	/��?�� *@�9F�J�A��_���7�K>���y���2��k��mo<#
M��K����߇V`{|�Ʊ����p����x�qS��N�����| ^m8����!J<�h5��ަ�>7����iys���s��		��������^�"������yD�3�:32��qY��zW�f�V�2�~��/^e]��3�Z����XPԠe�]��
��)2-��D�}؋�F�V��Mk�?ߠ_�h`�y�B���]?S�hG��{n��������C�J�����rD}:�M�>�1�p�Tag�X�~�+L�����l@�����B����*��5�L2���螚N�U���}�3�zء���;Pٜ��z�@m�3CdvIp�����Npd�|�ܡϠ�t������-]��8�n]te@|�P�3��긂w���n�i�v����r[���da�#�2q��&�%�?'/�D�Ul�ȕ��*c������˯���L#��l��y����G��|x�*Gd�1�"7h���xs�Ɏ�����,'�oB5ث>B�&�V/l6�b�~�Z�O����mEc���gS�E>��[�~e��i�8��{�2�ͩ�f"�ic�ȼ���9�XO�H�I9��� +'ڪI �O-M�T@q븖<�Ь�9V/�T�4k���T"�r�p�0��O�^���z��^��T�����h�Tr�S������*�8{N��S��W�����$��gYx��_��e�5�2�}��`�S�VS���JV9� y0�F�PմSߋ�ڑ��)DP`B<K�	�6�K5�ಲK�p��aQiU`ʎ#�x��4���3^cE���qN)Ǖ ��w0e�t+G<:���d�v�7�pg|^����w�=d�u���Z�Z�"]hoA����w|�p+s�"��E�,�%sni�vVݔ
���)Ѝ�,�>�qGQĩx�t���r �;-�
�a��hOT���:V�;��0���a1�K�L3{��%�e���C�����M�hgӳ\g���z���#P�����l=����Ȭ�[������O�,l���a�?/^�R�L�؏��G"�a�_�[�sf��������^�jZ�g�:ݮ�6}S}z��fv�ew�r�ϩm�J�|NUP�pe�2K�!a��W����h���1Q���(�u?��ҵ�^�Y�Y]�&�t�َ�O���+���H���|�{�1BkdS�AE(S������Ҫ�����q �$�����׍M���&���T0�$�}�cl,F�ǑC\&}!��|���>��)�'�q�J��4�r�#|�a�j��G��I�hIzG�d8�׎��; 0At��_� �����yיd�K"��k��W�S��|.'a������`/6�z�O"�z�C��<�s�S���F��&*�a��S�Ǻ��}��\y*%�m�ޒ,/Yq̟S�/�*�ｙs��m���k��nI/-���������|yڈR9}����$n3��᱑it%�Kj��`T���uxW�V/Z�b��R�u�`��,ş�q�+���1���?&ԕb���4�����1P��n�i)�����Tj��ک�Úg�0���dҭR6�/���9�,U/��!�jg3É��E���#=�@o:����V�A��o��{V[��c)��߫c�hC2lk����/�a�e�����Q�\@�?ە�k�1��7�N~��O�� �n����wd��YzS��~}�u��D>���(ƍy��:�*���rפ��L�c�l{��`3�4�;�ӱE�Sb왷�~7K��6�;�^蛀y(�KU,���JL�L�p�V���/f���0�2��ɶi3�H/��	+�372��:�Q{B�����.��HÒ��f��۽�	Z;���ħ?pW����:����U�Z˰n�ƒ��$&�]UzQ��1�"�*L�ʏ��7�K(%ȋol����u���Q��7%�dKN�ʗ�O/�T�ʘN�L��D�Ng{-n��c�=ۚ?nwqGs���	��t\��.��xk;D��o՘�o�T�zx�:�K	��ua��k�=�@Z��Ǟ�sB,���V�.|S�zʸ],�s�����sT�������%ee�w�?���(�����#���:�]Q�B�$<p-�V
����p�L���o[��"��q��)�d�y�;4=ߵ	�����j�%�h1����3�����9��_����Fk��0�^�s��0{9Wv(��^)^Ld)���rs7�Z2��8N�@��ғA�N�w(1��[�����VJ�?$m������f�����iަ*��r:��۩g��������%;F��2���g��Y*
�����V�|��/��Q?g���~��U��PH7��Y��y>����ץ�����⠤�gH~�7!��
�+�.����f���x�VP�v�����˹�ؗ�u�(0|�nX���u�Я��w�!����>�&7����o����VYZ���m�{c��_�h��1sTp�^Jp%R�h�ؒ�tS�PP������)���Q_v
�Ê��t)V�Id�4ib�]~�T�˓���<u�+R0m��V���#�g�/�e��d/k1EY�7��4�tX>,�K������x���*��Z�"���*�S��q����ŭ���%$my(cn�����#9=ŒX'�7\��!��v~:�s��_qX%��nF���v�0�=1MX�y�@�M��w��Ḍ�0k �JW�) �-6dR���c����B� �P������i*O�1&39�i�8�!���g;|�zj��A��m_�Ӌ���4�h)8��*6/�P,(ޘ�qw�݇�@d��J*.s�wYB��Z����R���]�'sp-K�t5�{W:߿��6��;T�_��i���*OM]�u%�_V9��vAYS�
e|�N�������z�%�����%z1p�sl���^��X��˟���3j�x��j�D~�b���o`�*��\�B |`��;����Ư�ݽ%��aQ{�o�:��Cf#�Q#��`��&Tr8H��ٲv�%�-A�k�;gl�|�ѪD�C�ٷ���\���1$��$��0�_�"Cv��ҹ�M#Nj����f�����[A��9r�n�c��>�^�w�><K,oT�(mG�}�z���5�Ɉ�9��^���j/I��_�������l���k�ԹɄ:��ͅ�j�}�S�(5)A�n^���*�Y���	c��ֲ�V ��Z�l���'@��>��=	���T�	���; 1�f������)в�6�.�X{��T�1���Ϣ��}����^�C�oP�<���X����9�>�pcq�T���H)�A��*١ԫ黉��K��8!՘1\}����pTf�'���1aX[�ya=�i���9�6�i�.�KQ�eX�@+��nr<}�&���3����[9x3i"<�J�v~�eOk��f��d�b��'.b�0��v�^��ɔ�&e���Kl��kj�,X�rV�%}��m�vHT�~��[h�o�u�i�0�P�!Yv�wF.����C0D��c�I��8�Re�.=�٫�w�o���P��s�O�ڝwO�����D-X/%�t�	M�~�ΰ�8{9��*��s�r�nZc�@غ�	�~q)� L9~6 �m�q)�"�4�K��.�l��HK�Y�l�U��X�2m�� qn����t��y��[�~�]�b��]�1�`a��]>8�yw��n�Dکs�SnXL㓈�<+S,y��!�}F��)�z
o+��囕���m���BQ���+���u �-�Ҭ'쏨�f��϶�}⟮��- �����^�b��b\=�#@��B��L�P�¿mtY*>PV0�b���.~gM�2oh#�d3�N���2]M�~=�L��i�qY[6^o����:���ר-��᠛�a���r�Ӗ��Q0k�賬[��¼jUR��È��+�+@=E�15��0D~�~S�=�2	��ˤ5�ſ�^W�D4��k�|�T��z����ךa����ҟUBܖ���Y��?�j ��DO� 1 Q�H4>���c�v���7�5�3S}�i�i�Y�5���> ��� �$�W�x5���h�1���P=ʷQx#;Ϝ[z"#bQߢW�	�H�����F/���I7�Ԅ��1����V������r6����>�����:�.1�H�i���my���vU	��v1D�ct�0Qǃ�>�$[�Ԓ0 x��	o���y������������H՝�����Hb������������S.�9K4@��A���м���遣�@�{�˟��I�����
�̀�W��u���A/���D�b��f,�G�#�cz���M���z�teP��)&�o� �;۱	���a"��c�[�n0��̎�2��US�+{����+4���a�����J(�*c@�cS���ׅ$�Z'����)�f����j��_l'�S/[���,+;�.:�#�0�.EyG��f!��F�;K�r$e}!+�s�q�$��o�A�Ţ���'��7��/�)��Qa+�S��j�k@Px��
�)��q��S���A�k0��hd輒���y���黿)9�k�L�e��V�fU��-l���`dN[�d:F��;ߜ�t
� M�r�$�XY��Ꟊo�Ԫ�@|���O��H�����u����m��	��S�ћE���<3�^ܕ��|j(��raOV���x�>9YxD�]�R��I8̇R�d���>K����Ř�U��A�z�u��J[��=A>�"-=�I%�y�s�}�ۇӣo�����u��x��a��-�E�1A��]>E(�<����l�ţ4��)��6籴!B��d
��桕��JAl߬R�/�;��l"1) �1�M��aT�w��+oʷ~�x��'�A�62�D�u�W̱Z� �ޞ�6`���x=˼�͕�G��a�}����b���&Lk��Q�A�����rj����t?-گ�Hz	�,����;�ǲ�{nP����Y�-��[k��R�GxGqM�(P>�%u���U��&�}ȖH���2��U�;�;�|�e�3H?`v/Ό��wk.���;�����H�̗w�ƺ�>,��G���D��^w�b('�ܢ/�#��)2������L��H�
���{��.��a���Wɫ�I�e��PWzu�o��&�p�6\zHt���d�\�&��6�(S�^�C�c��T?�dg��������O��I69�;�'��=����a�Ň
5�&F]�����\eڳ���*�� ��^���]��d$��S-�K�%`��QP���"d~�ɕFs�Ϲ��D�5Vo_�>C�Zt��]}��hY��d���4�:�u�/�W������rZC�ɿw�	�Ϩ��qSTT������h�|�aq}���*|�=���;l6
� ��{��\\[�1�d�DY=`���?��'u�F�/�c����R��-���]^�M|g֫���K�lAh�~���2
ݦdQd-�˨�S�A0�0�e]A��d�e
�̸ҩ�P�йH�k�MsX���:._�(�E^���".ܼ(�p��5�D�(�����y��Ej�� -�␚D���f��,%#֎(�d��b��ģc����]�n��J�fs.����2-�hH�/�7*O�"i�<~��Lj�ѐ0���,Bgl�/���UG��L�i���m�f_�F}�0��0�Tx�R;���Zg��[�mϧy�&���	u�~����2�%<Y��h��wq���j�/\�'puU���;��k�OlQ���i�L擊v�~��7;�ח���l��4�h�Q�<��޸?�5�o"�ȃڄ"�`%F0�?w(g�xB䂍�4!*q݆jz�K� r"�W+3 ��U�m����JUp\V�/ȆC�$��;�.�vTQR|)S��m�N���4iS�V�ÛP=R|��|H8
�Q��VDb�R3�^Vs��^u�:�I�	R�|��p��О���u���r?j�~-]��g_Q�e�ިF6`�i����v�4�5~���P0/���:e�.�M��=z���D�z��[���8�OfmR� b�<�j��W�e9J�>�P=;�?����~�E$��p:sz�.�[��@0%��>D�D�h���?c8j�%��̍�|��;X��(�E4�H:t����?���gC�<c�ƛ<q���P���2W��[D�����OMz��ʁxx~~T�6-�0�SQ��-,Ŷu�웧�a�O��[��Xm7�q�"z &s���.�z�-����Q�����.Oy���X������W�y0ѹ�Z"�Qq!�`\�RE��lƪ5�oh��f�����,��O�ױ+��.��a���[꜁Ahv�Xz2Xim���{��-�p�F{��H� ��aA�_��OY��ݎ�>�~�����yy�]��B���+pe�$]��]W��i��u�.�����1��u;���ٹJ�L����ȳ���6�[���ү$1���B��b��{����~�c2&68��8��}��U�X�qg���d�}���Xͅ��|���@�?j/X�9�l��\]K�ɽ��x��OM��قp_Rݫ�a
�ڝ��;��R�M����^�Z����ϩ���B,�T] ��_�4��/J��t����ؚ�Yx�z��	/'���|>�aCq��Ρ��;]G#ύ��6e��o,�bTÒ���"8�.`�_�@Qˍ��1��(��Z��c6�e�N���I��#�e�bm�w�k���״�0�RhJ��ˊPQ9��sCK�!��da��H�X�};�Q���[�ìH1��{R�U#�Nf
ί�a�p���F��t)<�6���0��n��"x�jV��d�a�=�d�z��C�S,�覣�D�a����J�=5�Wl�K���o�������u]eu��c��`w�n� w����w�"�͐��k�� �g|X3���K�QA(������;�a������I�S�1��X��R�׃��$Q6����V�R�B�oV�)v���<u
}��b�87G�J��
䗔M����&��>�6�B6��<�m�:�*&^ krP�����_�f_��e��1k<�x$�pA�ڃ���J�ʈh)5׺��G��(c��RS(G���,H;s���JY�e���T(��R[�H�.8�]�F�.o"�!/P-꯹������.�Eq~�S��l�	1��0uQ:r�<XK�S-���>��ʒ�������W��:����QKA���u����# .h���U���d��� �5v\U ���k1@N�����{��|�A$.���ٜ�/��x��hݴ�}��3erT�֛�t�=5���.�q�ӓ����������N�����;���v�ϺA�8D�%oE��!�_�N/l
�[l�,����v#*5��29l�M���ZM
�iQ$�􂫯� vFX;W���?���D?� �Hxss%�A�0߳7d��y��O]u�>C�67t�_S�A%-��}��g2!�G[�mJ��
u���C�΍(h^������ �{
|
-�w�Q��7�"��*��E1 e�Aq�����;;���Y��2��!�u�Bfd�k����@zS�=�E?�㗖�l��`g����Y�Tj�ܪ�L�5���ᰃ��׶�k�'��5|���)|��<��2䪤��{NHA~�+�z�����c���u���<}����Tw'���*3�4{���eKxY�z�$а�3J��B�]w�@5�Q��'I���v;N��_��W�;����u�O�x�����b�LF= 43���2�jjv�Z�¨C�RX�u�1I6�<�3K��4p�e���)z&K����F��~rӗ�@T����k���|s�m����=���W<l�2�Sf������~��KSz��"�a�*�:J�L� n)�l��f?B��^.�\��&ʪ{���91Ѧ��ԺbH�!nGO��X.ݢ��C������"p�>p
<t`�0��p~���:�s�a�Fo������hËp������;��E!wա}�zncz�=6yA�%��qˏ�n�cup�Wh��B�)�]ȧ��ꢶH%EǬ���������נc����	o���x�ڜD�ua��f���n���Q���fj����o�~^m��Y�0
�o�G��f�q�Pv0�x�|��rS�ah1��c�s��XT��	[A<��B�'YJN��|L�Ԁ@j�"d�l�_F}޳�!z�2h�у�ͺ����7c+ӌ�G�ƟݝF�*ß������,q�V�&�L��"�����܋�JBoYF�e�uG������}����u��:�;������c�Q�����mد��_�eO� ��#n�t��FN�O��F� �k��H�z{�:B��i+w9�U�P-�qƵ7ݬ1O�΋�)�-Hxv�r���mX�M���Yڨ^�_��,�EMg+��1����%�_���ڜ�)%�^7>NZ�}�pG�� 
j��|��,�fkC#�"�V{�h����6Qn�~�� ��K{3k���m�� �7��5�"5��O�'ԙ�h�r�EpO���IK��imUyX���R渾���9�N]�!��m*|���d}4?�:�?�hy8��h��n۪ߖБ�j�eD���/�i��EǦK�+���Y0@ڊmz%_9��Ě�։�մ��𛮜�>n�0P3

�-a�7�B��6(�q�F�W 	�C#K��d�c�n�+ڒO��p��m�4�$��h�ӹ����n�[hdR�[�ܗ�_��a\v�~���WA�,���a+����X�o�h$A
�74i)pw���,m��A�9���;Ӌ�ŉv��|`�A�g�R@U�?��O������@y���u�f6�j�(>f�������}
6�0�o�x����r���f��f����|ެAƱw+$�J����ɤSM�[�*ߨ�ɱ,M=��p��|�k��)�ׅ���p�e�}U���ߟ��Yͣ#�S�
7.�������i~E����)�p��vxm1���x-����C��i{�{�� ߻B�Z@���D�E����G����|��4v��lDӛ���l�E�)�!��� ����=�������Mϔ.�	@�c H �q- �Ѭ���74�4l���ra��ڳ�$���w��Y�B����L�5bփ����c��ZL|�~��7J]��/�Hcdθ� Z�*�ʉ8�<ךQ��k���� ˷�y��s�(�f��5gJ ������>��c��ja"��FY�P�JF00����,>>
��g?����-se9.�~�'�s��'�|�CӋmÜV��=I�U�?��U8��*@��+x<������eP��-���gjY(L�>Í ���F��|n�" y]}m*�z'P0Vmy`d�Ok�%���p �Fu��0	5�S�]���\c�f�V ���j��m�T�*s���Zs\��(�t�0���0>����b�%s��{���;�1�#�㦵��tL�kD�n$�i�`ډ�6��͗���d�	�k%�=��I� �͞��:!��MRM��֬֩��$t��<$Á��O�d k�u���rY�k����� %]%<�g3�Z~��'��{��W����9X��'�����=A��0���XPV��R�&Ă�?�B�����eI�y����߼>�m����M�����Fx`������e=m9)�k&P��6���
4>�/�-#j��hØ�5w֊���j%X(��}!CT��{+r�#�e��m���u��?��ߞ>�V.c��|e�ZJ�I��g����g�����*��hx� A��t,C�Ǣ �O2��`N�o= ��h�&ZT��ºB�� ����eM;O�U� @��U�ϵ �G�����nZ9~��T�ڠ��fAk��3p衇��N>��>ЬP�l�y'� �Iu)���Џϴ	�g=HW��� �����^B����"Je[��Lx���g�-�(k��ѝ�e�Z�tY,$G�b�����e�3.�ÍFH�#�	�-�$l��ʢ0sse����V�rq���c��ZqK<?>��3�ϭ����O�}٥@jN��ቮ�g��zjo
���T\�3CWPj��o����5���f���į�`7�9��4 �}Q� ����B=8�g"�u#hn�y�G�Y�^�T�踇�����+��}�=i^A���Cv��8���?��p�Ù� K��;�Ѣ�+���k�B��=�Vb����:����<�w�v�n�_,��5в�Ʈ���A۴�M��߱f[�Iw�'on��^��f= `�9�g��@@
4�'��@;iB;��/�;��̍u���o�֞� ��@|	�F��y��X�!�����ε�]�1�HX+n�g�f�C����} ��#	x<ki�s�B �3˿�=�yiV�${�b	Li3c�������4X��d-���\��9U�����	R9ui����EC��<�9%���Z��1kkEMȬ3���RUp�Ĥ'i�CР0�wi1.���e�Ô.A��TƤ~�����8y�O��E]n�d$�iv���i�C��X'��c�g?�����BX�Z2����0x�ߩ�iɠ��e  �u��g���p�~�S�W�L<A�\���]�kB����w�*�9��Y�G�>טU0:��녿O���*haX^�i\��{�v��gN�F����1�m��=�L�m��t���W\��?��_��� С}B�c	��`��'˫����omu	����Ȁ<b�`q���lC�9�|��]�oOJ@`��bG��m��'C 0\�Ղ���{ܟI�ř9���q�|<��/��-�V�
@ Y������cj{J��z�����6`��6�G�!4��	�כ��DÄ�zs�?��?�,)-�[�Sџ8W)���{����0���f�j{ӛ&	�Iց� h���3�DW��<�oj�5�aë��B�o��yڸ6�l��Zk�uK�H���VJT����a�~�s�=�b0s����X
��L�@k �� A�#�4X�t?������@Т�ǯJg����& �b�p6mo�M7m-��$(�뺹����#@��!2:��6A����Dp#ص�*8����Z����=�����ͪD�?� ~����:$%��'��O�#
$����������ݶ��wS�$�\�J ^�d���-WoBڤ�4�������ƛ����t�]3�����s�ɀF�� �(�߈U❩�p����� &$``�X
^����d1��)U��;V�������B�}�E����M2bj��߿����>��ϗ窀��Z�ȚY9��1=>1Ls���`:2�I��$mc�]�o:�.f؞�T�u��f���N��CX���k��@��x�^s�e��_�;��=��B@��jS�<���gc�]�6lZ���$`�a���|Ң2~, �I�c3-��*�RΉJ�.�Dy6c5���TT�>�n�&X��u-�.���k¤���i�M�\�Z]k0}f�X�������VM�~�ӟj�c�����vh�����6z��ײ  j"[����G�	 �Ɵ貐�cU`��<�E�$��X����J�I��u_�m���,O�x���������֔_>)�F,��
@�,��R���b�z���0���x �x��9�\�=2�0�(ʢN���������/-��;��(M`�F|A��Ϋ���J���L�Xf�M��e�T��yf��ɥ�Lk}��;Q|�(�O�]_��Q�h��� �������'�{�V�Sp:������g��I1��2 ��64�3�! вo��1�d=�Z�APh��3����6�R�}�L�(�˂��Y@���N��i.�y���TA������5J�,A�d0h��j�gN5�lH�n�g3.�B[ǗOA!^T�v n��{���VZy��\@/��%��
���`���!��l��&��?nmay��3�L�8�<3txw��:�}ߟ`�#�"9s�1�[�0֤��;��(��dͨ�L�͈ѣ_�����a� 	�iQ�YT�����x�K^�,��e!N�X�W���Y��d�c����#ZYcZ���?�f>�B����{o�o󛂃���y&�y(8Ԓ'�7���09�;���`��g���'� !�0P�)��˳ό���s7�{��CEYH��I����E�P3���ԴTA.�����]_5AsJ��\�9��~ӥQ#��^S�oZ
��/4'��I�uI���6��A�`Ư� %}M��=)��pi�݉+�x��G�=�Ѯ��:��\ݏVNf�@��H�B"��ذ�T}�V�R�+��b�Nd%��sF��~Z�j֝����?,�F��!�b�(v�T����U4	�]c��9	�k�p�Tt�N )YǿN9�&�����ǹ�D�J@ AcR�b
����EQ�a���Y�"�j1�QieE�㒞�����Ԓ��ީ�(��)0�@�ފ	�zd4�''�j���V��_S�&iz��j�da�Ԏ����o�a*X�R���Mzv5�j��oJ{���Z=�U��Y҆�����`;R/�O=�a��e�c�2�T�V��ұ�W@��Bs=��4�.5���X�p(p�4e���Yw�鬏�����դ�A�^�pmk��#ƣ�9��PY���Q���d��另��3)�FO��
�!�Y������f�mFw��n����k�B!�q*"�x��O���� ����gp� �'U�V
bRD�i��K��mY ������}�;�|�� f#8��[�2	W�T���O�����:��~O�)��_X7��(��S�ӉQ{I,k���Lt�4��Q9�_3�;1��
�R�1%Ɠ�0��q/��}n����D�?),��z�\��ޯ%G�h@�ōux���¤v
C_Y��F}��[� ��̳�xsB�)�xk\�w�it(T�;mz���8�����}�M�E;�#6U�l	c���9>[!:2yo�jƦ�������J��U�����?���M��x��$�@��� }��ʵ>�Э��am���}�=�l=�E�Z��ht�-�؄4�X]��~���*�����2ʴMQ(��<c��=�Oi� z�L4z��_,� u1ָ�/��ŏ��g���;l���	X3 .X7�*ip�T`P�M�,�u�~��hYr~�w��M�g^�����IO|kb&�.�����X��y�R�7��̓!��L��L�>U�M�q��\ jl~��\�qe�S>�������94�+s�a�{&�������H��Q���סL2W-~8l5��m�#��Ƭ��20��,�me�$Е�o���g�Ս�֚k�X�ƛ �T��g���븆�z ���) �j�2o��ZO��������5'����!p�|?0k��g��\T:3�����:W�K�ꂀE���$��qꎩ�H`4\CP7�u��uZ�2Z��[�̜��凃���1���G��f�̙� ���S&�� t��
A�����p
"���8� 0A�B+�!h�~1/��9�,���=�*`r��d��*��Yi͵�ya��Y����&( [a��0�������O~v���,����d1<*&�W��$�`X<�Q��*H��Ȥ�`M[L��ω���^��W�<��,��&rt..�e�OYw+�a>4��ό����Fh�0���4xU�e�6o) PU&��i@`՘��� A5��fX��?{H	7��oEQ�6�y�)޴`K��h�G6�y���I�2cc�4�
��m�au1���yP+7�:���3|�T5H�x�r�}ՂB{1)��ĸ���8 ���֟BO�G�"��&b�?̙�k����3W3� _r�S�_�/�w��6�f�<Zx�����5 @ib�	�����1kF!=��A�I.�2u�0Z�ygLưq� @Э��5Ƙ����񥗿����K�\& D�|DRJ�-}'& FC6&S�J�P�iZ�1��ͱ(`�pQ�&Ő��~���=����hBsnB�����'f�-��uHRWԮYG���P`ɘ���[
djh2W��T5�V�1C@P���� ��%�1��B@��F`�%�~����u��h��q?|��]�[�	 ����}�@�� ������jR��U8)�	���&�Z�����I�r�^����V]�̏�9�Re� Xp`� z�C�.�HI}������z���7���]ceBxb� @` �7��
VT�8]�Ҝ�X3ıU �ܹ6��N�Zy���U�ö�%�%�mϬVh��.9�t�"e�伿�ۿ}~�w�5��� t��D��&�߉�`�5`0����h������PF��%��P/OJ��_�◼n�{�~�\��ޟ�C��3w���>����t�0��eT��_�h�}e�UOa�U���a`�ؘ�-3�ڵA����]��FS+m۾LS;���s�k]�j�E�r�:�x�L�
ȡ��n �(�}�����*tc4˸�!��O��|�9�*� �����u�,��"�xU04Ԃ'�(0��y�k��J��k�yҥ
 @ӧ� Z:���Õ �Łtg�uV���Ŵ�wh�����g�*�Ј偀E^d >�<�̶ΘG�CU��y�ۤ�9-����16�x��x�+���)��h5�7��:���Ě����X~P�ӟ���>�y.u���%����^�ʹ#�-��^��@jL��`���-��o�}АqL�?|�s�󦔬<:Ϛ���_�(��A)���0�{g�m�zd}*(* ]� ���=�����a#�S)0쓂dh5����,�U��:c�EZ_S�{���g���M�^�@����!h��a�� <O����CF �7��&U����Ҝ����V!ﶩ�C���h�T�k���i$8�ٕVC3z�o�~������M�?.)0-	H� �9C���Y�!�XXZe7��<p��>�^*r-i�<�L��uf8�I aҘx�����;+� �R6�@bMV@f-�$'Cf��o��!�#� ��y	�|�\b�˔�@�f�<*�j�2����J 
�s�j����	��	Y���)�{ Y(�O��b�����ͥ��}�[H:�F�>&��ƶSz��e2n��I�bh!p�_e�C!�4�qd���7���4I���#����*��n�OZ%؇<W-掀�eji��������=� �WXM��4f�k$?�5_��;q�&H�����%n�ц�c�b�v'C�q3	oij���o����*ȫ`D�S���}�Y �,x��#����<�ﾣ��߿r�5��d�f@3N�ٖ1@\�J��:��o�vt2�W���Z�gLƠw��59ܣ����8�B���y~2rƩ�+�XRKU0��8��F��g)p=��un�_]<��k��^�Wk���<s�L�PpP�����VO��������I]���MTMg���,��{{H"��������?��o����s`^{�0�E��M��u�_��T>�� �$�<pPҰ�e0�Z�����=2��dkd�
X�{�=���FV �X��6��M�0�����;��V+���	�L����� pp/{�	��-����8�O h�������k�ua�G����۹�o�&��>�w�g��5'�z�b��� >d.� �� 'i���i�Z}���
 !,p�x�!��z���'�᚟��lM͵��`9�h$&������`~b�8K�5�z�eV%�!��=1e���ꜳ�W�ׇ�
�Zf>����s��9�p�L�j�F���	-c����@3*�V��HX�BO|�ߒ�O{S���:&P r�d�<�2���K����Ф+�V�I��U?�A��1��ʸ����ys����B\�ÞQ��� }@�@c}t��}h�� 1}���a����^�b�x�Z��#�iUT�y�����jX�,h�kȋ(��ʊs͢���CkI�KMU�B�k� N k��6�l�f1 @'1�SmPZA�-�eD����n��=�����
�#:�A00�Z3���\����	�O�`F���^dlĽ�]��w���/Պ!m�Ͷ��7�tz��	K{��e.���җ������ߔ�%�9�i@ =cn�G���)��l��eBL�H�	�T���R�!�M>d�aTY�JD��S|�98d�V�Zk�?r�S�C̢q6B*��5�6g�_Ô 3}J+T��7�L�7	X����t���Ȫ�`8�m*h'�����S`{?� �h@���yDF[hq<�v+���ސ���j��S�=����z�Ǜl�I���eB��	Y�n��W������>S�C6Z-��w�X���.,l��5(REI0D ����"π�^
���'�E�\��&Y+��&�Y;���,��;��K��鳯y��_��V�q��O��h��믟��Va�=�l�����z��=m	��������?05~�0�/�ߗy@ 㳺�G>���tH&x�v0I*�qb/I͕֬�Ƣ�y��S��aq1Ѽ�|tmRe����A�_[ٟ�tS ���q#<9���wռ���`�j�;9�I5�?5��4�6�3(�Bm����u�F�o2V�A�
�j���n�媠����(j���4s1�Rs5�����p��c��Wզ �uŨ���Lhz�����k=># Ѐ�����ըi^�P��[r�� �8��!�i�sk�>Gӷ�u����yh��nC���,�o����\�%26,�?��G�����ִ�r�t����?�,Вvi˂J�6� 8v�
-�w-=
ߺ)[���~�i�']�9Hj#�������w��9$��5�K���
�f/<�	Ox������n� Bg᭓�^�bO�&tg���d}F,A�~Eѵ��?D�hQ.N�y��s��Ї>���zֳ�����0�s�q!���'��W����]�=�I) d�
l�B�
)��TSk�{a�����}�)wh���� TP�5C�>�6n��-�X�t-���;6�5��,����
�+�j𚧡��n�&n<��7c �9^�jq��i	���T�7�-�.8�3���Z��N�7�H�?��ܮe��ӵb��t�8��J`���s�վT��;7�e��3�s�ڄ�i*��� ��K@�w\ �A��vMV\zɥ9������z����!��j)���n<�˺.L�[�� ���u��?`��%͝R>���
S�$�fs_ճ� �	a�e�]$��Ȥ�\W�NU�a�,c`���ǅp��~��/L���sj��>��7	�_�(���/�zr��p��>��؀�n��u��*j�6=d��GVF[M�2P�C� ����at�9AA}N�F+hђ��D8�f��Mb���j��^+��?��KP ����T�� �]�
^a�]
j�jz�m�\�O�+}}���j��7]�<��z�Cն2�� H���SSk�u�n�Ƭ4�M���M�`���׀ ���]w��%-�֎��D��ג�<[ @@�J9w~�j<?���M2��6�q�{��F��}���2�Fz׻�5z�#ji� ��Q�����	���ޭ��}���nQ v�_���_���n ���^��?	�(��<7pO����OB��J_{͵S)$���|�|/�42�M@�UW^�j��W�K�+A5�JQ��&#��E=���e�9��/�S��Ĝ��d%��6+#�g�$oxm�
��5
f
Z0�pPOT���I}s?i��^���
_��<�=J?�K��I�G�p.u�3����V���36�
�hg��E]����
�1
�ٮh�<��R��f��\��*�g��z�LV�^�_�s-�km:�7�Zw*(`N��+��r��3h�*e�0����&�>��������R�!�>���x�����}*���K>i�я|dţ?o=��O���L��!�8���H�J0�ܜ_D�f1�OSIU�sl����(D�X�	�'ʣZ�;^m��nrP��G��D{����D�b-��L���+~s*|}*֊�Ѱz3� v�e��3��Z�j������������ɪ��3 qA�2�;L�Z��5���ı��OX��߾0�� �i�D�3@N��� ����C�BNMt�U+@+��N7�����L.�0��D[֖�Tmu� �Z�V�I�q�3C����>j%���*�k�����þ5�մ�TA\�X���
꺪}T���V��rk��V�����f�`�����O��
��W^~����n�z��G�>��Ѯ��}�ʊ��.��љ?���#?1:�������������E����.�w�誕�5�]����AS��\I'���%1D�e��0�^B�ە���8���K��?&-���<2�X��z�"��s��SG����p��&���C��I8߭���]����W��I9�_N{w����Kh�/-��Z�^"�OM�w�9�'���na��4d}�W^�p���ʨ�&7Ɍ̞���u��J��ڟi�jH�d-ì�ǡ+�C�x���8n�b�CPR���x��y�������e�V�j��3@� ��7� MW����9�~�	���L��Fuɨ��V��	"k{��]�#}����@�߆���3'����q��Z��?�ƹe~ ��
��P4�P,���b��5W���.�=�!�]�[�7�4�臿9s���9��g�0Zu�F�?����z���)�L��@\qm��^5�X���<������` ��6H�,�=�dI��- ��)�qv�K�uj��|JLJ���V���F�BӏkPU�(.Zc�l�i��Y,�p�:���4�'��m�txt�m/\��?{nS �Ï'S�[�l=>V�'dm�=�|u5\֚V�[2�j��Wf�@q�����ι'_\�?{F�� e���n�QM�z�2UiY�B���jm
H�����Uv�����
r5o��_���KM��Y�i;C�2�4����;i�'i�|g��
[AΤ6d�%k���3��@0@�8d̯֜���Ļ��2Vn�咋Z��g<��Gw�z�\6t������G��4�ˮ�7�߁ͻ���&�o::�'g�8�v��j�!�9W������6�]d��I��s��#o��aR����]	�����)�&�������9��a�˵Am  }�������
��l|������yg�y�w$�z���������+�f��=���E<���2F�$�����@�����Ԭ�gm�- u�OպaH�T;$Ee�0�ژt��,��e�_��9�he�D�����.j�C�2I;����+��[�Qm[Ư���ԥ�J�T���>jm����G+.�h��� ph&�dIpN���:�*|&i�Cp!Mk�|�xT��?i+�.�mx�´�:���K�֯}��V<I���=�\�����5VͿ&1a������>���%W^2��[�毸�����p���sMN=]r�%�k92qk�����K.�G4!+��#2Z�!fxi�@��v
��eI��۵����;-&��^�/c�}r��� 4��r�S�-XP��\tnJ�0�k��W�0iq�k�������T���oz��x�?���?/�џ?�)�٧f��C2f���ccm�'�g3���$3p����3���f L�v<�Pp04#׽`eړ4�*L�Y���z��Ma^��=<�=�^5O}��־�,���V>��B^��@�i!46w�l�Ң�����5֟:�3ͽ����J�M��b���I@���b ���t}��-�EV�N}���஌���.�����#?}��w����;~���:Z���G�E�_2/�^�L�uW[uta�>�Ol��5Ȳ�6�[\q�he���̂d,�Bh���8�_����?)R����#耠�R�aj�Ρ?�9/�"�	g���WN��<�4ʦ�9X�B��E7D�0���@;�#�_v����=�8�ē���7���a_�u���bb<K�c�^)�T	����ᓲ��%BVM�u��e����
���F�i]�(Ht	(�41�~�����y�n5�L�|R�y
*�h�C�P�F"�U��x�5��>�W�Ҵj���:پƚk4I��A-U+��U���͌�u��r��n�b��>�9\�U!�v�d��XY��0˥��J�8i]���\A���χv��������M�
Z���7e5���o���O���.I'\-k���:nt�UW�V�����$J|�5`9�?������Z�:�$� ^�$^�`�;l|�v�U��"-�Ǯ����_��5�H�Ж9Fz�\uʒ�G(�uM߇���P�ha��翊&�UXx���ḶN��+�,X78�k�b`�n3�|����~v��^��=>���}�?���R��lƙmOKj����
�*&g��1n����/>:�����m��r0rR�X�
��� K���,X`�
�����Q�d��o$�)o2���$�@V�U�2���7���7ϯ������ WK�>۱��i�j�F����(�R�َ� j��LT�?��gr%T 7Ip/hW@XA�� �V�O�y�C�8��a;uXW Ig��dy2�Cz�)�1̴sy�F䫯��h��J��a�G���9��.	_.�}*XF�����#-q�h�����W_5Z%�d��i�6����>��$&��so�ƚ٧.I�����"��t��J���� w������,j����L~����X�|��0��m�����v衇~4E/�7���$J�ܧ@���^�i9��۟��'��w��;��4���$+�Zhe̕��[�I���b8�6�!�"Ȩ�l(����0Ts4�`>�S�û{�� �6I���o`��Dc\1B��m�V�4�iZP?��
X,�S��
�$�3Z���x�]:)�����d5��W�=��d]�~�b�����\ӱ�Ԑ|y>�?%3�j�^�R�dU,g�]1���F������;l0Z� ��Sѐ3o8x�U׌�8�ף����h�-�4:�q�����'�~z�Y�kr��9��@SP���(0�f$w��b���Kf;I��@�m�������j���}fҽ���*h?�D��&�PY��d&2��
��)�|kNQK��$�q��N;�^)N���l�zfƭ��~��F�Xp3����X��җ����"wc\�@�*�"U���Q�ȼ�fj~��z
h��Y��܊u��W7���£Z.&}��'ȩ}�;���y]��5U�Nj�
�*p+�P��,nŌ��?�8P]wu|d"�W�ǵW�_1i� L���zv3Y�*��ka��E�n ���O���@R�6�c&�=-3ί1�+��;����k��ų�5>)���q�M�U�-|�bpEJ_7o�d���o8Zc�UG���w�y�X.V������]9:�w�$�`4zի�u�=�=�;'��N=���u�P� 0������N�ؖO�W]�<���P?�t^.�X�?N��' �1Y�[��x�z�x|�մ��jn7�LŅ�;�� ��f�v���<gל���A�o�x���$M�ܧ@���8�|�O~��Sk�I�=8Lu�0界�W�M�3	���O25�N�fo�<7A\ ��/��itC��l)\����4��
X��PsU��m�{ ��t̪��P�qp~�
f�i}V; �	籽��أ 0 ������'�����-���$�Xw�f��  ��@�XP���˵���"ԧ��������<W�뵬�B���G;��(��v�2'+V�TC['�TƤ �U��*���ο�B�sr���^<Z9��|ΟF���h�8V]a��&���%�]�bX��W�5���.��'S}�r�!�[�qc�rW�ZpF�r~�ώ��1��"�-�l�;��A���j@�p+s���A�U3�ڐg�%/M���x��r�Ƨ��~.�,���zَ;�ȡZ����㒦�$��v���*��V�V V&^M畖��N^�+��]�f۰O�e�A����a�������&�}r��6@C��fcz��?h\[�{uW@�����<����
�0��y B��52&i��X]C�������a�C� KB��I�|Wiq������\�ߢ�@ |�G��R�N&�o�NSU/�v-gBPI0�P-v�T�0k�`ݰ�v�m���������~{�{�;�������qT+�r��*��� �^)֙<gݵ�m�ܝG���9�_��7�\5���VXc�?��jS��x]��qUiW�w�	u�x�y� 0�i�K4^���!)�@)+�Θ�������p�W��Z�.e�Uӕ��a:��� dzj,2`�^�G��M����{��|���ߑs�O�C��N)p��~=>T\_���ON\ʎYS���X��C#�V�*T���l��uWS~��)t|W�f5i]<ד�0�jj�X�>i���i�&��h�
v�c?-3l��+������ �7���mNʕ&�L`A���ŎE���� ���kx����gC�3IS�`��N��T��}T��μ�W=D����6�4�)���l(!�M��kc)���I����2�:sv2м)ǝ��ٟ-�P�ˍRɳ����غ�8�ˬ}�b��i0�pC `�'����u�;�c������H�-�6�,\���4�}_9Y ���x��n*ק�`�z�xNoH: X�xt���jJM�*>�'��ܞX&.�|�`erf!�3P��4�fN���6`l����_��_'�p� �wr�!��,��W���H��p}4P��꜇<%kl묻5բXg�@����\��8�5�#�@��8V6%��Ϣ��<��/�m�xl���ׂ�X��4���U����Ղkܿ�n�(+h񷪹�-���$:����pK�f��Ⱦ���'<���9�ʵ���;����?�"�?���������CT<��d]\7�b�;���G�r:h���>K�@�Z&��fv�1)��[' �~̻z^�z����7��̣Ѫ�:�W>_v���S�=��j�$�k��������E��^�BpI�J���b{�N;�tr���s|��k�j2Y�="U&Rͱ"F7��$��c&[.t�7��M��Zp�'��s��N���T;<'����>>k���?,@vۤڮȺShU��$Ͳ��'�o(���h��� m���/x���m�X�� V4���$��K��u�Tp (���u̱����U}�ҫ�C���*���jڼ+�<����3�pM|�&/b
TB9��T~�ıTZ-��P-
� ��}���J��ේ������R�ʖ)�C %�����0��	XHV7�v~ƻ�f��8���QܸS����ʌ�;�Q\���?��L���\S�����u|�o�eo�u�nc,������+��d�]��tb�r��޸����g1b�;6��n�&���������gs��j�4�������n�Z�U�m�8�o��O?��������1	:|k:\��b�������Da�Fz\f�a_�e���le��>��Э����o� �K�M}�|�1�����D�c�֕��Y��`&��a�U��W�"��yW(D�V���>�
!��v�@[�`��лZ
�CbCz7�4�G�O�ڴka���P�A5�W pK�_u�Tˍsw B���\�/O���3�S�8֐8"\Wo�M*�N�)�4��g��8`t����,<2֮Q@�(%��f���
�� �qUA,o��
@�&	Ndl��ӧY�ν����f���Д���u��)�zu�" |ɯ�._�����0��3�k�@C"�W���(���AL#s���A�)�.�ʡZ�`���N���&Eq���ߙ��υqR�n�W��r�r�n��71G)����R*�}'�ُI��S����6@R8�֒���j�%��]� � /�$M{��Z��7��`�Z3���u{���
ɺ�?�?V�T��Au	H˱0��x�{_�T�7U�)���>��[�o�^T�D�ׅ�o���TK�t�5��� ����&����X���؀��) � �tY��:|���{���A	��^{$po��ҫF���Ì���q-#ᚴ�?�a�e�����]�f����2������O�n��c� +�T��>`-����cYp}��
K���""}�'vď��r�QG==i^��ww�Z��E���z"T�L`��Pּ>�c�(�n)�Y��ڪg�s����z6�/�˷J|��a���|��;���_�������ļ�C\{������7����n[�|Ͻ��^��1'���Y'�g������Hz����e<xMk�-@�F"M��q��$3�/�2m,k���x0�9���Wm<�]�}a�'�P�)�
K��V;���- Ѣ���P<h}�_�_�$ �v[]5`��:L��(!�*�xnX���[�]::
�!P��I4Ԛ!�q���;p�%i�+����)H�Xe��F+���!CY?��|�kG���������F��h��6���:>������wG?;�W��O;#����.8�r>����j%�3t#MA��^���F��G��3��uo���1��SY��X�\3����q��2,������|�z\r�1��=;���zz�����[��ʤܰ�����bA��Q�	'i�4�|5-�pj7F\�c��]sD����g�i�����u��O9�=ӿ�r��y^�[��)&ڋ�z׻�8���'X� �~�"^KCs�r�y�?I��oy�OJ��e�47���2i°��7dj�u̆���&�̊�d%���?4��Jh��8-l�s�
P��F]A�Ev<�[���
�I��n��yp~7�|}ִ B m@�����J�*4�*��k�
e�a�0���p���9�����?�8> |ƻ��&dw�i��3���і[�it�uW%��ף�O��������KF{�y�v�C��G��
P�|:�u6c�
� �9d�G<��
���c |��p�wZj��-��em]Ϳ����nʆiR\�#)(��w���/>�����t��a,��5U�r�F\kUÐ���?]�#�Lr\&v���|�k^s�h��g�l������??�&� t�^��_�c�= �щ�x]�q�yz�K��}B,?�Z88�'����$7�Q�����U���4���L�����>�]�ߘu�ƭ�[��m��C@`��s
6��L2�W��
N��0R�]M[�?Tt�kŠ5�Zo�P��4ǟ�$0�Ϝ$܆��p��-�ؘ�)��5I3]�	���/��
)���c��A�ں�~���妣�r�E�qtڙǧ&�ى�?�t�uFo�n���'�Ϡ��׃�?�-���gcub]���K�C�Lǥ�&���~�(J_8���96�����1�#JY�5��%���6$���oz�i=#��'�q�c�5�Z�E�q�l~���,4���L�ЦͶE�2�`�dCn����9��oH���|�D��V
z<��/~��/}�K�y�ӟ��D�~��7=G)&xU��� ��}��TNzr ��ôV�iZ�H&,�_��a����`���<$�?3��B��&f���Ǫ w_��!���\A]�Lë���Px��
�}�Y
�jƯm�~���*M	&��0+���J�j�A�UWk�}b�D�_r��M��(�5VZm4?���S!���_�9� ��W_ct������|t�e����u���h��W�A�$����^we時G(J7��_м ]'\˘X_�X[���o�x�3Fq��5m�����\3&Ϫ�k�Z�k4+�1�ߙ��sI�6��K���mL�q���o��T|v�aL�НXl~MMVMH-ւ�20�X�Cpp�'̱����K��Q����0w��Z�98ѿwL����Rp�7��2�H4�~��m�^�b���N�ޘ��oQ�0k���ӻg���PۮL�
���
�J���0d]cC��ܛÿc&����
m��?|A���jA�A�����WM�2�I. ���[���{���0����
3�A�FGR�<yp@p�m�R���T���|j�p�C�"O��1W\�ƚ�� �&��Kf��@��|&L�4JN\m5�
W��=���˯��h��s^̼h�W&�*���ȁDg��� �1��	��r��,�-o���f>ﴉ���t�`uѢ+/M\�kꏭ"�1�����r���RB�Ԡ��砤CSz�)1��;��b�,*��iQ.,�n��s�-�8�����b��a����VW�#F��r�j�����}�����>�a�b4�����������Z?�]?P�?k�9t���v
��o)k�0u�NX5�t���֞U���{��5����7�A�Z���sZb�uO͸3Q����S������g5}��V��q��
\j{�G����D�A�5ر��±�7!�ﾘ�&�*���:��� ZW��P]5���r�����9zD�!�S�q�=�.�UW_��S�z��.������]2����G	H*�j�u��"qݰ�h���]�<��Xڧ,!���#0x1F�`]���Ru�Q��˘��ŘXk�Ě�*=tm=����S��!6�4un���b{~��!�7���n!���5Ҙ`?����M��S���,����r,6Nc4�4D����4��o<��ͯ����bfʈ��*m�	x��/���,5��	����L_�̅{$
}���g�]v9y��7��Q 5㿑��?L���s���nw�Z"F�&��My-ХI�5|s�]kz�U���b1`mk-T��_��������>����5+Ap�5n���#�[�gZ;����[�-���dA���L��'~��V������Zȱ�S}�|�T��)A>��i}����J��>%�W^{t�E�\6�h�MFW\z�4�#c!�aaCn<��VX�}$8��䡀J�1y�',z��%��Ue&K���j�	ݗ��F���.�E�[l��/���L��_'����\oHK�7�ki>dϰIt�YȜ��Q�$�S (��a*0̤%��vFӦ�(�OB�j g�j�Ǎ`��d/�������F�l�~��)�[��������#��%3��_����y�hN��n���dӬ[5�[2Vک~n�`�hun��M�w��`�m�ϟ�qW���_K��8k��|���U[���K�S}�
f��}�������a[��W�����6V@�6LrG�d��Yu�X?������a��������aNS` �Q�A�9�\r��̐�WϏ��d�b���EX_tU\
�����K�@��,� �B!#�-�f��� ���ik-k!��--��i@�����U�O�j��; �%�`Y�g�v�a,/�ַ�u\������O6��71�:]<��Zۤ�lX͏nbk��  L��ǰ X���y<F�@�B�b���؃0���������ߓ"H�O����Q ��ԭxu���O~�I�����*�i%�4�G+c
�ِP�t����ŀ��:&���jN�4�I~_��a(T�A��Ǡ�l����
}���`���5բa�$� �_S�.�*|j�����L�sb�6�mH8���~�7����;���B�ɭS�|�1�/��S�e��+�e'���W^q����0i��A]Pwi�����qv�1@�b�W^�
M�w\�&U0'#�(P��X{>��"G(P���k�O:�~������z�礵�<��aW�FS'2-�W�,A���\�_�<)Q܇'���ad۹ ��+���RkP�������:���D��ԻQ*N�X���M�<e�,T>������}��T���ۿ��v���S���X>��}`Kx:o��O�2��R����;<����p��zI�IB��͵_�o����$ .������S��	����{'�U���G��Z��wBu�-�- �}R����*�����&��~W�9� ��e�k �����SB�c�lV>q�!&,m�$�k�~��d�.k��|���ŗŚ�f��5kB;	q� �Xn��BSV]:C:T�����$����{]_��KnS����g���\�$�$PsėOCO�
��↍6�h�mw@pk��"�7i��^��W�}� ���"��� $��5��wMo��j_U�ps�I��=��٬���'S�z��O��ϝҮL���,�\� ��s����S> ��I %�g�u;�����b�:>���N����y���� ���>��N�;�yM���e����U�gͳnY� m�����^�ނF>����C���U��w��
�ZGط��ׂ�(�t=�5�i�U�"���06��y��I�Q�(H�V�q�T0�X��Y���y�9�h���|������DdG��*hn�����Ayᥣ��I�?��dDwB��ÞbI�]�nMƇD�U9I��]�G�;��k�0�W��Um����h�U�7��t���^9�'���`�E`M;Wm��6K�(�fÑ�5	�;)����P��ӳ�w3ZAs?��z5��9�6�����\#4(��lk���t�v�8V��xa ��0��e	�lr��	��l��r�����v����x�v�7L`�q�����</ߞۯĥ��7z\���"�x���qN|3����n)�[���p�o�>k�5K| P�:Vh��4(��j����� >�jٌ��S�j�������0>@zV�S�}p�;a&�	���"����ϔ�Xb|�Z�h�6OCI=���rPӔ�_.f�?����C��Q���o���XV�l1/<nŸ�^SA������7':7�>\��	˩�T��rO�Խ`��g�)<�Bt�����ۍ��?��o���%J�������߱�S�3�u?,�ns��Y�ڇ�TZ,�8`t"X6׳x���`�_߀ �Ymq������8X��G뮳n[������{������IM{G�?����"[]
��e�Բ�B�:<q8��hZ�k�j�7�k��=>��j��6����h} b���
2x�s�[�gA��3I�xOSu���>M�H\���
c5�ڏIJ�Q��� �U��B��� �a�E��}� CY��p���{�]О�����@b�꒙b��v�m?z�[�:�6E��;���7���QBǩ���O�0!+�@����1�{hݘ$�'!�u�5_e͸�����ja��@� 	� ��}�sC�[�e�K7��,�kc-�A�OW�hYOI��{G�Z�n(�Y�n�z��q4(��.w�K�d,L�v�`j�,j�|�$1���X����ƪ�g|�9փh��+&Na�W���w0�?��}�1�2ȋy�̕ǥ6)�'|����Kw�Pޜ��:R�,�b0I˓!�c���� �X�_��]0�"X@��MP��ϫ�u�q]�'HXT-�{�/�V���I��U�S���/�:~3�Q����&�	yK��p��<nfC-��8z\����1mnS1�R���mpC\J|K���yC�'����Y������}��clI�j]��I��ڦʐ`�g�>k����%��ŵ|/ݰ��� � ���|���v�s���_,A����Y$�vA4��S%�)��,ޭ�0s.H���6�D��f#��ȫ�-�e���Q��5�|�������',jڠM|��Ϫ��	$xsO4���`�}s��O{���p��ٌ�_��Q���>*�]_M��aɪyb���ф�ׇ�j�3Q��) NU����U������0�b�KFm�����4�ڿ�՜�{�I�
U��c��8�8U�)�ݓ���f}T����
�&�C��ŧ��5$�D�� �D�A� ��S�5���y�E��Ѥ�"���T������ ��s}R��X7`�
v-1�/�S�1�LZg����ϊ�Z��!O;Z�xmn�3
�Gy���?��9�7�Jl˟��`��y�و¨~�E��=����0�'$0�YP[l��4�<^�,44�ܜ�V��k��Gs&ߑ�#D���[0�)���*h�����Y�+��s�6�]L��I���:�O�4��l��醳�������O?�c�9����Q���U��0L��$aπlU0L�r�u״5�����u�ٟZpȾL2?7�7�]+�K���jР�Q�A�t����TAEv
�j��ou��椱��L@������s�j4��e����?��p����fy*^�O)u�p�J�>�!0o��wp}�V-�QBZv�[�z�%$�LϮ1 C� ���gIy�1W:���T��-@&
�)��e胒�X�ks�9y)K��-K��7��Y0�e��s�==�c9��^t��@��� d�����x�N��]���j������4��vK���9�@.�q2,��H!�=��_�e����Jx���w�/�<
���
��N?�X��k_��w(l���}\� v-�\k	��M2�.�6���Z7��G פ����q-��藂��)||n-7��oګ!HЍ�^������%Ml�j�
q��Z(�CҬ�
��Ծ��XL�ݚ��������L!�	Ҋ"�$`��؄�Z�ݮ!"�E_zY2����ظBAd L�,��>W"���v�u�Q�Qܮ�����j��|��}Ҕnu�!r&}��8xz�H|�y c�k� ލOQAR����ˢȅq������w@�0.2�i��Y����,*fn�b#��� Z���,k��Y伣��i��E��f���L00������� ���l�_�Z���H�&�/|�w�i�G���������9H�ޥ�@�8�a�'�B��Į�#t�v�����oI�fj������ ��߲O f��[���o�����m��lG�^��`~�F˻.��uZ6� dH�IV�!��c�7�� U�
�@J��H�3�d0�EqL</����e
\�j8zt�&���^�@Dx .�R�{��F�{��FYS�y@tЭQM��j-�~��HXJq�r�1���o4����f�5��;p�L�6��ҪS`w�)J�[���=,j�.������I��,��"��`�`ZjnF��"�ev,zL���F(x`���5���E�n&��Q�>���&v�(l�z/�	|�Cz����c��.HW��]?�]�� ؆�.&���,f
dM�s�Xr���t��$��	�p�6�rm�fU8U�U˕q�!U�x5x� 4�-�*dհwp��k��$��q��jE�+(�[͔�
��T�l���@�ZTط�hsh�j�C_imڥ�lTz���k�SUuҶqAˊ(�B��wRS�Z�Z�YQ*&��� s�Z����G�����AzP������#�aL<��G�D��&�Q@ �-}��_�@�x.���E��}s:����`b�">/��3�Y��E�|�U0/�,���h�4 Fъ�D{`���<��w��X��\ev|W������ɠZpP6 ���6]�pv��?��H�⷟��g�?���󲁒Ut��0���\&sI�v��\@�.��.w�M��\e�U�x-�en�-�E�R�M'�|�7����0�����m�l��n�8�.Ua<�L����)�5����C�
.�i��:A��M�;�>ۯ�����l�[����r}���� د�������kƚ
���P
&��O?j�	���u<��&>�Y)�5)�����3��|��=��q�a���N=��5v�m�Q��F�{��k�\z٥�8)��}u<(FX�
 ԉ[ ��~?�Q�Ū���b�sYX�;c�hf\��C]�1�\�.�+1U�B0�2G��о,���'%��ԅ���4A�G���r���~3M��Б���+cS��8xןi�V��� #�F^'��1?��Y��R������3���a����馛��IOz҇�A�+��[��z�m��y�{��kO=���~�S���a��Hn��`\�	�.�RMka〾��*|���
A?ff�ci�E8a- }����B8��4CױV�\���B�=��X|���3Z醖�^c&=�g+��炈

Z�� �'�O��'�ZM*�	�����
�a3��6��k��6f|�~��7z��?�����QN�l�H�R�R�r#�3VC�wܰ�Y��%Ω� ��J[�5�Sq��mˣZU(��U@��h�X�A��˟*Ν���-��ඤ�m�6� ��o83��0�d�L���t`hn�id�_X�GY�A�^LהLf2M�2Mp�mt����ԍ(���]��f-�?�8���_6����V0X9��?��r�G|,ϝ���x�o�?��ḇ�K&��q%<.�1��І��Z'�5W5t�SAq%X���Z���5�>�-�2�bF�h��VP�e���x��L��P[
Kv���3���H��g��u��ڦ����~)�O�hY] "�+��iY�d�.`��V\�Y.�ް�{���g����g��Gx�F�}�sG)�>��}��y�F����9��c�a���T�L��ǳ�����~�@qO��G�y�c��Tj{�8�M"��ouƕ���κ��n�W)dN: X�Yk� ����fqm�Bw�k��	]wmS��Hܼ{P�̎�Se����E�mJ�� ��n��@���մ*㪤���a�bl�Me������.,�z��g]��ޗZ���'<&途�^�5�����E��@�;��>M�<͓����Bj.�e�,�*HQ�ׯ?�U(O�{�k��)�5�W��3�KC><�ZI����_�	�18oV�
�A�7�&ு��G�L.��?��mBChJ��1���K^�#����?|�����?��3��ㅦ
�j5�h��o+�"��y� �S�"��6���@�J�[o��4�ѝs�6.�,����c�s���r����;�F��0�M5ձ��,f�3~���0���KrV0�{��}�)�Z|ilr��ǕA�.@�<&��]�����m��k }��!��]�ςi�	of��=�qO��JgD�8)�G���]��K�:Ou�?e�?���-��T�|d���fԘ�!�����&�Ø��$���A���2 8 &�Ht�J��6`��Ų�F��ij��w��_A���vI�չ/�]P��0싼@���=�j���S�pOޤ� 'Ep�6��cz�&�<-1��*�j�2�rD1��x�;ͩA&}pi���a�D$V_el�#(�	OxBsA`m0}��&旾����o�7����֔:F]���ɤ�O�E1S��iɚ9s�l���L��~������1>��b�Z�Ma�@;�;����wj�,LMe>VfĂ�t+��d�4���y����Ԭ��2Q����+���;$Qմ�u���w��B]p�/���i6��NLN�i���xcm�[H�~ے����u�$�����7�a1��7�t+��n1�����EK�t�|�Ѯ&xA��
�
�����ƛ�ȅGkԔ��·@eH�
`��Uk@Zխ�RP-�7��{M��L���k}�mp-�6=Z�=7-x���5�:P�y�=�m|�^���oD@'|-ǮOH�������)~�:�ȣx�
  N����C�FUF d������-�� �dZ��+�5����\��G��dv��}jse&na?n�~2���À�o��h�s�f1h\���4���f'c�:�*PX.fQ�y�	D�[~ʔ�K��B7�q��aL��%�]�!z�<{���6J���RyD~�2���� ��F�����~j�}g@M�Y쯥�k��&��|9�!u����d�<'���N׫��������/_���ކ,�����.c/xz"{x���9{�X����j�
�I� ����A��X�|Z �+$�{uC�l��Z�ܣ>þ{�%RP�u�Y����T��O"��Z��5�i���YpHP��F�JT�làML�}�CGG<�Ѿ��۔%�Ό�����on��|�+G)�ր ��@w�$�3iCH��!A� �d3̙����R�g�h�m�ʂ���������_�*l �+)42	���A6*����M1�+���[M��hOD�4��`6'���=��g���\����C��JM�2}@�/H�r��F����ӟ�t�Tƻ"�����~��%�JP�7s��OC�����p�B�I���'��7�#<.>��v�`�X6WmSm^�UBU���4;M��U���ܸ��� ���l-B����?�6��R�Ts~���*`��f�nk>t�^t���.@W)`,��e@�a�`�B@;�GpaCP�ޖ��oAi�ٽ>��o[�o�þ��j�x�	��<�{｛��G�5K����*p�G�rrk�<�Z �ԢKf�,�Ui�>S�0`���^{�$<jNT)�`b����}����s ��:88Bq+L_,@ѳ�FFӆ�ŉ�#�wc�sK����ܘ|O��Ģ�E۶ˆ�l������.�_u���ҶY<Vs���kD�|f�64s6��g96.�۴L����%�M� u��qi@�i/zыN8���K�ۏØ��-�ez(1�Y�D�:��O�+�1��.�眐;U&�
�I�_�@���)qUC�*���� �f���߻�j�C�2�@A�}s*�����Cם�B�k��ϫ��R�X��e�1�W�6,H@ֱMZ�Zh��ɫ�)�i�|T�Q�!j�|ǜ�9@f����_.h��,?�GEQ���:z��s����]Ղ�y5�ǺzK^��tÎ���������[2�s�L�a2��Y딏��ϋ�ދR�,b��n(��Q�,T7��զ�1M�oY�PfSͨl,�4�U���ج���[�D�LP뢏���U�Z?�-�T�? �#��~s����S䙀M�6�.n��v�O��>q'k�O����X��B'?�i��9:�[�����	�_Ja�'�=0��.�Q��j�֪�Y���\��x-o\�&j��ĭ��k���`��j��e���y���g����Z �WK��E�Цu�}pX��a��mK�*��g�)�XCS��-\�s�U�N��7�|�;�ҽc��[�-��,sn��9�y�(���@i��=x��O�5�\�Y<cim��g�}v���=�!gP9ߕG7�$�c7�#��EQD~8�6qsi6A_�K3���lЗg���)�Q�X���AA�
g���ؠF�Y���15Y�Q��F�b���U�$V
ж~Ǫy�W|�0
���`�h&��(荡Zf־�P+�ȬymY�$�_%��8�6>餓�FtD�N����13~3��Դ9�_s����w2�''᠔�~z��������g 2�ꧯZ��dM*���B+��i�4p=�=�Uk�gj �.����Wf��`W_���u���?�p��U8WA?�$��+��Ep�5��J�+�Ƴ]Hs�B;�s-dh��;c��X�{/|���-e7���\�����E��"�9�V�>�1[\�z�w���_�*Ҕy �4���[�e�9�a@�; ���]ʮ���A�O;��cc<"B�,d�!<�,P6��M�	�j�\��1�`e|��� T�����F*�2U]��F,�����04�Z�\Q7��D��m�����V
�6	s���o~�����9�N�1�_OV�7S���lIܮ��B����5m����Y�-�PM�uXM��Q��֋�+�C����k�O�=��&~�{���ep����"د���ѹ�۴���o_��$����4�U`	
Ԧ��Gj�Br
i�XR�����j�����N�F@�t��J�}݂f�����Xhx��R��F�'��������5RGQ2)�	X�HN[3ѿ�%-J�|���(ps������Eߑ,����;N;�'�cv�/g]@�U�`� g6��E+�ԷV}z\ѿǆ��F�,
x��9�a�{��s���6�U@��Lk �b,h|ƍ��0��I�2�]fEh�`�'p (�N�D�.V���Vh�V��l����9#�ҿx�!�|1�I'T��_s��Gl��I@�?�O<5�k���~'|��%�n�g�	r+phUػ�+�u�&>�]r���.@0�l���־[[�F�Y�j��z0�+�k�Z?�rB�P(����wݗ�L>�۠~?�} -xA[�o_5�[<�}��68�wx��R�p��I�^o�)��q�|sGPݐk�{�I�g�6x
A� ���}�T���!�V�+_���ǥ?s��z��IK�5)^��0�#r��a���'�����&�;oy熔S	n�G0�GT+Cc�#<��`E��4�	G�n���M`�!E�uʹ�$�V	6�Fبlh4y̭�~̀�̖0(�BHb��Q{3xh`8�tto����F���r@�n1Eo���|�ɇ�NNk<&A�ߊ	��K�RYf�����թ[p,� i�
���2�P���rP�jj�C-wh	P�*8k��+]u?�v�##,��?�������J�ý#�m���p����`F���X	iQ��P��7�ங
�qA���u��g�����
�!8�!�fD���S�������f���e�#�4�j����m�z%Ma����7y����Z�<k�pF�H��㪖�!����զNfd<�=������_�k���6#�Q8<#���j?I��EK: Bu�w�q������Z O�kjlu�����PL)�a0���� 6���</�6Q���Ы6�F��6+υA��gί���?��7��(T�)��~� ��`c��I�~�LODK�sTš�&��]?|�k_��D0*���F�؛��H�����}���=%������@W׀�5�I� k�t��v���Yk�j��'� �&�&��k�;mѾC�)pu!��U�4��_�Պ��Z���$�7���s�xM�j���g*D��c�S��]����;��i�38� � ��}�ŏ���r2�X�Z�`�M�� .��q���}��gt�_����i��O�)�S�U���lT���|�U�ߐ���V.�E~{���s��0�kһ��u���F�><�k�$��d�V���JS˄z�o�q�@���(c|���@����I��w�/�Rj���
i�GC`A�f��@�lh4y@ ��nHM���?��V��A�C�U7���0�X(�Kq�$Ui�D'?��x�'���'~|���a��3"���#�����h��&#���n���
ơ S��ÂW��pH�� ��"�=���[^�E6������(�̻��
�� u�~�5�
�|iI��F��l���]$q����{w�G�5�����ozӛF�~��H���8D��{���:� X8&Y �7��ߡ�&p
_�����5>� �x��L�w~f���X5�Nlÿ�8�����: �����8L#��p����|�Օ`8�x�&�&�W�V�(h�>86�7l͢c�Ap�A=7��=f&�H4SVA,c�W�w�h&���F0�ZB���@� ���P`yY-��x�1|����n|4����v��S����/~�?3�Ǣٜ�l��ec4Y�x_�ЗR��I�yTή������hY�
�*,��W��L�R ��xcX�7�U�,���]ۦ�c04QW��)��e���Z�j[r��C�5R��3�R���?=�=��}b�&~g���=�� ���~g��?(%��Og���@`1�G��R����?�CsG�\��<Ү\kj���Zj\'� އb�g\pt�ޚ��SfC�%qMK��s��a&�p��h��b:�_��qܝ�d�>����ŀ�^}�l���D�
QM���-z�"|���$
T+c�s�$�}���M�qI����� �>����0k�_m�ͬ<�jW�C��Z�ޔvW�6�c\3�$��ѯzի>~�a�}2L�g&́�?�B4Fb?�#k�S1'?%ŪԎh�
n�E�Ռ� ��^5�If|H��kn�-}��� �^L��f��>��1����a��P�U���A� �
k�u�1�g��2��공��+�- ��g_����K� q� ��J�o�t� Sb��E� @��q�5w��;���(�s��B�k(�k�f|�5]��I���\�2�ǧ��=���D~����A�8�����l�W|�����1G�T�O����&Bx����:l.��AM
a��]͛6h���lL^��FD�����px�����  	h �;���H@��m�j��Z8���*x�{����h�0�ø���J/�i�����Ƀ>��1w�lq�q��(pȼ�,�_<�c��t�3�w���C����)}vO��jVt���\�g��)X�xg#0r�~K!W�Q���Y�|3C�� H�np��o�K���4��U���T��ʾ'�� ���&K����Nkӭ�m��t�8�v?�Ӣ��8N�h#4����@K!	IȾ'�T��R�}����y߿�M��]@TBj��p�u�����9�{Ϸ����l�Ƴ2J�9N���ڗ��e�W~D8n�N<8����>�n�����N\Ih"�\%�.��{悠��$,p��/})j"}(��D���@�/t�d�yM�ϤZ�ͷ�z�Q3�'xf5�k9�;!8��k�i��������w>��2Sy���Prbd�'i���Q�i�"S '��+WY�8�9�q`f�pD�*L���	UdE*LM�Ze����s�S#e*���b�i������n�ʇ��.��&l�sBT��4-���c5���_��\�@���埱���i`]�����e��Q��97#�� ��ٿ�:�}���ʙ�f
��կx^��}��}��b
J��hG'�]��W+e����J8�4�2}'D���i��"�:gh�1	U���q
��K$�,{,�d��LmIv,�
�
��%@"���䟤\�A����QH���Uq"*a�������k��{"-("S�sEN�}U\�&�O�V����"j?L��Gfć@F�A�`0=�S�V�ت0�|���{0�́�!5��5i���>�6�I�����Aȁ����h�� �JG6|�
M0����XI#�}y-M.�6���iF�����O�*�D��H��{�񊚐W�LzR�j���Q��C��Nv�v�΁	�� h�Y�b�����7�FgO�xv|&?a���[Q#�# ���/*�<�ץ�
m� ��vB�ʾ#�"�)b
`��y>i�:�U1�"�I��o"aā�U(���З'�R�k�cQcG�4����f}i���KP�T���/3?R#���h5�1OS��Q������(�~˖-3bI� ����@�
9?���=��y4��7��B�N�?�y�{pl�2����O'hMAO�?ڻg�_����6��w&m�����I�ZB��EjwNJ
�*R���Y�@H
dG���\iez/k��T�K]���z*QJ��I��ڪB���U��PԄ�|(��z��Rt?KK�}tR�r�C�Iźu�n�*�$7��.ޏɚ�����<�|�Cۧ@������x�E$�̷!g��^&�"��kh��٫������+�	/�9�W��$��
�͞k���־���1� �>��?��r6D�D�Rn�_����=9�Xg�$ "�O� W�$��wb����|,��9�X�t�p̦�)��h��wUN�<.:�-�D���3��~���<��u����A���Hq���`�=�r�F��_bм2��a} p���Ȝe��pTR#<0�I�U���#b��/R�s(&X�k j�й4�i�"�V��I�
� f�<'I_r`�'X���$���K�sJ�(� ߵ��jFD$4�/'n�3@��#�����G�����|���p:��]x}c�L
)�9�9ʦ.�j�x[�"���{�#�4r�^};\����!���K��g�z<��}�v#$��>x^�x-��9�3	|H��ʄ��� ���~720��40J�F�9>�����oD�������FE��7� �����>��h#�b�c>�ҒR[�������=(��rnꛟ:������q,�z����A��Nu�1h��9��.x��1��܄N�R9�i���W=ZQh"��;R�j�^Aa��K�W�29H��&#9LI K�(�+GG�8pU��q��A@bC�,Ձ\	([��f@Z�pŤ��d���m���((y�fac�NrX՝���}�X�\�����4�2���6X����O���Ƙ��+��r��Lh}���I���D�g�q��ߙ�S.�+3C�q:Fd��Ri�9��;�/����ʕO>o���a���"�'�5vB��'�$�-�I�U?��#���p��v	�'W��B(s�L-���~|��If������Q�"���;ڏ�@��s�q�����M%��L?�9~�q\}2�=�qB0��in#+�A�~6�נ���^��'ܛMo�:�`�*@	>"�hO�D�$NV��(MAh�ЪF�U�����P6O� ����8p���2ۤ���E�L�n�XB?+M*�!�~�{V6M�|� �˩P5�p6<�L���/���p�s��_��G��-�8�-E���,_�>;����S��ꇡ��wU!�o&p5��Rq1���1��!	6��^�m	��[�G��?3��s�����L"¹����q<��h~��5�=�\����7�4�ﵣH�<M�99 �Y��'  J�IDAT(�
��G���0���*��\(h�8�1*S'�-p|�BC3�� �@t���s���`�=���^>:Y=����0<t?A^��3�怣�� Ԥ(3�����q¢M���\+�G�?��߀&]�W��B���BY�I:q����Ī�C<V�T��){px<��{ �a����Uu��8q2�3&����<����7����4=r��� �~Jb�&��A�o1� �z,D?��
�a���ӽqV��;���Q2�q؏�7�!sn�t@o{Fذ�Ӈ���}T���R�k��#��j�NFK�s�p|��6�  ��� ��G���Ì�3�i">�O�:xȖ\�$">4��-�G��`{Ix��z��G���EU�2���oĶ�$�y���wN��S��Ԑ�C0$멽)��z���ܗq����〢 倖�ov�{r`j��;H���Y����s@r��N�X�!h2����JէIR�'�K5�j�U~
s�d$��	��&�N�uP�5ǉM���2?�T41��!SG8��M<#"�Y�0���^j�����@ $�+�;�f���
�&���o�H
�P���E����A�fe��㪛}�2��(T�69�d�i�%�y9.� �~2f�f � �:ȴ�L&��kS&O��#gJ��'��gq#f�C�ڣ�I������@ā��y1~�AV 4����a����`��5��靦�cp��$�s�<�Z��}����
��b�Ze�\�s
P��9a��+��,g$M|��7�hB!��y>9QpK*��!�5Q�y�|ʙ�6��ܟ�HN(Z���
9.R�ɗ'V��|$$$X�-��l����������Z������
�n����s0Vr�"gߐ�������\J�9�M�����ƅ��웪+B<�E�k:�r5�ߤ���� ǕT�!i	���l��p��IIǣ���/�DŃ�W���y�Q[�J�|
��u�
8��c_��LgAEhAjUB�!ϣs�{�Ib�j� ��� �|����o�1�7'C���7�A��LD��9"�ք%r � ��y����P��I��r�^�|��ݩH�)�o^Wj|�3\i�����tp����<��i4��z
�'Ai1$�y<?W;y"ᑽ����sߪ$���]���8!x���<#T�LF��_�$���0����~%��Q���:Y�Pm�{���W�[��\����E���_$�h�)6<O���4���@��ۧ���l�(_���/-#�9�>�9�Hp�ZẆ�Q�B�x���lkʿB��6�(�@s���	���+���I��S�Wڹ��'2ڃ����-p��D��DDZIh��A:�e��	GU�ys��F��I+�=m��*E��x]9(r��$�I����ኅB�!M\-h������ϧ�VLrbRGid#e�(�y^z�Z�&c��6�OEx DrAf�.�M��x�����/��յ�^��3��3�a��]�T�� $!��X�u� Ia�N�PE�ʥ"��:�T��|�	a�V�3�u��1*A�N$�|qUwTr"FQ{��i^`���ѕ6}���7����#Fm��S9��=!\�M7-Gn��%����W�n'o����/p����q�D��Q��%[9��KBQ���5J��l�k /Q�by_ˑ0l$����2ղ�\�w�ȹmڴ�D�d��9��Єb�h� R@a�?s5��2�j��q�ҊHUT㪮�B�q�1�6�(>L�G }��m5�p��Y��+�ރg>N6q	.	�7{ϼ��S��Z��/G$X�[B�����Tѓ+T��54�$�lsh��&!������s����;�M� �sLp1�W�W��!S�3�A"���o��Hc��K/�0C�G�4'��$+�D�,q ����;@��]�'2l���a�������0X��`��+	v�2���ohվ����͟W�D����l����d����j_&9q�����T:`i�����m��֟�����&|�C���0W><	� ���p���W��\%�mPG��z��=��ݓx�/"z�z�0�s۶m��GGe&�:Y4��w	�Lr��ҖIS�����~HL�=x�(�a�}T��
UT�D����	���s̪���Ӹ��Z8�X	i~'AEy�����Ҿ���GE�X�!�a �!)���{�{c�u"z"��"2�rΈ�D��"��\�@�{sB0����}��<�+��VW��9�x����Vx����4�ej8H� _�i{grj
8���$�4�e^��ˑ��)).AܡE�̩v����"��j��'6':�P���1��)B>"!
e�$�'^NP23��$4%��U�}h3qB�{�ցs �K�>s�o@
>��s<��A_ɧ�HB6���:�޲�?�i�H2ٟ�
����!i�92�Z�R�X�89�RȲ�����γ$o"���	M l#���q�>��p|�h<H���Ixs,�����aXBS?��Qr�������Du�)��/|!/�x��}�� nċ�:��@#�/K�,�M����ޖ8!8��꫃����[WL��F���ޕ���a��l}�߇�H�����(l�Ҕj�߫,l�mЄ�H�ZRT�<��D� �9Q����x=�i����՝�N�M)�C͉��+*A���D����	5$;8���uG���'@jI��)䝸������p.�Q6�ǒȀ�[��oL����ϖ�P^X��qy�k��|$�4���|S�p|p���r|��v����p\�/���cD9 d��M�T���96d"�8��?�sC�U���[x��� �������v�hh$��H�y�Z5�Aa�";}QJ������+@z�y���8!��{#�D:�1�0��V�����#֏շV8�`'��h�`R#�0��$�α�cV\R��/W&�V%��	Q�l��B�b�M�r��7@��s��2�ីz� ׄ�I���%��Ä(<N�@d�Imʕ�� ܗ���=���q>���{�ҁ} �Xbo4T?g*d�\g�� �19ױ/�߲oj|ɾ/���r�!Q�F,LN��$$���$/l��c������i����1)횾Ǆ܏}�������c�������������{�g��XQR1e$�����I`�7���k������0x2}�	�ɠ��� 
����wB~.�3��H�j5��ܜB۾��VΑ�����*c� �*�o�$��g�2&IP��|d��9Û�VW���Ɍ*R�69���e���$��
!���ĔM�c������S*UN��Y���	�;���^{����Q�_��1	�Eb��a��ð�_aw�V�7�C�r�O
�"����B�s�̠�A�^�+w�꩕c[��OLS�I��2�5����
��B����@�9����;����6q�R�S��\#���T����F)�Ip+�>��B���`��6���8!x�!>'�DP���?�3�YPݗc����s� $��8YP��[�͔)#/}�;�?�WY��'��Xi4Q�����d�� ��C�l��ٯ�}h��ID���O��Ɍ�U�M��D|Dr4I�f��>˜ 	������o~�~�[��4��O�7�6}�QO [��x��j��$8��X��ҋ/]��7�l_�U��Qee���"�������~&�Cg	���5�8�To�c��,��(�4d2���'� �W><������<w2�;�(�yn�1gFp^�&B�:���y��:��V�� H�vw<�ੋO'��M��+�j服7."1 ����tL&������";����Ç��L�Y�i�A�)5��V�<���a~Z�]�SZ���P��D�AP���s_n�W���4	��d���
L&��4Q��A�U������*�O��@��U�������ܫ;E���n��]��������/A��
�S���S��q͌�W���" #�>Ԣ�HS�+lV�~�����3����Pd@�V�Cr~ǿQ�>��O�]�˶�����w_�E㪟��a�e�]�Ñ�K�>�0��ϟ?~c�	�N��$P�[�@uׁ_X�g5j.�})��F�1i&�8"}�}R���䢤C�凫��l�R�+��˩��~j
�r�D%�+�7ߕ��+�H�I��#P����Ofh�VW��V><F$B��������͐m�6T��@^rak�v��R_Bv?J���}th!��݈;�V�/�n�M(�s���R��K�������ȯ�4�W�_�0W�H��c8��W�
�M:��G�� $�zZ"/��xBd�`:�yO���xi�"��~H��_�T!�1R?��2�zûs7�!xwp�WAȃ��C{��+L�d ��$$Ed����V5��_��;�ġp=N\Mg�Y9�i2��犃�P
{y,��U�<�'�݃���E�Hu}�QyكE�����<���a��H�<r��785"H�������H���\�eg7!9�vW���?� ��g�����OQ�J3F���$U}-�M��J�\���V�����#gCi&D6�o�8Bm�ƅ�;:a���d��|
~���jh��9��U���Z=�+��u�]\��+��^�N� ��зG NRK���/�8ߝ-�i��5��4�����&3���֕%`C�*I�
��L!(UB���`T�-�
յ�r��ה�U6O�H����O��p��k�ebԄ'�H�L�ꎿq��*
��t����_��൷2��`E���+V܁p�[�J?+�e�$�&)�K�@����0_���R��R+�7�t�q�?B�+B�C��H��=M#�'x�e�%��4��= ¯!���W_u����&��s ��	�@zC�-�����7>���<�+ �N�B1�y�����pM
t.�&��j��2�Q��:
��ꟓ�2��'3��8�1���A%by~�/����J�r�ʌ,��M�ѻ*��w�둔�N+jF������AR@5+���������]wݯ�`w�[
@�sYj� <�P�Db�>ʾf��a�� $�;t.Ծ�Hi�/JP��q8ތ���D�E.�E��PfA9Ck�!�?E���Q���C�	�;����M�*��F��gϞ� pc�R#J�"�C $Z��a|�.H`�A�U����s��$ItR��FU<��FE��
��R>�$�>����Ve~��T������G��|��DD�0�@�5K��K�#��I|ݺu��-?���+l�k�S}����G��U�V]�><}3ƾ�Wh��@�V����O}U�i}f_T�?����f�Y�?j#������ٗ�InHty~�z�9�D��'�X�!F�`|%���}w�Н
�]���հriA���~�����w!=�?79
q2�
Z�T�!ho�ʑ��2�,�窛��/eT��R�|�s�l��Lu\�9Nmf�(��oΥz�����a����9�*�&�pr��}��!�
q�=r�����`�x&2�}�sB0FJ �
ҽ!�K����W^����o�ܲ��W\Z��Ƙ�#|��ʌ�O��x�u��21�|�DL�����="��������¢��a�XO�-����></
g�;F�w����:'�00���^!O�N���A��L�i��d�U:�Q0����r�	#��`�1c�,����.�ɖ����䨘k9F�Lr�R�^S���8sb�$<2�{iOH&xO!�����X�x��}-�.Ap��0n�ūW�� h	��d�/�ewI��	��V��s��ߑ|2g����{+�5v�<+"���}~F��{�w�y�C�\rɯѷ=r��e��b����� �~�bsl��D�eMc��
/	�PE�	�������r�K�+q�T�ޙ��Q��Ģ��\�qJ��7iD4�Ʉ�|�|�|���U���H����Rؘ�4'�<$$���A�FGp"eV9�W�{�ʕ+��9��A� ��}�y�K����-[�,��FKN���G�$����!�1:���e�����!a#t8�i�C�nC���Hz����|	���#<�����?�.���m��G��kY����[�2�	���[�@�X	��W!����!�Y\ag���yMew5r�
W�9�,.���V��Iq&����L��J�Y��V���ٳϴ���~�ܹ(sn��K/�l��>��/�R@�qO*��lO�2����f���Q8�vh�¸;c�T>,�q��*Hc��I���Pc#$���0���ԫ�������{�?���#H;���{�v��tް�Ӊ�0�6<��������0	,��!W���r���\i�s�a���][(��PE9#�X��*ELR�j��/3\K�6▊��B�� S�VJR�r��պ|�xE�	���}ץʔΐ��i�kҔ�6
��3g϶�3fFm��JXWG����\;���J
�(/>-��Q��]�:�oa�$߇闈H������\�����F>"��aLhr�y�S�g��БQ������@;�3��m�����Ӧ��Tç��:!8=���	jݏ��o}��_�"��LM�m�d
�P`rB��Q&��*^Qa8��8Q�$#��@KD0 �uM�QE��������8�%����P��^d�`[�R�d���l�z�T�+U+	m����#�pJzw�:c�MC�������Τ�s��� ���r���=c��-W&�:���֝n��<�U�o"4��g�y斧�~�V�跅*$��pY�[�ܐ)�߇$��#�Q����X��8L]@V|�x�s�Y�D��vT'��a{��o��'C�G�?���h��C;e&0Z��{����	o8FW��Ī��)�?��x.N\���k+7�����CǪ(>��B���>�䔑�פ6��$�PH!�W�8�Bm #H��g�$�0S���%�QZVwS9Ɗ
z�*D[w
�D*L�ҔO���x��O?���^����ee#�J�q�7��=x����H�x��P<i.�q�� ��LpR�*i��1!��ƤƘ�4�85e'#$��{?|��Ň�c����)�};�x��i~ ����#?���}k�Ν�Μ93_� a�@� Zy�7i
ҩ�&����I�X5����u�� М�T>��R�*TP�ahй�>	J3˙Q�\���G�un��+�o��~M��>+�Q�sr�Js SĎ�Y�@FY9�ě���u��cȋ�_`=�^tt%���>�ۋ��W]v���/�7��A�q��z8��Nd=��=ga<�4>8F��R�+�V�?a��g��V򯺺:^��A���<~K��88!8�bX��g��?��F�����D	Ae4$0�΂��$hE����uvtFd��8ё P����dfC	�t%�VC� ��������ս|DXB��#p2e|5?�-"$|�̶�D���� !  64o���Y7C'��D�O�>�Q�XXVn]�Il�!\y�7_�hᏮ�p��-.*�X�a9���i8����/~q��>{=�t碯�Ps�>F�O��r\�|F�;��ۃ���s��Y����/���^�{ �?'��&1����o@�_��R�+e���H�V ����M��T�W�O�}_L~T8��%@��HO����9%��d��
��V���秐B��l��4@UjW^y�>|�~��_F���S��Q3 ���J�#�T��˧��H�K��@΄,�KHA�����ZW<�	�tܺ��x��!�N��t��ߜ3�����~�T�<�g?�هPD�ZDǜ�>�C��~,_�Z�Wi�N��K�%���F'B��Dx�5�<�l�^s` wB'����Amy#��}�\�Υr���s���購����Gaϐ?&&"��J��oNd�W?<���)M�\�SN��l�>�I6���geD�@W� e!$Y�'57^��v\��	~T�4dq4��0YFZ���RdV�$ɬ$�GHC��4���K�e[.�@��-V ґk�+��"��im�]֒�L��<�_j��vkn:"S���g?���˿SR6�+$��v��>� D��׾�w>�J�Wk$4�����ζ��>9k֬��{���@�G�|N�ʾ��D�	��D߯}����?��_���L%C��^Y�S����?eJ� mlj4�7Se���AO�a1i8�)�P�$"$2���Q��R�ܔ��D`ܸq���p�Er�w�<�w�x�P(f6r�"?�&@C���mI��p\:?7Z�%;�f�my��N&,��j��x�w�ؙ�l����t�$���v[m�aK���`dŪ�]�Յ������D �u!�!I���������}"�'ǐ6�5��$��&�~"���������g5�[JR�O��O�����X�O�[*w��)� 3�5գ=Z�{�p�⊅��{��@A�� "
MT8�r�S�З0��N���4Pk��p��k�@)�)��ƘD�Z �i옱�_л�R������I@��
rX &GB�p�lkg���]�-�(�pz�y�A�)�B���C�y�;�t�����u@
j,��ά��+'��޹�����1cz��o�@� ��.@DЇ�cp-|`� Y͡Ƌ}���>��Ϋ���Q8>����C�	��{fC���_���>�$*��`���T]PE��#�@!� e �u�����@�x�=vH�(yUGD�����7D�T�r�zTy���e� `x`Aa�����y�V��A�k-8&�"��y��KK1s�e{I
)!Hd � �`6Ē��ȱ����*G����l���=��ں�W6ۊU�۶m;�3w�l�v��"Dq��uv��Qkjm�݇�6�?����=��y/����֘���C �={۶m�/_~���)a�<RgW]t�E/�x�+.�첧0f�
� �5N����j����D̓O`2��ln�:)�sa������䠩�)r��ʝ�� )�)�i�W��V����_�]IH���F*�|�%�U�	�G���THR"G�x<���IJ{�(q{{p���(2o��4ÿ�0
1�4y��a:VU��)"���>Kf7J��>js�c��e�P��?z̞�pО��ZO0b�DU�g��:;���n�b�����;l��}��εںc�wp�\~�E?8aܸC�����������#5�b��4���E��G����m�"��`�>���p�1����x���?�a�@ʔ%��^9��ҡ2�@� ��"(\i2�F�B�+n
h~GR��C$�c!C�F��� �I*TP���U�4�ݟ& ����s����+��D�,/?/�;�M��D�ۑ�%�H��7��I�pLt'�0����hw��$����	�@^��(:��� jH}b���m��`oԵ[C�D�qs�����$1�>����;ltO��92m��Nˇ�����η��;Pu����]�d�7�͛�4�W%�#�i<S�~���� `�"G�� �����¶��}
r
������ΩP�`
ii ���$Qr��T�*�D� ��ߨP�A~��guA��|$�&�P%@s�Q�C�
m��!H&��ϑ9�7���Aɋ���n�J�_�fE5�}a��A��}�&��x��N�l-M�Vw�&�I��D��B+Un�5��a�;ڕoSf�g��α�t���2�#�,667�� �a�P��ڹ�&��ؔ1��ƈ�]�9��g4�4_��/�@F��C5��5�j��N�rG�p�I��;�. ���w�}_B�����_&.R*�0���Ps@AR�
��������R�@"@�<�I�p�6}�H>�/?�(�dH���ꫯ����L��N��Ĳ�q���^��ȉ���r�����nh80�Xo�	��	M´�q��I'G�8{���ڡ#�8B��qla���-]h��eV՞e��R;�B�Bv�TJD��ѱV��B�o.B�hUx_�H�L���E��b�I�^���w.\�(x��(�����uN1�!8� ���0@����}�+_�!�&|I��R�*,1�BPJa�赯Z"�w9*�QD2`~He���{�aB$�������=I�ҥKm����裏V�'��0��$T����{6(&NEۛ_����6�q74�]��ݱjo���|��y�`���j�N�<�*'��y!���Й@��9��r��(���&���-X�wk��eȄX��)�J wA�ڛ�B���"�F��撶L	 .g̚��N灐M�6d!�'�F��-�S��G` "����T�M�	��˿�oܻ~��@���� �bH���W�"T�3)�|�C@M7e9T��0�!ϝ@�]}]�о$t�P�;Q����.C��H�@m��/��!z�
F���eRajh@A8h�&���� �"�P/���)�l�����ȶ|�b�w�D�!�#�#AON���(��Sf�,������?| D&m�3���ܹ��OANr�G��,��k�Z-�����E��1�1H@
��9����L�)wFf�&���a��,X���0�xE���B�	�z�C�V��������������IE磊a�!���:���1���� �;	:�I�@�ǿ�@S�j&�B�r���_�x�}�4�\E�����O��IP�[.�-\!\c�� �v؈��v�+.C�&���g�h�%h��a5��SI�d�k>Vo[w�}�@T�2W�HF4���l$�Z��H]u9Z����Dd��4�/u ��X<eyp�Jt��=0��� ��A8�وCA3Fr2�#��f���Z���Q�G=�x�{�3kƌ�C����9�'��I����~�C=��U�V}�|&	�87e$��@1�t2���g�#��iRP
b�2�qt`k�<�F��H��`����;�R$�{�+VD
眳�F�WXIQ1��vKuwA���q�fXy�xˆ�Ck�6�j�7�5��jc���_i�]8����}����Ax�`�`�^2Sm���� �cv��֎��Y�E=�=�β:��$<sP�.���OA���4Z@�Gj\#� �3vu�G�����C�(�������������z��JKKZ�H��p�-�C0l��q���a��6V��~�ӟ}���k�B%�����k!D�aw/F� ���P���J���F����ȉ�A���=�X�s@�PBlv�d���GɆHFh�(�(�r���`���VP<�벗~���l�����U0�μ�Z+�j�'^�e�;��&ڸ�����5�H����2�D���Vr1�(bT�u����Y1��~g2m��v�'BjE��o�[T>��C����C��ބO C0�4Cь����ѣ����/�&�H��yf��9��Վ�	\C��aP"�}�s�=w�O~��#'��D����'!�ڟ+}�d�~p���skKo�A��y���H��(41*ܗ�HI�Y@����oH�jӦM���v�ZC��ȷ�D����r�-H��#Y��(�"��Xw�(�qH#/@�H8f?h��{�(��F�mta��,���h� ��Q:ҦL�em���sѣ�0�� �$-���GH$�A
B��Џ�C�7�K�cAT�977�K�@Ѭ��� #F��xT�� ��q�Wl]����ݻ�ኛeg�F;�@��k�#J h�|]����~�S�Up-�u�����/��� jH- �Fe�Y��sh
(X�/��S�7I��x	���2�E������$Pk����{��"i;V����2+5��%S�	�
�ae�w�p����$!vܺ��8V��K�� I��ǭ=� M~AO�5�b�$&Y����E���<+�N�|p�� Z�GY��/*�Doì��A�?L@���II���8g�\�5:�>�F��ںڼu��?r�������3S&N:6(;�7�p�x� �ol����`;�~Ϧ#�=1�	���o���_@aNM5\	˗���T�M���0�J2G�LGLB��H�;vD�M���m�F�[o��(w�f�jh!�Xń�6���,;����,+d
��p<,�n��H8������-�w�!0������e0]oǎ�ŋ��!��?bu�k�� �*F���x!�	;���B�I�r,��	�L��[��_BGk�&0C�Q��sϞcS���j�w���.[w�ݎ��c9��t��xNq���M�zG`x#��������#��a��>�3��|� �`�^�\��H��J	�(p��dE$ E��
� ��cH#(��ꊊB����^e�e2�F�/
~jh�Pb#��H�2�L���˯خݻ,�рRȕ6��yyeX�3
Y�+��#/:v": Z������S���'l����(H��+�o��m�{�Hñ0�Z
�FH�&Csko�a
���hE��Dj��c+'ڬ�����B+f�##bڪ�l��F۵����ف�	(�4�FfU[yQ{wv~��!��71\pB0\���od���v�����ރ�+��>�利� �ʟ��ؽ{w��G�H��.2A^Q�">+�Q}B�xn�HH�-���7�		�i!��x$�!�N���\eSwL�V���۷ظ	S!��8�j�@d ��B���׉�=U�i|e?����� o��� M�VSs[��(��b*V�|���,�����l�ڿ�5�Y� � �9FMkSfͰ�2�>@]n�ȏ���z۰�����@�H\o�%�ĨQ	y��Y�*�TI��'���9���E�	��}t����5k�.�{_z�gQ��8.F��1��$�)�f����j�`�C8������PY��V@�@Z^�	��[�>$$��ۑ��6c�L��aP�������U�l����-@Y�(T34�R�s1��G<�����4�$,�D?�=� ���v����M��؁��L�� :�� IQ����*�bVY09���gX��U%�� 箮k��:l��.;p�6�R =Yq�e�������	�hD�����*��8�'���y�������͛�>��S�"���H�{�#n��a��ٳw���P�㧃���q�=�8,�,?
|n����� � "$�
yԹT�(��8���jd�2u�U�T������fN�i�>��ܻ�{��;��L�R$_B�A���� ���f���©0�H�4�B��\�f ���o�:�)4#=qww��5i�֚�5}
%-@�(�gP�ʋi�S������MV�Yh�9#�;f��:�e�D8Ƭ䥽��mZm�s+��l+:��8�'���y�����k;R	����
Qrca˯A��Z��޽u���W�\�Y$z?T��J�,M ro���XU�/"�����X��d@���F�^�]`�?T�t��G��ț���7m�h'L��S��4q�͛{�͚9�klú�v���R��܇4�0�9�ڀ.��؅s6w�㻘��� �!A2R#�s�	���aH6�!;a4c�l�S&��1�A�Y3��� ��@��n�����[i�8�*B�dF��P@��,�0
t5�Y�*�ݺ���h��_�y�G�-�%s�}s�������ԼͿ_|1��e�]h^G�����/�p7B0�J#�������!�����ޜ>�E�����~��YB0���T��aB��6$)�8a"^җoK�-�g�4[��*d<`壒(K��"�� 'Vd�.���|�k �m��ݰwuXckc$�s�n_t�96vJ3CaLQ�������Voo���u@:6�Re -#iz��"�(��%`b �i����j�:;�k�u�n����?l���Ҧ�\�P��p-N��������k�����g���իW_�
��������$�4@���3ܐa����؉z�h#%�cџ��3?��5ccHA;<�۰�� g�P�O�	�>`k~��~��Uk�8���M �B���򡶏��,�tI�:!�;�X��)b##*F#R�l�g�� �P[Cc��q��6�i�==V�S�R��+�@̓�j  ���{Wc�j���T�#;^��]k��v�i�q@,Ղ�ᛀ������9������wo�� @���['�mH;|L���p&�ǵw�#�_n-�<%$�<�Ah6��k���w� : F$����F!8� �Y�����544!$d ڂ8�&]t��8u��ꩧl
M�4I�pL�*���apd0�i��/��S�Z��@6x��RVէl˞۴����0RV�%��]��T��@D@`~Ȯ7km�ښ��g���Y��v�u7��zdODHd2LŘ��6�Bҽ�|s�A���A�����p���lٲ��^�t�kk��:4��@���� ����P�̇yJJ�R������@��H3 2��H	y�-���<�&[m���ֆ��S�M�(��������m޼���k�έ�2�AވZg "sTB��_P]�:���v;��e�w��n��!w@O��a�kG�B!"��L�f���ցj�-�����뭮z��6�jYSMV�Յ��Q��̐UَC3A�FdI@�An��7G��8!����n 0w��=��8%�B�B��/����i��L?p�����p������ύ��ׄ@2@�fUAV���1ȇ?+:�o�5����i�l�h�>�ib��e6y�����ȡC�`�<{�³�r�8�`yO"�H���	�'�W��Yu�Ⱥ�P,���H$�	���BȌ�s@^��:��[��=V�s���[K݀�hg����@3B6ڟ̱ڝH��:t�Z�� ��SwV�5�F��k8�'�\?��A !�͸���@�X�n�)�>s�[����G$�U�dN�|#� ����C�!�ޔD��a������YaA��?�n����ցBC#������&�Hm�m��joT%�)k�I��������hCv�؅���@t�챖��XgG�l����Un@dD����$�� ��P&�!��Sր�X�(�م�21�s���;����;q�'^�px>w��S� ��Q���;w�)ÄPA����	���'�!�Q����1��CZ�dV�� +��?q�H�D��l)�֐HE��km��zd(̳v86�K-�ͬA���]h�Zl1�H�Ls��]V�c�5Wm���=�Zw Ս�,���S�ɉ��87%H��q�o@� B7��s�&-\����{�c����>��p+N��vX�8&������Q�`B��Qd	��(�7��&���'�Ȥ�@�Q�0�:�TI�:�ɟ�I��0f�L�$��l�:X�`6H[��Pa��JZ���Z����l��u�~h7r	��!��M�Fzd�2�:!*J"�� ������@	e�4�Lg�C�|~��KW^v��+'M���>o�#��4NN*����@$��e��HZ4%�B`�F!k�!��p4@#f���L� �4r��ܒR�7���<���֔;�:�1h�E�a)���ƩK@z��[��>�"y��׬�n�u4��·O@64,?��5$ N���Bh r�	�X帥�a�)D ��,<眍7��G�-�tٳ3g��YPP��
�9��PA�}�ʓ��p 3�$8�R"�����u.�_A�*)��E)F����"�4
0!л �^��]��!Mq�%�؅j�ݹ(2C����.K;fG�D΀W�~�fk9���B�_o全�XG6Ch#HJ@��]���M@[;�	��11eʴ�e�^��n��1�➪�� G�xGpB����'q�G �D�ۓU\��w����5�ǌ�a�޼L���ʝz�"��aJ�LX��cq�$.����ȵ���,H7G>�7�X�Vk�	8���Ǭ ~�a�F!�4IF�)��;�t;�f�V�%
ik���;���n��3�d���]�:����7��ٹ�Wy%��w@�4R\�����1�І�����B��������)#�jd�={��VJ�T���Y5f�\�Kr��W�yL<��\y�=�nY[����h��;�e������n����\t�):���5I�t��gV약ٚ�z�в "���of��4^̱�=�0�[����uuU'��+R����U����9(d���^���p�u�G��?l<v_�zu���Z�}�N�������}0��#�E|��?��>o��#�,��~���o��%,�}���%W������w���0m�L���'Sڬ�EUs/b�)p=�m�c�).z�5��x����]�f-?7s��E����������+�!���[v~�]�>5�Z���dN�g4���;�)�B�|��W�J~f�;V�{ߧ�b�������մ�f��f����t���9����V��l�I��Y��(��y�/c����K�T8��Z���Hg��O��V��<=���go�=	g[�'�� ��ρ��s����ݢd�wgGn��i�*���Y\t�}iò����yq�K��8^��
�(aJiZ,�D`����ˁ�㮱�u�^��KчѶM�qBW^��ri���nMb��%,��\������i��On.���Ρ��{��fNg�/�tI�4p��tf�k9o]\R[�u"���������4&;V��7�W�qx��c(`5h�9�t��������o.q�=W5����B�����t�@f�ƞ��'7?;w����w}�ө��e��[Q��o�����U�m����h�hJġJ�޴�n��7�wY�~o�u׷���Q����>M��y���?�]ӂa��[�����@����WUC�.ݵ�B6m9Mg���}]��}�~L�٫����;v���B���s�ښ8�!� ˧O�+��_�rc��E}���;��љ���W��hM���2x6��lݩ�b{�f�=�\Y���g=/����b��{�W��n�2I\�oN��E��/A]0F������aA����~瓵�!(լo�}k����ь�8�?pˑ�j��
aQA�O�&w���"��e~T۔C�E׫EEEy��l�c�נlp 4�t@~�y�%��CO�oߊ��V�_��e�߇����_�_h���#��i)1=������߸zݮ_ᗁ�:_n�5'�}����8�8rT�6�s�����ʡ2����Ƕ���������R!�.�߇��^������=}~�ivvٶ٬~'ж`r��4��?��Ud�ee���,|۶m")�3tlܪaY��qw��.`e��Qj��F��N�x�������`�5�<]�\�9%4 PK   j
mWN3_�	  ,K     jsons/user_defined.json�[]o��+=��� ��y�s�qbıo�"(�_��*ZU��A�{g��r���PB��^�-���%��pf��>Z~������}��gQV��,F�їrq_73�)O��~��?����������g?\&�H��D%��]�����aY�5�o����'�?�?�Gu�O�;�9Ɍ�%SN�	[0_S� 3q�{|��r�*�^弼��|��W��s"|:���s�zv1��������y}?��o�f�s�N�%�g�����vL��k���aeV��_+|��Eq�\Ԉ�K������7���-*H�UF��65���W���,��,����NCV��L��u�c�M �|~����/����#�N&�r��	^�=���6ƇU�(���E3/�z��V�y3��I����{}��\�{߬fE2if�2_6��C��f�bJx`�J`�(`Pf�\٬(��?� ���ƹ�?�Eʟy���(�J��Տ����2=�[��6`����}��IF�]̖�bV.)��e��Y�3Ud�|i/x�L�iW�
<A5���s�T2����W�0F��K�2��a�ě�� �fD	����_k�%q�E)�S�2�y.Xڃ�
�;xJ�Rg��NK�T�S� KreR.A���$�;n�y�|-@��`+ \5���H���;��ȣ�:d2^�d��j~�Գ�zڐb�%8ȌeJr�|�c�����p-���#O��(ޤ�z]�������x\���֖L`��oX�nc�u~W�M�;������gob��9^__%����&Q�H�J!�/Ӑ��ZdMv&��,�^�sv�|�%��\�����)VӒ�tBZ��P2ȌG�$�X���d��B� �NG��8fiƊ�4��X�6�!�(�`,��F��I3��6�Ƹކ���-A�v��m\�,"|��`7Idx(}��j���32S/�$�1���dݟ���'��S8���.d�2y����瓳"̱$�xs�k*�6/0�J3��	�RNcl~�7S�iՠ�B�No�����%7� �X	�*-Ş�8���oL��t�L�k�9L˟��%��j�M�%��Ѷ���SHf*-�*+�7EQ!�*Ue�Ǵ(�V�I��} ������k-�X��
�Ҿ�PDa/��l�%B^ۮ�a�ʗ�T��w��^~K���=���i���&\�q��͐ �g9��*;F3x�f|ꥵ�S3��؀�`(���
a�{ؓ?���pu�!F<�?qX�ñ%s��D�/19���8"�A�"٠���9�\�dE��L��e����ܶesf������r�$)�0ά��]���+~�����P�N�\'�%yY�&Yo���$/Ů1�Wa�<P���d�,
R����*��k��!j'+��(�B+e�1�v�ŕ]�I�y��Xt��к�~f�_�{��z���˰�)�Z��I�A�$[rW�g�����233V�97�92hV^A��O$���A_�\�Ϛvm��&�Rsk�ti�4�M�U�[�>𝼉\ij����e�==��
Q'���'��ڞ��(�6SA�
��2�aS3�lXV���)𴦉w�w_�،E��4��)�	��
-)����5���	����u��o=^�dv�l
�;�ܺ�G+�K�cN-W�L��1��lY��W�9wL�B���[�j�s���XtI�1TcdK�����m��}�Gk����Z�z�۫�����՛�'�I�>���(FAQq/8k�=XT���*H��J[P�>&�Q�)̦^�y#��X�b�Kqk�n����n���#��my5�O�8��%NG?)���Rњ�my��1n��7ͣ�x��?�-qN���8��nJ��&a��@'`�n�w��|���}/�*�]�|u}%!���/* :c2���K���c�W�
�����m
<�N�I���/O�[uH�	��rr���Ri��s�r�ܮ��6�Ї�ͤg��p��t��$٦�<�C�\L���GP������P�f���)�ma���n7f�'�(d*���RPݢ5��w��o�����u���zƐ����c����bI�x��ɋ��o�)H�E�U����� UǕ	�v��N�����d���d�Ժ9�n��_�>�%��e 
�X���&�k�R:ˏ�$�d�E�}@��2)>������޺a9���<b�ޕ�~�G�Gy�ˑl��Or�C���"��p�&}�y�q�x�1���lŌ�4�̔/�c/
<�5)�7�{�)�齭�]��D���X٨�+c�t(�O���Rp����g��~G��f�5�a����EP'�}��ޏԏ� �ӷ��l��g٭���,t��䅾�/�v&��x����w@K��p�ɧ��7�'a���+�Z���2W���J�,H(����p��1�U(�R�%y�7�c���N��{�A�9�
#ݞ��|�sY��.ܐ�>���B�D�	
���bu���Tk����?PK
   j
mWݵ�2>  ��                  cirkitFile.jsonPK
   �cW�����8 �I /             _>  images/13784fae-2b69-4ff3-9746-a43cbc14e23a.pngPK
   �cW��*��~ ̋ /             \w images/243361b7-2241-4a0b-aa59-149fc34d5bc9.pngPK
   �cW�>|�2� � /             �� images/2cacff52-a01f-447b-a47f-67011eb49dd1.pngPK
   �cWL̔���  � /             � images/37b4a41f-4938-46b6-a864-47b2117c0019.pngPK
   �cW�[0E  /             � images/42df0910-34e4-4e6b-8fa3-2ad2f5724f59.pngPK
   �cW��cH�1 &7 /             �� images/4657de38-a294-4f46-8901-aa5929bd88a8.pngPK
   �cW~�޴� �# /             �� images/51dc5037-8d6b-4f3e-a32e-636e17d8257a.pngPK
   �cW]*�Ļ� �� /             �� images/5241023b-b430-49fc-8631-1e6053993f23.pngPK
   �cW�����  -�  /             �� images/6bda90e9-5ec7-4d98-9c70-49b6fbff5641.pngPK
   �cW�{0n_C N /             �� images/7ec862db-5bbc-4dbd-b9e6-0d0e46cb58fd.pngPK
   �cW	��t bv /             e� images/a4ba225b-3a91-4e5e-8458-60f0fa258431.pngPK
   �cWh��~� ˴ /             �L images/ab527b7f-4192-4732-8642-2eb32cc47bdd.pngPK
   �cW�Q9lpz g~ /             �� images/b53b9fe2-18b9-4e15-8ac2-a2240bce23fb.pngPK
   �cW�ADE O /             �s images/be117233-6f51-4efb-b1df-934e4f712848.pngPK
   �cW���/�� Z� /             Nu# images/d3087b83-655e-4811-b17d-9d66f7a3b2a5.pngPK
   �cW<�� � /             <& images/d3b60164-5006-402c-a3a5-273a0eda4daa.pngPK
   �cW>R���5 �= /             m!' images/e1c0e916-28de-44d8-b600-7ef9d9f2b881.pngPK
   �cW�!ߔ�� @� /             QW( images/f1137482-0179-4042-abd2-21e421d54476.pngPK
   �cW䬂'�G �U /             U!* images/fc51afbd-40d4-4045-8777-933d8523ba7c.pngPK
   j
mWN3_�	  ,K               ii+ jsons/user_defined.jsonPK      i  qs+   